/* verilator lint_off UNUSED */
module IDU(
  input  [63:0] io_pc
);
endmodule
/* verilator lint_on UNUSED */
