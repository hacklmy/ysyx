module AXI(
  input         clock,
  input         reset,
  input  [31:0] io_axi_in_araddr,
  input         io_axi_in_arvalid,
  input         io_axi_in_rready,
  input  [31:0] io_axi_in_awaddr,
  input         io_axi_in_awvalid,
  input  [31:0] io_axi_in_wdata,
  input  [7:0]  io_axi_in_wstrb,
  input         io_axi_in_wvalid,
  input         io_axi_in_bready,
  output        io_axi_out_arready,
  output [63:0] io_axi_out_rdata,
  output        io_axi_out_rvalid,
  output        io_axi_out_awready,
  output        io_axi_out_wready,
  output        io_axi_out_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] Mem_modle_Raddr; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Rdata; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Waddr; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Wdata; // @[AXI.scala 26:27]
  wire [7:0] Mem_modle_Wmask; // @[AXI.scala 26:27]
  wire  Mem_modle_Write_en; // @[AXI.scala 26:27]
  wire  Mem_modle_Read_en; // @[AXI.scala 26:27]
  reg  axi_awready; // @[AXI.scala 13:30]
  reg  axi_wready; // @[AXI.scala 14:29]
  reg  axi_bvalid; // @[AXI.scala 17:29]
  reg  axi_arready; // @[AXI.scala 19:30]
  reg  axi_rvalid; // @[AXI.scala 21:29]
  reg [2:0] state; // @[AXI.scala 24:24]
  wire  _GEN_1 = io_axi_in_arvalid ? 1'h0 : axi_arready; // @[AXI.scala 49:42 51:29 19:30]
  wire  _GEN_2 = io_axi_in_arvalid | axi_rvalid; // @[AXI.scala 49:42 52:28 21:29]
  wire  _GEN_4 = io_axi_in_awvalid & io_axi_in_wvalid ? 1'h0 : axi_awready; // @[AXI.scala 39:56 41:29 13:30]
  wire  _GEN_5 = io_axi_in_awvalid & io_axi_in_wvalid ? 1'h0 : axi_wready; // @[AXI.scala 39:56 42:28 14:29]
  wire  _GEN_6 = io_axi_in_awvalid & io_axi_in_wvalid | axi_bvalid; // @[AXI.scala 39:56 43:28 17:29]
  wire  _GEN_7 = io_axi_in_awvalid & io_axi_in_wvalid ? axi_arready : _GEN_1; // @[AXI.scala 19:30 39:56]
  wire  _GEN_11 = io_axi_in_bready | axi_awready; // @[AXI.scala 56:35 59:29 13:30]
  wire  _GEN_12 = io_axi_in_bready | axi_wready; // @[AXI.scala 56:35 60:28 14:29]
  wire [2:0] _GEN_13 = io_axi_in_rready ? 3'h0 : state; // @[AXI.scala 64:35 65:23 24:24]
  wire  _GEN_14 = io_axi_in_rready | axi_arready; // @[AXI.scala 64:35 66:29 19:30]
  wire  _GEN_15 = io_axi_in_rready ? 1'h0 : axi_rvalid; // @[AXI.scala 64:35 67:28 21:29]
  wire  _GEN_17 = 3'h4 == state ? _GEN_14 : axi_arready; // @[AXI.scala 37:18 19:30]
  wire  _GEN_21 = 3'h3 == state ? _GEN_11 : axi_awready; // @[AXI.scala 37:18 13:30]
  wire  _GEN_22 = 3'h3 == state ? _GEN_12 : axi_wready; // @[AXI.scala 37:18 14:29]
  wire  _GEN_23 = 3'h3 == state ? axi_arready : _GEN_17; // @[AXI.scala 37:18 19:30]
  wire  _GEN_26 = 3'h0 == state ? _GEN_4 : _GEN_21; // @[AXI.scala 37:18]
  wire  _GEN_27 = 3'h0 == state ? _GEN_5 : _GEN_22; // @[AXI.scala 37:18]
  wire  _GEN_29 = 3'h0 == state ? _GEN_7 : _GEN_23; // @[AXI.scala 37:18]
  MEM Mem_modle ( // @[AXI.scala 26:27]
    .Raddr(Mem_modle_Raddr),
    .Rdata(Mem_modle_Rdata),
    .Waddr(Mem_modle_Waddr),
    .Wdata(Mem_modle_Wdata),
    .Wmask(Mem_modle_Wmask),
    .Write_en(Mem_modle_Write_en),
    .Read_en(Mem_modle_Read_en)
  );
  assign io_axi_out_arready = axi_arready; // @[AXI.scala 71:24]
  assign io_axi_out_rdata = Mem_modle_Rdata; // @[AXI.scala 72:22]
  assign io_axi_out_rvalid = axi_rvalid; // @[AXI.scala 73:23]
  assign io_axi_out_awready = axi_awready; // @[AXI.scala 74:24]
  assign io_axi_out_wready = axi_wready; // @[AXI.scala 75:23]
  assign io_axi_out_bvalid = axi_bvalid; // @[AXI.scala 76:23]
  assign Mem_modle_Raddr = {32'h0,io_axi_in_araddr}; // @[Cat.scala 31:58]
  assign Mem_modle_Waddr = {{32'd0}, io_axi_in_awaddr}; // @[AXI.scala 28:24]
  assign Mem_modle_Wdata = {{32'd0}, io_axi_in_wdata}; // @[AXI.scala 29:24]
  assign Mem_modle_Wmask = io_axi_in_wstrb; // @[AXI.scala 30:24]
  assign Mem_modle_Write_en = axi_wready & io_axi_in_wvalid; // @[AXI.scala 31:48]
  assign Mem_modle_Read_en = axi_arready & io_axi_in_arvalid; // @[AXI.scala 32:48]
  always @(posedge clock) begin
    axi_awready <= reset | _GEN_26; // @[AXI.scala 13:{30,30}]
    axi_wready <= reset | _GEN_27; // @[AXI.scala 14:{29,29}]
    if (reset) begin // @[AXI.scala 17:29]
      axi_bvalid <= 1'h0; // @[AXI.scala 17:29]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      axi_bvalid <= _GEN_6;
    end else if (3'h3 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_bready) begin // @[AXI.scala 56:35]
        axi_bvalid <= 1'h0; // @[AXI.scala 58:28]
      end
    end
    axi_arready <= reset | _GEN_29; // @[AXI.scala 19:{30,30}]
    if (reset) begin // @[AXI.scala 21:29]
      axi_rvalid <= 1'h0; // @[AXI.scala 21:29]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      if (!(io_axi_in_awvalid & io_axi_in_wvalid)) begin // @[AXI.scala 39:56]
        axi_rvalid <= _GEN_2;
      end
    end else if (!(3'h3 == state)) begin // @[AXI.scala 37:18]
      if (3'h4 == state) begin // @[AXI.scala 37:18]
        axi_rvalid <= _GEN_15;
      end
    end
    if (reset) begin // @[AXI.scala 24:24]
      state <= 3'h0; // @[AXI.scala 24:24]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_awvalid & io_axi_in_wvalid) begin // @[AXI.scala 39:56]
        state <= 3'h3; // @[AXI.scala 40:23]
      end else if (io_axi_in_arvalid) begin // @[AXI.scala 49:42]
        state <= 3'h4; // @[AXI.scala 50:23]
      end
    end else if (3'h3 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_bready) begin // @[AXI.scala 56:35]
        state <= 3'h0; // @[AXI.scala 57:23]
      end
    end else if (3'h4 == state) begin // @[AXI.scala 37:18]
      state <= _GEN_13;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_awready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  axi_wready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  axi_bvalid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  axi_arready = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  axi_rvalid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSU(
  input         clock,
  input         reset,
  input         io_inst_store,
  input         io_inst_load,
  input  [31:0] io_mem_addr,
  input  [63:0] io_mem_wdata,
  input  [7:0]  io_mem_wstrb,
  output [63:0] io_mem_rdata,
  input         io_axi_in_arready,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  input         io_axi_in_awready,
  input         io_axi_in_wready,
  input         io_axi_in_bvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  output [31:0] io_axi_out_awaddr,
  output        io_axi_out_awvalid,
  output [31:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid,
  output        io_axi_out_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  axi_arvalid; // @[LSU.scala 19:30]
  reg  axi_rready; // @[LSU.scala 22:29]
  reg  axi_awvalid; // @[LSU.scala 23:30]
  reg  axi_wvalid; // @[LSU.scala 24:29]
  reg  axi_bready; // @[LSU.scala 25:29]
  reg [1:0] state; // @[LSU.scala 28:24]
  wire  _GEN_1 = io_inst_store | axi_awvalid; // @[LSU.scala 36:38 38:29 23:30]
  wire  _GEN_2 = io_inst_store | axi_wvalid; // @[LSU.scala 36:38 39:28 24:29]
  wire  _GEN_3 = io_inst_store | axi_bready; // @[LSU.scala 36:38 40:28 25:29]
  wire  _GEN_5 = io_inst_load | axi_arvalid; // @[LSU.scala 32:31 34:29 19:30]
  wire  _GEN_6 = io_inst_load | axi_rready; // @[LSU.scala 32:31 35:28 22:29]
  wire  _GEN_9 = io_inst_load ? axi_bready : _GEN_3; // @[LSU.scala 25:29 32:31]
  wire  _GEN_11 = io_axi_in_bvalid ? 1'h0 : axi_bready; // @[LSU.scala 44:35 46:28 25:29]
  wire  _GEN_14 = io_axi_in_arready ? 1'h0 : axi_arvalid; // @[LSU.scala 56:36 57:29 19:30]
  wire [1:0] _GEN_15 = io_axi_in_rvalid ? 2'h0 : state; // @[LSU.scala 59:35 60:23 28:24]
  wire  _GEN_16 = io_axi_in_rvalid ? 1'h0 : axi_rready; // @[LSU.scala 59:35 61:28 22:29]
  wire  _GEN_19 = 2'h2 == state ? _GEN_16 : axi_rready; // @[LSU.scala 30:18 22:29]
  wire  _GEN_21 = 2'h1 == state ? _GEN_11 : axi_bready; // @[LSU.scala 30:18 25:29]
  wire  _GEN_25 = 2'h1 == state ? axi_rready : _GEN_19; // @[LSU.scala 30:18 22:29]
  wire  _GEN_28 = 2'h0 == state ? _GEN_6 : _GEN_25; // @[LSU.scala 30:18]
  wire  _GEN_31 = 2'h0 == state ? _GEN_9 : _GEN_21; // @[LSU.scala 30:18]
  assign io_mem_rdata = io_axi_in_rdata; // @[LSU.scala 72:18]
  assign io_axi_out_araddr = io_mem_addr; // @[LSU.scala 73:23]
  assign io_axi_out_arvalid = axi_arvalid; // @[LSU.scala 74:24]
  assign io_axi_out_rready = axi_rready; // @[LSU.scala 75:23]
  assign io_axi_out_awaddr = io_mem_addr; // @[LSU.scala 76:23]
  assign io_axi_out_awvalid = axi_awvalid; // @[LSU.scala 77:24]
  assign io_axi_out_wdata = io_mem_wdata[31:0]; // @[LSU.scala 78:22]
  assign io_axi_out_wstrb = io_mem_wstrb; // @[LSU.scala 79:22]
  assign io_axi_out_wvalid = axi_wvalid; // @[LSU.scala 80:23]
  assign io_axi_out_bready = axi_bready; // @[LSU.scala 81:23]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 19:30]
      axi_arvalid <= 1'h0; // @[LSU.scala 19:30]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      axi_arvalid <= _GEN_5;
    end else if (!(2'h1 == state)) begin // @[LSU.scala 30:18]
      if (2'h2 == state) begin // @[LSU.scala 30:18]
        axi_arvalid <= _GEN_14;
      end
    end
    axi_rready <= reset | _GEN_28; // @[LSU.scala 22:{29,29}]
    if (reset) begin // @[LSU.scala 23:30]
      axi_awvalid <= 1'h0; // @[LSU.scala 23:30]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (!(io_inst_load)) begin // @[LSU.scala 32:31]
        axi_awvalid <= _GEN_1;
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_awready) begin // @[LSU.scala 51:36]
        axi_awvalid <= 1'h0; // @[LSU.scala 52:29]
      end
    end
    if (reset) begin // @[LSU.scala 24:29]
      axi_wvalid <= 1'h0; // @[LSU.scala 24:29]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (!(io_inst_load)) begin // @[LSU.scala 32:31]
        axi_wvalid <= _GEN_2;
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_wready) begin // @[LSU.scala 48:35]
        axi_wvalid <= 1'h0; // @[LSU.scala 49:28]
      end
    end
    axi_bready <= reset | _GEN_31; // @[LSU.scala 25:{29,29}]
    if (reset) begin // @[LSU.scala 28:24]
      state <= 2'h0; // @[LSU.scala 28:24]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (io_inst_load) begin // @[LSU.scala 32:31]
        state <= 2'h2; // @[LSU.scala 33:23]
      end else if (io_inst_store) begin // @[LSU.scala 36:38]
        state <= 2'h1; // @[LSU.scala 37:23]
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_bvalid) begin // @[LSU.scala 44:35]
        state <= 2'h0; // @[LSU.scala 45:23]
      end
    end else if (2'h2 == state) begin // @[LSU.scala 30:18]
      state <= _GEN_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_arvalid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  axi_rready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  axi_awvalid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  axi_wvalid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  axi_bready = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI_ARBITER(
  input         clock,
  input         reset,
  input  [31:0] io_ifu_axi_in_araddr,
  input         io_ifu_axi_in_arvalid,
  input         io_ifu_axi_in_rready,
  output [63:0] io_ifu_axi_out_rdata,
  output        io_ifu_axi_out_rvalid,
  input  [31:0] io_lsu_axi_in_araddr,
  input         io_lsu_axi_in_arvalid,
  input         io_lsu_axi_in_rready,
  input  [31:0] io_lsu_axi_in_awaddr,
  input         io_lsu_axi_in_awvalid,
  input  [31:0] io_lsu_axi_in_wdata,
  input  [7:0]  io_lsu_axi_in_wstrb,
  input         io_lsu_axi_in_wvalid,
  input         io_lsu_axi_in_bready,
  output        io_lsu_axi_out_arready,
  output [63:0] io_lsu_axi_out_rdata,
  output        io_lsu_axi_out_rvalid,
  output        io_lsu_axi_out_awready,
  output        io_lsu_axi_out_wready,
  output        io_lsu_axi_out_bvalid,
  input         io_axi_in_arready,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  input         io_axi_in_awready,
  input         io_axi_in_wready,
  input         io_axi_in_bvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  output [31:0] io_axi_out_awaddr,
  output        io_axi_out_awvalid,
  output [31:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid,
  output        io_axi_out_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[axi_arbiter.scala 18:24]
  wire [1:0] _GEN_0 = io_ifu_axi_in_arvalid ? 2'h1 : state; // @[axi_arbiter.scala 51:46 52:23 18:24]
  wire [31:0] _GEN_1 = io_ifu_axi_in_arvalid ? io_ifu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 51:46 53:28 57:28]
  wire  _GEN_3 = io_ifu_axi_in_arvalid & io_ifu_axi_in_rready; // @[axi_arbiter.scala 51:46 53:28 57:28]
  wire [63:0] _GEN_11 = io_ifu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 51:46 54:32 59:32]
  wire  _GEN_12 = io_ifu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 51:46 54:32 59:32]
  wire [31:0] _GEN_23 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_araddr : _GEN_1; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_24 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_arvalid : io_ifu_axi_in_arvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_25 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_rready : _GEN_3; // @[axi_arbiter.scala 46:46 48:28]
  wire [31:0] _GEN_26 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_27 = io_lsu_axi_in_arvalid & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire [31:0] _GEN_28 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wdata : 32'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire [7:0] _GEN_29 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_30 = io_lsu_axi_in_arvalid & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_31 = io_lsu_axi_in_arvalid & io_lsu_axi_in_bready; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_32 = io_lsu_axi_in_arvalid & io_axi_in_arready; // @[axi_arbiter.scala 46:46 49:32]
  wire [63:0] _GEN_33 = io_lsu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_34 = io_lsu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_35 = io_lsu_axi_in_arvalid & io_axi_in_awready; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_36 = io_lsu_axi_in_arvalid & io_axi_in_wready; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_37 = io_lsu_axi_in_arvalid & io_axi_in_bvalid; // @[axi_arbiter.scala 46:46 49:32]
  wire [63:0] _GEN_39 = io_lsu_axi_in_arvalid ? 64'h0 : _GEN_11; // @[axi_arbiter.scala 46:46 50:32]
  wire  _GEN_40 = io_lsu_axi_in_arvalid ? 1'h0 : _GEN_12; // @[axi_arbiter.scala 46:46 50:32]
  wire [31:0] _GEN_45 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_araddr : _GEN_23; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_46 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_arvalid : _GEN_24; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_47 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_rready : _GEN_25; // @[axi_arbiter.scala 41:40 43:28]
  wire [31:0] _GEN_48 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awaddr : _GEN_26; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_49 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awvalid : _GEN_27; // @[axi_arbiter.scala 41:40 43:28]
  wire [31:0] _GEN_50 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wdata : _GEN_28; // @[axi_arbiter.scala 41:40 43:28]
  wire [7:0] _GEN_51 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wstrb : _GEN_29; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_52 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wvalid : _GEN_30; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_53 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_bready : _GEN_31; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_54 = io_lsu_axi_in_awvalid ? io_axi_in_arready : _GEN_32; // @[axi_arbiter.scala 41:40 44:32]
  wire [63:0] _GEN_55 = io_lsu_axi_in_awvalid ? io_axi_in_rdata : _GEN_33; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_56 = io_lsu_axi_in_awvalid ? io_axi_in_rvalid : _GEN_34; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_57 = io_lsu_axi_in_awvalid ? io_axi_in_awready : _GEN_35; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_58 = io_lsu_axi_in_awvalid ? io_axi_in_wready : _GEN_36; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_59 = io_lsu_axi_in_awvalid ? io_axi_in_bvalid : _GEN_37; // @[axi_arbiter.scala 41:40 44:32]
  wire [63:0] _GEN_61 = io_lsu_axi_in_awvalid ? 64'h0 : _GEN_39; // @[axi_arbiter.scala 41:40 45:32]
  wire  _GEN_62 = io_lsu_axi_in_awvalid ? 1'h0 : _GEN_40; // @[axi_arbiter.scala 41:40 45:32]
  wire [1:0] _GEN_67 = io_lsu_axi_out_rvalid & io_lsu_axi_in_rready ? 2'h0 : state; // @[axi_arbiter.scala 74:64 75:23 18:24]
  wire [1:0] _GEN_68 = io_lsu_axi_out_bvalid & io_lsu_axi_in_bready ? 2'h0 : state; // @[axi_arbiter.scala 82:64 83:23 18:24]
  wire [31:0] _GEN_69 = state == 2'h3 ? io_lsu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_70 = state == 2'h3 & io_lsu_axi_in_arvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_71 = state == 2'h3 & io_lsu_axi_in_rready; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [31:0] _GEN_72 = state == 2'h3 ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_73 = state == 2'h3 & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [31:0] _GEN_74 = state == 2'h3 ? io_lsu_axi_in_wdata : 32'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [7:0] _GEN_75 = state == 2'h3 ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_76 = state == 2'h3 & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_77 = state == 2'h3 & io_lsu_axi_in_bready; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_78 = state == 2'h3 & io_axi_in_arready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire [63:0] _GEN_79 = state == 2'h3 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_80 = state == 2'h3 & io_axi_in_rvalid; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_81 = state == 2'h3 & io_axi_in_awready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_82 = state == 2'h3 & io_axi_in_wready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_83 = state == 2'h3 & io_axi_in_bvalid; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire [1:0] _GEN_90 = state == 2'h3 ? _GEN_68 : state; // @[axi_arbiter.scala 18:24 78:39]
  wire [31:0] _GEN_91 = state == 2'h2 ? io_lsu_axi_in_araddr : _GEN_69; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_92 = state == 2'h2 ? io_lsu_axi_in_arvalid : _GEN_70; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_93 = state == 2'h2 ? io_lsu_axi_in_rready : _GEN_71; // @[axi_arbiter.scala 70:39 71:24]
  wire [31:0] _GEN_94 = state == 2'h2 ? io_lsu_axi_in_awaddr : _GEN_72; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_95 = state == 2'h2 ? io_lsu_axi_in_awvalid : _GEN_73; // @[axi_arbiter.scala 70:39 71:24]
  wire [31:0] _GEN_96 = state == 2'h2 ? io_lsu_axi_in_wdata : _GEN_74; // @[axi_arbiter.scala 70:39 71:24]
  wire [7:0] _GEN_97 = state == 2'h2 ? io_lsu_axi_in_wstrb : _GEN_75; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_98 = state == 2'h2 ? io_lsu_axi_in_wvalid : _GEN_76; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_99 = state == 2'h2 ? io_lsu_axi_in_bready : _GEN_77; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_100 = state == 2'h2 ? io_axi_in_arready : _GEN_78; // @[axi_arbiter.scala 70:39 72:28]
  wire [63:0] _GEN_101 = state == 2'h2 ? io_axi_in_rdata : _GEN_79; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_102 = state == 2'h2 ? io_axi_in_rvalid : _GEN_80; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_103 = state == 2'h2 ? io_axi_in_awready : _GEN_81; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_104 = state == 2'h2 ? io_axi_in_wready : _GEN_82; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_105 = state == 2'h2 ? io_axi_in_bvalid : _GEN_83; // @[axi_arbiter.scala 70:39 72:28]
  wire [31:0] _GEN_113 = state == 2'h1 ? io_ifu_axi_in_araddr : _GEN_91; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_114 = state == 2'h1 ? io_ifu_axi_in_arvalid : _GEN_92; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_115 = state == 2'h1 ? io_ifu_axi_in_rready : _GEN_93; // @[axi_arbiter.scala 62:39 63:24]
  wire [31:0] _GEN_116 = state == 2'h1 ? 32'h0 : _GEN_94; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_117 = state == 2'h1 ? 1'h0 : _GEN_95; // @[axi_arbiter.scala 62:39 63:24]
  wire [31:0] _GEN_118 = state == 2'h1 ? 32'h0 : _GEN_96; // @[axi_arbiter.scala 62:39 63:24]
  wire [7:0] _GEN_119 = state == 2'h1 ? 8'h0 : _GEN_97; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_120 = state == 2'h1 ? 1'h0 : _GEN_98; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_121 = state == 2'h1 ? 1'h0 : _GEN_99; // @[axi_arbiter.scala 62:39 63:24]
  wire [63:0] _GEN_123 = state == 2'h1 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 62:39 64:28]
  wire  _GEN_124 = state == 2'h1 & io_axi_in_rvalid; // @[axi_arbiter.scala 62:39 64:28]
  wire  _GEN_128 = state == 2'h1 ? 1'h0 : _GEN_100; // @[axi_arbiter.scala 62:39 65:28]
  wire [63:0] _GEN_129 = state == 2'h1 ? 64'h0 : _GEN_101; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_130 = state == 2'h1 ? 1'h0 : _GEN_102; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_131 = state == 2'h1 ? 1'h0 : _GEN_103; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_132 = state == 2'h1 ? 1'h0 : _GEN_104; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_133 = state == 2'h1 ? 1'h0 : _GEN_105; // @[axi_arbiter.scala 62:39 65:28]
  assign io_ifu_axi_out_rdata = state == 2'h0 ? _GEN_61 : _GEN_123; // @[axi_arbiter.scala 40:27]
  assign io_ifu_axi_out_rvalid = state == 2'h0 ? _GEN_62 : _GEN_124; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_arready = state == 2'h0 ? _GEN_54 : _GEN_128; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_rdata = state == 2'h0 ? _GEN_55 : _GEN_129; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_rvalid = state == 2'h0 ? _GEN_56 : _GEN_130; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_awready = state == 2'h0 ? _GEN_57 : _GEN_131; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_wready = state == 2'h0 ? _GEN_58 : _GEN_132; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_bvalid = state == 2'h0 ? _GEN_59 : _GEN_133; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_araddr = state == 2'h0 ? _GEN_45 : _GEN_113; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_arvalid = state == 2'h0 ? _GEN_46 : _GEN_114; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_rready = state == 2'h0 ? _GEN_47 : _GEN_115; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_awaddr = state == 2'h0 ? _GEN_48 : _GEN_116; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_awvalid = state == 2'h0 ? _GEN_49 : _GEN_117; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wdata = state == 2'h0 ? _GEN_50 : _GEN_118; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wstrb = state == 2'h0 ? _GEN_51 : _GEN_119; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wvalid = state == 2'h0 ? _GEN_52 : _GEN_120; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_bready = state == 2'h0 ? _GEN_53 : _GEN_121; // @[axi_arbiter.scala 40:27]
  always @(posedge clock) begin
    if (reset) begin // @[axi_arbiter.scala 18:24]
      state <= 2'h0; // @[axi_arbiter.scala 18:24]
    end else if (state == 2'h0) begin // @[axi_arbiter.scala 40:27]
      if (io_lsu_axi_in_awvalid) begin // @[axi_arbiter.scala 41:40]
        state <= 2'h3; // @[axi_arbiter.scala 42:23]
      end else if (io_lsu_axi_in_arvalid) begin // @[axi_arbiter.scala 46:46]
        state <= 2'h2; // @[axi_arbiter.scala 47:23]
      end else begin
        state <= _GEN_0;
      end
    end else if (state == 2'h1) begin // @[axi_arbiter.scala 62:39]
      if (io_ifu_axi_out_rvalid & io_ifu_axi_in_rready) begin // @[axi_arbiter.scala 66:64]
        state <= 2'h0; // @[axi_arbiter.scala 67:23]
      end
    end else if (state == 2'h2) begin // @[axi_arbiter.scala 70:39]
      state <= _GEN_67;
    end else begin
      state <= _GEN_90;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU_AXI(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_pc_valid,
  output        io_inst_valid,
  output [31:0] io_inst,
  output [31:0] io_inst_reg,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  inst_ready; // @[IFU_AXI.scala 19:29]
  wire  _GEN_0 = io_axi_in_rvalid & inst_ready ? 1'h0 : 1'h1; // @[IFU_AXI.scala 20:41 21:20 23:20]
  reg [31:0] inst_reg; // @[IFU_AXI.scala 25:27]
  assign io_inst_valid = io_axi_in_rvalid; // @[IFU_AXI.scala 43:19]
  assign io_inst = io_axi_in_rdata[31:0]; // @[IFU_AXI.scala 41:31]
  assign io_inst_reg = inst_reg; // @[IFU_AXI.scala 42:17]
  assign io_axi_out_araddr = io_pc[31:0]; // @[IFU_AXI.scala 31:31]
  assign io_axi_out_arvalid = io_pc_valid; // @[IFU_AXI.scala 32:24]
  assign io_axi_out_rready = inst_ready; // @[IFU_AXI.scala 33:23]
  always @(posedge clock) begin
    inst_ready <= reset | _GEN_0; // @[IFU_AXI.scala 19:{29,29}]
    if (reset) begin // @[IFU_AXI.scala 25:27]
      inst_reg <= 32'h0; // @[IFU_AXI.scala 25:27]
    end else if (io_axi_in_rvalid) begin // @[IFU_AXI.scala 26:27]
      inst_reg <= io_axi_in_rdata[31:0]; // @[IFU_AXI.scala 27:18]
    end else if (io_pc_valid) begin // @[IFU_AXI.scala 28:28]
      inst_reg <= 32'h0; // @[IFU_AXI.scala 29:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst_ready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  inst_reg = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module I_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_ifu_araddr,
  input         io_from_ifu_arvalid,
  input         io_from_ifu_rready,
  output [63:0] io_to_ifu_rdata,
  output        io_to_ifu_rvalid,
  output [31:0] io_to_axi_araddr,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [63:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_0_0; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_1; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_2; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_3; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_4; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_5; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_6; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_7; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_8; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_9; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_10; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_11; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_12; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_13; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_14; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_15; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_16; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_17; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_18; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_19; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_20; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_21; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_22; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_23; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_24; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_25; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_26; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_27; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_28; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_29; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_30; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_31; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_32; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_33; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_34; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_35; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_36; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_37; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_38; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_39; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_40; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_41; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_42; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_43; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_44; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_45; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_46; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_47; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_48; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_49; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_50; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_51; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_52; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_53; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_54; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_55; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_56; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_57; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_58; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_59; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_60; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_61; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_62; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_63; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_64; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_65; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_66; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_67; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_68; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_69; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_70; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_71; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_72; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_73; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_74; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_75; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_76; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_77; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_78; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_79; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_80; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_81; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_82; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_83; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_84; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_85; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_86; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_87; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_88; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_89; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_90; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_91; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_92; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_93; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_94; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_95; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_96; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_97; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_98; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_99; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_100; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_101; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_102; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_103; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_104; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_105; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_106; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_107; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_108; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_109; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_110; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_111; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_112; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_113; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_114; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_115; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_116; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_117; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_118; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_119; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_120; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_121; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_122; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_123; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_124; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_125; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_126; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_127; // @[i_cache.scala 17:24]
  reg [63:0] ram_1_0; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_1; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_2; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_3; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_4; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_5; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_6; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_7; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_8; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_9; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_10; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_11; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_12; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_13; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_14; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_15; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_16; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_17; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_18; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_19; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_20; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_21; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_22; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_23; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_24; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_25; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_26; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_27; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_28; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_29; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_30; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_31; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_32; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_33; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_34; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_35; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_36; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_37; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_38; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_39; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_40; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_41; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_42; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_43; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_44; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_45; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_46; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_47; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_48; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_49; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_50; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_51; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_52; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_53; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_54; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_55; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_56; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_57; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_58; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_59; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_60; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_61; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_62; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_63; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_64; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_65; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_66; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_67; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_68; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_69; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_70; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_71; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_72; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_73; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_74; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_75; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_76; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_77; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_78; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_79; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_80; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_81; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_82; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_83; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_84; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_85; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_86; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_87; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_88; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_89; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_90; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_91; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_92; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_93; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_94; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_95; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_96; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_97; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_98; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_99; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_100; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_101; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_102; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_103; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_104; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_105; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_106; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_107; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_108; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_109; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_110; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_111; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_112; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_113; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_114; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_115; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_116; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_117; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_118; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_119; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_120; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_121; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_122; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_123; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_124; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_125; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_126; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_127; // @[i_cache.scala 18:24]
  reg [31:0] tag_0_0; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_1; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_2; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_3; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_4; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_5; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_6; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_7; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_8; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_9; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_10; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_11; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_12; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_13; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_14; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_15; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_16; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_17; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_18; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_19; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_20; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_21; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_22; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_23; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_24; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_25; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_26; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_27; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_28; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_29; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_30; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_31; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_32; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_33; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_34; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_35; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_36; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_37; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_38; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_39; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_40; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_41; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_42; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_43; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_44; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_45; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_46; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_47; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_48; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_49; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_50; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_51; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_52; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_53; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_54; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_55; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_56; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_57; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_58; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_59; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_60; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_61; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_62; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_63; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_64; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_65; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_66; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_67; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_68; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_69; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_70; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_71; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_72; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_73; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_74; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_75; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_76; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_77; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_78; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_79; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_80; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_81; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_82; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_83; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_84; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_85; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_86; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_87; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_88; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_89; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_90; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_91; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_92; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_93; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_94; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_95; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_96; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_97; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_98; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_99; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_100; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_101; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_102; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_103; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_104; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_105; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_106; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_107; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_108; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_109; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_110; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_111; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_112; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_113; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_114; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_115; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_116; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_117; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_118; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_119; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_120; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_121; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_122; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_123; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_124; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_125; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_126; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_127; // @[i_cache.scala 19:24]
  reg [31:0] tag_1_0; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_1; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_2; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_3; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_4; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_5; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_6; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_7; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_8; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_9; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_10; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_11; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_12; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_13; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_14; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_15; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_16; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_17; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_18; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_19; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_20; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_21; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_22; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_23; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_24; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_25; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_26; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_27; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_28; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_29; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_30; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_31; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_32; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_33; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_34; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_35; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_36; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_37; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_38; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_39; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_40; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_41; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_42; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_43; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_44; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_45; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_46; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_47; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_48; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_49; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_50; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_51; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_52; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_53; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_54; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_55; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_56; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_57; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_58; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_59; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_60; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_61; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_62; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_63; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_64; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_65; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_66; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_67; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_68; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_69; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_70; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_71; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_72; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_73; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_74; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_75; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_76; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_77; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_78; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_79; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_80; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_81; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_82; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_83; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_84; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_85; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_86; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_87; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_88; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_89; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_90; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_91; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_92; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_93; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_94; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_95; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_96; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_97; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_98; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_99; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_100; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_101; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_102; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_103; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_104; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_105; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_106; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_107; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_108; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_109; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_110; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_111; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_112; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_113; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_114; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_115; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_116; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_117; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_118; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_119; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_120; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_121; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_122; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_123; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_124; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_125; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_126; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_127; // @[i_cache.scala 20:24]
  reg  valid_0_0; // @[i_cache.scala 21:26]
  reg  valid_0_1; // @[i_cache.scala 21:26]
  reg  valid_0_2; // @[i_cache.scala 21:26]
  reg  valid_0_3; // @[i_cache.scala 21:26]
  reg  valid_0_4; // @[i_cache.scala 21:26]
  reg  valid_0_5; // @[i_cache.scala 21:26]
  reg  valid_0_6; // @[i_cache.scala 21:26]
  reg  valid_0_7; // @[i_cache.scala 21:26]
  reg  valid_0_8; // @[i_cache.scala 21:26]
  reg  valid_0_9; // @[i_cache.scala 21:26]
  reg  valid_0_10; // @[i_cache.scala 21:26]
  reg  valid_0_11; // @[i_cache.scala 21:26]
  reg  valid_0_12; // @[i_cache.scala 21:26]
  reg  valid_0_13; // @[i_cache.scala 21:26]
  reg  valid_0_14; // @[i_cache.scala 21:26]
  reg  valid_0_15; // @[i_cache.scala 21:26]
  reg  valid_0_16; // @[i_cache.scala 21:26]
  reg  valid_0_17; // @[i_cache.scala 21:26]
  reg  valid_0_18; // @[i_cache.scala 21:26]
  reg  valid_0_19; // @[i_cache.scala 21:26]
  reg  valid_0_20; // @[i_cache.scala 21:26]
  reg  valid_0_21; // @[i_cache.scala 21:26]
  reg  valid_0_22; // @[i_cache.scala 21:26]
  reg  valid_0_23; // @[i_cache.scala 21:26]
  reg  valid_0_24; // @[i_cache.scala 21:26]
  reg  valid_0_25; // @[i_cache.scala 21:26]
  reg  valid_0_26; // @[i_cache.scala 21:26]
  reg  valid_0_27; // @[i_cache.scala 21:26]
  reg  valid_0_28; // @[i_cache.scala 21:26]
  reg  valid_0_29; // @[i_cache.scala 21:26]
  reg  valid_0_30; // @[i_cache.scala 21:26]
  reg  valid_0_31; // @[i_cache.scala 21:26]
  reg  valid_0_32; // @[i_cache.scala 21:26]
  reg  valid_0_33; // @[i_cache.scala 21:26]
  reg  valid_0_34; // @[i_cache.scala 21:26]
  reg  valid_0_35; // @[i_cache.scala 21:26]
  reg  valid_0_36; // @[i_cache.scala 21:26]
  reg  valid_0_37; // @[i_cache.scala 21:26]
  reg  valid_0_38; // @[i_cache.scala 21:26]
  reg  valid_0_39; // @[i_cache.scala 21:26]
  reg  valid_0_40; // @[i_cache.scala 21:26]
  reg  valid_0_41; // @[i_cache.scala 21:26]
  reg  valid_0_42; // @[i_cache.scala 21:26]
  reg  valid_0_43; // @[i_cache.scala 21:26]
  reg  valid_0_44; // @[i_cache.scala 21:26]
  reg  valid_0_45; // @[i_cache.scala 21:26]
  reg  valid_0_46; // @[i_cache.scala 21:26]
  reg  valid_0_47; // @[i_cache.scala 21:26]
  reg  valid_0_48; // @[i_cache.scala 21:26]
  reg  valid_0_49; // @[i_cache.scala 21:26]
  reg  valid_0_50; // @[i_cache.scala 21:26]
  reg  valid_0_51; // @[i_cache.scala 21:26]
  reg  valid_0_52; // @[i_cache.scala 21:26]
  reg  valid_0_53; // @[i_cache.scala 21:26]
  reg  valid_0_54; // @[i_cache.scala 21:26]
  reg  valid_0_55; // @[i_cache.scala 21:26]
  reg  valid_0_56; // @[i_cache.scala 21:26]
  reg  valid_0_57; // @[i_cache.scala 21:26]
  reg  valid_0_58; // @[i_cache.scala 21:26]
  reg  valid_0_59; // @[i_cache.scala 21:26]
  reg  valid_0_60; // @[i_cache.scala 21:26]
  reg  valid_0_61; // @[i_cache.scala 21:26]
  reg  valid_0_62; // @[i_cache.scala 21:26]
  reg  valid_0_63; // @[i_cache.scala 21:26]
  reg  valid_0_64; // @[i_cache.scala 21:26]
  reg  valid_0_65; // @[i_cache.scala 21:26]
  reg  valid_0_66; // @[i_cache.scala 21:26]
  reg  valid_0_67; // @[i_cache.scala 21:26]
  reg  valid_0_68; // @[i_cache.scala 21:26]
  reg  valid_0_69; // @[i_cache.scala 21:26]
  reg  valid_0_70; // @[i_cache.scala 21:26]
  reg  valid_0_71; // @[i_cache.scala 21:26]
  reg  valid_0_72; // @[i_cache.scala 21:26]
  reg  valid_0_73; // @[i_cache.scala 21:26]
  reg  valid_0_74; // @[i_cache.scala 21:26]
  reg  valid_0_75; // @[i_cache.scala 21:26]
  reg  valid_0_76; // @[i_cache.scala 21:26]
  reg  valid_0_77; // @[i_cache.scala 21:26]
  reg  valid_0_78; // @[i_cache.scala 21:26]
  reg  valid_0_79; // @[i_cache.scala 21:26]
  reg  valid_0_80; // @[i_cache.scala 21:26]
  reg  valid_0_81; // @[i_cache.scala 21:26]
  reg  valid_0_82; // @[i_cache.scala 21:26]
  reg  valid_0_83; // @[i_cache.scala 21:26]
  reg  valid_0_84; // @[i_cache.scala 21:26]
  reg  valid_0_85; // @[i_cache.scala 21:26]
  reg  valid_0_86; // @[i_cache.scala 21:26]
  reg  valid_0_87; // @[i_cache.scala 21:26]
  reg  valid_0_88; // @[i_cache.scala 21:26]
  reg  valid_0_89; // @[i_cache.scala 21:26]
  reg  valid_0_90; // @[i_cache.scala 21:26]
  reg  valid_0_91; // @[i_cache.scala 21:26]
  reg  valid_0_92; // @[i_cache.scala 21:26]
  reg  valid_0_93; // @[i_cache.scala 21:26]
  reg  valid_0_94; // @[i_cache.scala 21:26]
  reg  valid_0_95; // @[i_cache.scala 21:26]
  reg  valid_0_96; // @[i_cache.scala 21:26]
  reg  valid_0_97; // @[i_cache.scala 21:26]
  reg  valid_0_98; // @[i_cache.scala 21:26]
  reg  valid_0_99; // @[i_cache.scala 21:26]
  reg  valid_0_100; // @[i_cache.scala 21:26]
  reg  valid_0_101; // @[i_cache.scala 21:26]
  reg  valid_0_102; // @[i_cache.scala 21:26]
  reg  valid_0_103; // @[i_cache.scala 21:26]
  reg  valid_0_104; // @[i_cache.scala 21:26]
  reg  valid_0_105; // @[i_cache.scala 21:26]
  reg  valid_0_106; // @[i_cache.scala 21:26]
  reg  valid_0_107; // @[i_cache.scala 21:26]
  reg  valid_0_108; // @[i_cache.scala 21:26]
  reg  valid_0_109; // @[i_cache.scala 21:26]
  reg  valid_0_110; // @[i_cache.scala 21:26]
  reg  valid_0_111; // @[i_cache.scala 21:26]
  reg  valid_0_112; // @[i_cache.scala 21:26]
  reg  valid_0_113; // @[i_cache.scala 21:26]
  reg  valid_0_114; // @[i_cache.scala 21:26]
  reg  valid_0_115; // @[i_cache.scala 21:26]
  reg  valid_0_116; // @[i_cache.scala 21:26]
  reg  valid_0_117; // @[i_cache.scala 21:26]
  reg  valid_0_118; // @[i_cache.scala 21:26]
  reg  valid_0_119; // @[i_cache.scala 21:26]
  reg  valid_0_120; // @[i_cache.scala 21:26]
  reg  valid_0_121; // @[i_cache.scala 21:26]
  reg  valid_0_122; // @[i_cache.scala 21:26]
  reg  valid_0_123; // @[i_cache.scala 21:26]
  reg  valid_0_124; // @[i_cache.scala 21:26]
  reg  valid_0_125; // @[i_cache.scala 21:26]
  reg  valid_0_126; // @[i_cache.scala 21:26]
  reg  valid_0_127; // @[i_cache.scala 21:26]
  reg  valid_1_0; // @[i_cache.scala 22:26]
  reg  valid_1_1; // @[i_cache.scala 22:26]
  reg  valid_1_2; // @[i_cache.scala 22:26]
  reg  valid_1_3; // @[i_cache.scala 22:26]
  reg  valid_1_4; // @[i_cache.scala 22:26]
  reg  valid_1_5; // @[i_cache.scala 22:26]
  reg  valid_1_6; // @[i_cache.scala 22:26]
  reg  valid_1_7; // @[i_cache.scala 22:26]
  reg  valid_1_8; // @[i_cache.scala 22:26]
  reg  valid_1_9; // @[i_cache.scala 22:26]
  reg  valid_1_10; // @[i_cache.scala 22:26]
  reg  valid_1_11; // @[i_cache.scala 22:26]
  reg  valid_1_12; // @[i_cache.scala 22:26]
  reg  valid_1_13; // @[i_cache.scala 22:26]
  reg  valid_1_14; // @[i_cache.scala 22:26]
  reg  valid_1_15; // @[i_cache.scala 22:26]
  reg  valid_1_16; // @[i_cache.scala 22:26]
  reg  valid_1_17; // @[i_cache.scala 22:26]
  reg  valid_1_18; // @[i_cache.scala 22:26]
  reg  valid_1_19; // @[i_cache.scala 22:26]
  reg  valid_1_20; // @[i_cache.scala 22:26]
  reg  valid_1_21; // @[i_cache.scala 22:26]
  reg  valid_1_22; // @[i_cache.scala 22:26]
  reg  valid_1_23; // @[i_cache.scala 22:26]
  reg  valid_1_24; // @[i_cache.scala 22:26]
  reg  valid_1_25; // @[i_cache.scala 22:26]
  reg  valid_1_26; // @[i_cache.scala 22:26]
  reg  valid_1_27; // @[i_cache.scala 22:26]
  reg  valid_1_28; // @[i_cache.scala 22:26]
  reg  valid_1_29; // @[i_cache.scala 22:26]
  reg  valid_1_30; // @[i_cache.scala 22:26]
  reg  valid_1_31; // @[i_cache.scala 22:26]
  reg  valid_1_32; // @[i_cache.scala 22:26]
  reg  valid_1_33; // @[i_cache.scala 22:26]
  reg  valid_1_34; // @[i_cache.scala 22:26]
  reg  valid_1_35; // @[i_cache.scala 22:26]
  reg  valid_1_36; // @[i_cache.scala 22:26]
  reg  valid_1_37; // @[i_cache.scala 22:26]
  reg  valid_1_38; // @[i_cache.scala 22:26]
  reg  valid_1_39; // @[i_cache.scala 22:26]
  reg  valid_1_40; // @[i_cache.scala 22:26]
  reg  valid_1_41; // @[i_cache.scala 22:26]
  reg  valid_1_42; // @[i_cache.scala 22:26]
  reg  valid_1_43; // @[i_cache.scala 22:26]
  reg  valid_1_44; // @[i_cache.scala 22:26]
  reg  valid_1_45; // @[i_cache.scala 22:26]
  reg  valid_1_46; // @[i_cache.scala 22:26]
  reg  valid_1_47; // @[i_cache.scala 22:26]
  reg  valid_1_48; // @[i_cache.scala 22:26]
  reg  valid_1_49; // @[i_cache.scala 22:26]
  reg  valid_1_50; // @[i_cache.scala 22:26]
  reg  valid_1_51; // @[i_cache.scala 22:26]
  reg  valid_1_52; // @[i_cache.scala 22:26]
  reg  valid_1_53; // @[i_cache.scala 22:26]
  reg  valid_1_54; // @[i_cache.scala 22:26]
  reg  valid_1_55; // @[i_cache.scala 22:26]
  reg  valid_1_56; // @[i_cache.scala 22:26]
  reg  valid_1_57; // @[i_cache.scala 22:26]
  reg  valid_1_58; // @[i_cache.scala 22:26]
  reg  valid_1_59; // @[i_cache.scala 22:26]
  reg  valid_1_60; // @[i_cache.scala 22:26]
  reg  valid_1_61; // @[i_cache.scala 22:26]
  reg  valid_1_62; // @[i_cache.scala 22:26]
  reg  valid_1_63; // @[i_cache.scala 22:26]
  reg  valid_1_64; // @[i_cache.scala 22:26]
  reg  valid_1_65; // @[i_cache.scala 22:26]
  reg  valid_1_66; // @[i_cache.scala 22:26]
  reg  valid_1_67; // @[i_cache.scala 22:26]
  reg  valid_1_68; // @[i_cache.scala 22:26]
  reg  valid_1_69; // @[i_cache.scala 22:26]
  reg  valid_1_70; // @[i_cache.scala 22:26]
  reg  valid_1_71; // @[i_cache.scala 22:26]
  reg  valid_1_72; // @[i_cache.scala 22:26]
  reg  valid_1_73; // @[i_cache.scala 22:26]
  reg  valid_1_74; // @[i_cache.scala 22:26]
  reg  valid_1_75; // @[i_cache.scala 22:26]
  reg  valid_1_76; // @[i_cache.scala 22:26]
  reg  valid_1_77; // @[i_cache.scala 22:26]
  reg  valid_1_78; // @[i_cache.scala 22:26]
  reg  valid_1_79; // @[i_cache.scala 22:26]
  reg  valid_1_80; // @[i_cache.scala 22:26]
  reg  valid_1_81; // @[i_cache.scala 22:26]
  reg  valid_1_82; // @[i_cache.scala 22:26]
  reg  valid_1_83; // @[i_cache.scala 22:26]
  reg  valid_1_84; // @[i_cache.scala 22:26]
  reg  valid_1_85; // @[i_cache.scala 22:26]
  reg  valid_1_86; // @[i_cache.scala 22:26]
  reg  valid_1_87; // @[i_cache.scala 22:26]
  reg  valid_1_88; // @[i_cache.scala 22:26]
  reg  valid_1_89; // @[i_cache.scala 22:26]
  reg  valid_1_90; // @[i_cache.scala 22:26]
  reg  valid_1_91; // @[i_cache.scala 22:26]
  reg  valid_1_92; // @[i_cache.scala 22:26]
  reg  valid_1_93; // @[i_cache.scala 22:26]
  reg  valid_1_94; // @[i_cache.scala 22:26]
  reg  valid_1_95; // @[i_cache.scala 22:26]
  reg  valid_1_96; // @[i_cache.scala 22:26]
  reg  valid_1_97; // @[i_cache.scala 22:26]
  reg  valid_1_98; // @[i_cache.scala 22:26]
  reg  valid_1_99; // @[i_cache.scala 22:26]
  reg  valid_1_100; // @[i_cache.scala 22:26]
  reg  valid_1_101; // @[i_cache.scala 22:26]
  reg  valid_1_102; // @[i_cache.scala 22:26]
  reg  valid_1_103; // @[i_cache.scala 22:26]
  reg  valid_1_104; // @[i_cache.scala 22:26]
  reg  valid_1_105; // @[i_cache.scala 22:26]
  reg  valid_1_106; // @[i_cache.scala 22:26]
  reg  valid_1_107; // @[i_cache.scala 22:26]
  reg  valid_1_108; // @[i_cache.scala 22:26]
  reg  valid_1_109; // @[i_cache.scala 22:26]
  reg  valid_1_110; // @[i_cache.scala 22:26]
  reg  valid_1_111; // @[i_cache.scala 22:26]
  reg  valid_1_112; // @[i_cache.scala 22:26]
  reg  valid_1_113; // @[i_cache.scala 22:26]
  reg  valid_1_114; // @[i_cache.scala 22:26]
  reg  valid_1_115; // @[i_cache.scala 22:26]
  reg  valid_1_116; // @[i_cache.scala 22:26]
  reg  valid_1_117; // @[i_cache.scala 22:26]
  reg  valid_1_118; // @[i_cache.scala 22:26]
  reg  valid_1_119; // @[i_cache.scala 22:26]
  reg  valid_1_120; // @[i_cache.scala 22:26]
  reg  valid_1_121; // @[i_cache.scala 22:26]
  reg  valid_1_122; // @[i_cache.scala 22:26]
  reg  valid_1_123; // @[i_cache.scala 22:26]
  reg  valid_1_124; // @[i_cache.scala 22:26]
  reg  valid_1_125; // @[i_cache.scala 22:26]
  reg  valid_1_126; // @[i_cache.scala 22:26]
  reg  valid_1_127; // @[i_cache.scala 22:26]
  reg  way0_hit; // @[i_cache.scala 23:27]
  reg  way1_hit; // @[i_cache.scala 24:27]
  reg [1:0] unuse_way; // @[i_cache.scala 26:28]
  reg [63:0] receive_data; // @[i_cache.scala 27:31]
  reg  quene; // @[i_cache.scala 28:24]
  wire [6:0] index = io_from_ifu_araddr[6:0]; // @[i_cache.scala 31:35]
  wire [24:0] tag = io_from_ifu_araddr[31:7]; // @[i_cache.scala 32:33]
  wire [31:0] _GEN_1 = 7'h1 == index ? tag_0_1 : tag_0_0; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_2 = 7'h2 == index ? tag_0_2 : _GEN_1; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_3 = 7'h3 == index ? tag_0_3 : _GEN_2; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_4 = 7'h4 == index ? tag_0_4 : _GEN_3; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_5 = 7'h5 == index ? tag_0_5 : _GEN_4; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_6 = 7'h6 == index ? tag_0_6 : _GEN_5; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_7 = 7'h7 == index ? tag_0_7 : _GEN_6; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_8 = 7'h8 == index ? tag_0_8 : _GEN_7; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_9 = 7'h9 == index ? tag_0_9 : _GEN_8; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_10 = 7'ha == index ? tag_0_10 : _GEN_9; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_11 = 7'hb == index ? tag_0_11 : _GEN_10; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_12 = 7'hc == index ? tag_0_12 : _GEN_11; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_13 = 7'hd == index ? tag_0_13 : _GEN_12; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_14 = 7'he == index ? tag_0_14 : _GEN_13; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_15 = 7'hf == index ? tag_0_15 : _GEN_14; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_16 = 7'h10 == index ? tag_0_16 : _GEN_15; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_17 = 7'h11 == index ? tag_0_17 : _GEN_16; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_18 = 7'h12 == index ? tag_0_18 : _GEN_17; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_19 = 7'h13 == index ? tag_0_19 : _GEN_18; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_20 = 7'h14 == index ? tag_0_20 : _GEN_19; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_21 = 7'h15 == index ? tag_0_21 : _GEN_20; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_22 = 7'h16 == index ? tag_0_22 : _GEN_21; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_23 = 7'h17 == index ? tag_0_23 : _GEN_22; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_24 = 7'h18 == index ? tag_0_24 : _GEN_23; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_25 = 7'h19 == index ? tag_0_25 : _GEN_24; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_26 = 7'h1a == index ? tag_0_26 : _GEN_25; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_27 = 7'h1b == index ? tag_0_27 : _GEN_26; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_28 = 7'h1c == index ? tag_0_28 : _GEN_27; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_29 = 7'h1d == index ? tag_0_29 : _GEN_28; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_30 = 7'h1e == index ? tag_0_30 : _GEN_29; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_31 = 7'h1f == index ? tag_0_31 : _GEN_30; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_32 = 7'h20 == index ? tag_0_32 : _GEN_31; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_33 = 7'h21 == index ? tag_0_33 : _GEN_32; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_34 = 7'h22 == index ? tag_0_34 : _GEN_33; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_35 = 7'h23 == index ? tag_0_35 : _GEN_34; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_36 = 7'h24 == index ? tag_0_36 : _GEN_35; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_37 = 7'h25 == index ? tag_0_37 : _GEN_36; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_38 = 7'h26 == index ? tag_0_38 : _GEN_37; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_39 = 7'h27 == index ? tag_0_39 : _GEN_38; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_40 = 7'h28 == index ? tag_0_40 : _GEN_39; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_41 = 7'h29 == index ? tag_0_41 : _GEN_40; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_42 = 7'h2a == index ? tag_0_42 : _GEN_41; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_43 = 7'h2b == index ? tag_0_43 : _GEN_42; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_44 = 7'h2c == index ? tag_0_44 : _GEN_43; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_45 = 7'h2d == index ? tag_0_45 : _GEN_44; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_46 = 7'h2e == index ? tag_0_46 : _GEN_45; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_47 = 7'h2f == index ? tag_0_47 : _GEN_46; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_48 = 7'h30 == index ? tag_0_48 : _GEN_47; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_49 = 7'h31 == index ? tag_0_49 : _GEN_48; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_50 = 7'h32 == index ? tag_0_50 : _GEN_49; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_51 = 7'h33 == index ? tag_0_51 : _GEN_50; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_52 = 7'h34 == index ? tag_0_52 : _GEN_51; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_53 = 7'h35 == index ? tag_0_53 : _GEN_52; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_54 = 7'h36 == index ? tag_0_54 : _GEN_53; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_55 = 7'h37 == index ? tag_0_55 : _GEN_54; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_56 = 7'h38 == index ? tag_0_56 : _GEN_55; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_57 = 7'h39 == index ? tag_0_57 : _GEN_56; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_58 = 7'h3a == index ? tag_0_58 : _GEN_57; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_59 = 7'h3b == index ? tag_0_59 : _GEN_58; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_60 = 7'h3c == index ? tag_0_60 : _GEN_59; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_61 = 7'h3d == index ? tag_0_61 : _GEN_60; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_62 = 7'h3e == index ? tag_0_62 : _GEN_61; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_63 = 7'h3f == index ? tag_0_63 : _GEN_62; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_64 = 7'h40 == index ? tag_0_64 : _GEN_63; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_65 = 7'h41 == index ? tag_0_65 : _GEN_64; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_66 = 7'h42 == index ? tag_0_66 : _GEN_65; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_67 = 7'h43 == index ? tag_0_67 : _GEN_66; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_68 = 7'h44 == index ? tag_0_68 : _GEN_67; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_69 = 7'h45 == index ? tag_0_69 : _GEN_68; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_70 = 7'h46 == index ? tag_0_70 : _GEN_69; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_71 = 7'h47 == index ? tag_0_71 : _GEN_70; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_72 = 7'h48 == index ? tag_0_72 : _GEN_71; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_73 = 7'h49 == index ? tag_0_73 : _GEN_72; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_74 = 7'h4a == index ? tag_0_74 : _GEN_73; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_75 = 7'h4b == index ? tag_0_75 : _GEN_74; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_76 = 7'h4c == index ? tag_0_76 : _GEN_75; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_77 = 7'h4d == index ? tag_0_77 : _GEN_76; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_78 = 7'h4e == index ? tag_0_78 : _GEN_77; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_79 = 7'h4f == index ? tag_0_79 : _GEN_78; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_80 = 7'h50 == index ? tag_0_80 : _GEN_79; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_81 = 7'h51 == index ? tag_0_81 : _GEN_80; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_82 = 7'h52 == index ? tag_0_82 : _GEN_81; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_83 = 7'h53 == index ? tag_0_83 : _GEN_82; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_84 = 7'h54 == index ? tag_0_84 : _GEN_83; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_85 = 7'h55 == index ? tag_0_85 : _GEN_84; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_86 = 7'h56 == index ? tag_0_86 : _GEN_85; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_87 = 7'h57 == index ? tag_0_87 : _GEN_86; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_88 = 7'h58 == index ? tag_0_88 : _GEN_87; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_89 = 7'h59 == index ? tag_0_89 : _GEN_88; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_90 = 7'h5a == index ? tag_0_90 : _GEN_89; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_91 = 7'h5b == index ? tag_0_91 : _GEN_90; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_92 = 7'h5c == index ? tag_0_92 : _GEN_91; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_93 = 7'h5d == index ? tag_0_93 : _GEN_92; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_94 = 7'h5e == index ? tag_0_94 : _GEN_93; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_95 = 7'h5f == index ? tag_0_95 : _GEN_94; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_96 = 7'h60 == index ? tag_0_96 : _GEN_95; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_97 = 7'h61 == index ? tag_0_97 : _GEN_96; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_98 = 7'h62 == index ? tag_0_98 : _GEN_97; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_99 = 7'h63 == index ? tag_0_99 : _GEN_98; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_100 = 7'h64 == index ? tag_0_100 : _GEN_99; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_101 = 7'h65 == index ? tag_0_101 : _GEN_100; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_102 = 7'h66 == index ? tag_0_102 : _GEN_101; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_103 = 7'h67 == index ? tag_0_103 : _GEN_102; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_104 = 7'h68 == index ? tag_0_104 : _GEN_103; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_105 = 7'h69 == index ? tag_0_105 : _GEN_104; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_106 = 7'h6a == index ? tag_0_106 : _GEN_105; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_107 = 7'h6b == index ? tag_0_107 : _GEN_106; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_108 = 7'h6c == index ? tag_0_108 : _GEN_107; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_109 = 7'h6d == index ? tag_0_109 : _GEN_108; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_110 = 7'h6e == index ? tag_0_110 : _GEN_109; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_111 = 7'h6f == index ? tag_0_111 : _GEN_110; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_112 = 7'h70 == index ? tag_0_112 : _GEN_111; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_113 = 7'h71 == index ? tag_0_113 : _GEN_112; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_114 = 7'h72 == index ? tag_0_114 : _GEN_113; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_115 = 7'h73 == index ? tag_0_115 : _GEN_114; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_116 = 7'h74 == index ? tag_0_116 : _GEN_115; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_117 = 7'h75 == index ? tag_0_117 : _GEN_116; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_118 = 7'h76 == index ? tag_0_118 : _GEN_117; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_119 = 7'h77 == index ? tag_0_119 : _GEN_118; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_120 = 7'h78 == index ? tag_0_120 : _GEN_119; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_121 = 7'h79 == index ? tag_0_121 : _GEN_120; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_122 = 7'h7a == index ? tag_0_122 : _GEN_121; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_123 = 7'h7b == index ? tag_0_123 : _GEN_122; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_124 = 7'h7c == index ? tag_0_124 : _GEN_123; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_125 = 7'h7d == index ? tag_0_125 : _GEN_124; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_126 = 7'h7e == index ? tag_0_126 : _GEN_125; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_127 = 7'h7f == index ? tag_0_127 : _GEN_126; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_7706 = {{7'd0}, tag}; // @[i_cache.scala 34:24]
  wire  _GEN_129 = 7'h1 == index ? valid_0_1 : valid_0_0; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_130 = 7'h2 == index ? valid_0_2 : _GEN_129; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_131 = 7'h3 == index ? valid_0_3 : _GEN_130; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_132 = 7'h4 == index ? valid_0_4 : _GEN_131; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_133 = 7'h5 == index ? valid_0_5 : _GEN_132; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_134 = 7'h6 == index ? valid_0_6 : _GEN_133; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_135 = 7'h7 == index ? valid_0_7 : _GEN_134; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_136 = 7'h8 == index ? valid_0_8 : _GEN_135; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_137 = 7'h9 == index ? valid_0_9 : _GEN_136; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_138 = 7'ha == index ? valid_0_10 : _GEN_137; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_139 = 7'hb == index ? valid_0_11 : _GEN_138; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_140 = 7'hc == index ? valid_0_12 : _GEN_139; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_141 = 7'hd == index ? valid_0_13 : _GEN_140; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_142 = 7'he == index ? valid_0_14 : _GEN_141; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_143 = 7'hf == index ? valid_0_15 : _GEN_142; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_144 = 7'h10 == index ? valid_0_16 : _GEN_143; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_145 = 7'h11 == index ? valid_0_17 : _GEN_144; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_146 = 7'h12 == index ? valid_0_18 : _GEN_145; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_147 = 7'h13 == index ? valid_0_19 : _GEN_146; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_148 = 7'h14 == index ? valid_0_20 : _GEN_147; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_149 = 7'h15 == index ? valid_0_21 : _GEN_148; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_150 = 7'h16 == index ? valid_0_22 : _GEN_149; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_151 = 7'h17 == index ? valid_0_23 : _GEN_150; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_152 = 7'h18 == index ? valid_0_24 : _GEN_151; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_153 = 7'h19 == index ? valid_0_25 : _GEN_152; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_154 = 7'h1a == index ? valid_0_26 : _GEN_153; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_155 = 7'h1b == index ? valid_0_27 : _GEN_154; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_156 = 7'h1c == index ? valid_0_28 : _GEN_155; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_157 = 7'h1d == index ? valid_0_29 : _GEN_156; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_158 = 7'h1e == index ? valid_0_30 : _GEN_157; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_159 = 7'h1f == index ? valid_0_31 : _GEN_158; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_160 = 7'h20 == index ? valid_0_32 : _GEN_159; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_161 = 7'h21 == index ? valid_0_33 : _GEN_160; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_162 = 7'h22 == index ? valid_0_34 : _GEN_161; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_163 = 7'h23 == index ? valid_0_35 : _GEN_162; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_164 = 7'h24 == index ? valid_0_36 : _GEN_163; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_165 = 7'h25 == index ? valid_0_37 : _GEN_164; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_166 = 7'h26 == index ? valid_0_38 : _GEN_165; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_167 = 7'h27 == index ? valid_0_39 : _GEN_166; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_168 = 7'h28 == index ? valid_0_40 : _GEN_167; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_169 = 7'h29 == index ? valid_0_41 : _GEN_168; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_170 = 7'h2a == index ? valid_0_42 : _GEN_169; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_171 = 7'h2b == index ? valid_0_43 : _GEN_170; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_172 = 7'h2c == index ? valid_0_44 : _GEN_171; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_173 = 7'h2d == index ? valid_0_45 : _GEN_172; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_174 = 7'h2e == index ? valid_0_46 : _GEN_173; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_175 = 7'h2f == index ? valid_0_47 : _GEN_174; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_176 = 7'h30 == index ? valid_0_48 : _GEN_175; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_177 = 7'h31 == index ? valid_0_49 : _GEN_176; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_178 = 7'h32 == index ? valid_0_50 : _GEN_177; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_179 = 7'h33 == index ? valid_0_51 : _GEN_178; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_180 = 7'h34 == index ? valid_0_52 : _GEN_179; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_181 = 7'h35 == index ? valid_0_53 : _GEN_180; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_182 = 7'h36 == index ? valid_0_54 : _GEN_181; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_183 = 7'h37 == index ? valid_0_55 : _GEN_182; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_184 = 7'h38 == index ? valid_0_56 : _GEN_183; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_185 = 7'h39 == index ? valid_0_57 : _GEN_184; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_186 = 7'h3a == index ? valid_0_58 : _GEN_185; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_187 = 7'h3b == index ? valid_0_59 : _GEN_186; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_188 = 7'h3c == index ? valid_0_60 : _GEN_187; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_189 = 7'h3d == index ? valid_0_61 : _GEN_188; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_190 = 7'h3e == index ? valid_0_62 : _GEN_189; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_191 = 7'h3f == index ? valid_0_63 : _GEN_190; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_192 = 7'h40 == index ? valid_0_64 : _GEN_191; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_193 = 7'h41 == index ? valid_0_65 : _GEN_192; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_194 = 7'h42 == index ? valid_0_66 : _GEN_193; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_195 = 7'h43 == index ? valid_0_67 : _GEN_194; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_196 = 7'h44 == index ? valid_0_68 : _GEN_195; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_197 = 7'h45 == index ? valid_0_69 : _GEN_196; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_198 = 7'h46 == index ? valid_0_70 : _GEN_197; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_199 = 7'h47 == index ? valid_0_71 : _GEN_198; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_200 = 7'h48 == index ? valid_0_72 : _GEN_199; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_201 = 7'h49 == index ? valid_0_73 : _GEN_200; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_202 = 7'h4a == index ? valid_0_74 : _GEN_201; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_203 = 7'h4b == index ? valid_0_75 : _GEN_202; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_204 = 7'h4c == index ? valid_0_76 : _GEN_203; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_205 = 7'h4d == index ? valid_0_77 : _GEN_204; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_206 = 7'h4e == index ? valid_0_78 : _GEN_205; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_207 = 7'h4f == index ? valid_0_79 : _GEN_206; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_208 = 7'h50 == index ? valid_0_80 : _GEN_207; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_209 = 7'h51 == index ? valid_0_81 : _GEN_208; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_210 = 7'h52 == index ? valid_0_82 : _GEN_209; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_211 = 7'h53 == index ? valid_0_83 : _GEN_210; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_212 = 7'h54 == index ? valid_0_84 : _GEN_211; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_213 = 7'h55 == index ? valid_0_85 : _GEN_212; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_214 = 7'h56 == index ? valid_0_86 : _GEN_213; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_215 = 7'h57 == index ? valid_0_87 : _GEN_214; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_216 = 7'h58 == index ? valid_0_88 : _GEN_215; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_217 = 7'h59 == index ? valid_0_89 : _GEN_216; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_218 = 7'h5a == index ? valid_0_90 : _GEN_217; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_219 = 7'h5b == index ? valid_0_91 : _GEN_218; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_220 = 7'h5c == index ? valid_0_92 : _GEN_219; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_221 = 7'h5d == index ? valid_0_93 : _GEN_220; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_222 = 7'h5e == index ? valid_0_94 : _GEN_221; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_223 = 7'h5f == index ? valid_0_95 : _GEN_222; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_224 = 7'h60 == index ? valid_0_96 : _GEN_223; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_225 = 7'h61 == index ? valid_0_97 : _GEN_224; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_226 = 7'h62 == index ? valid_0_98 : _GEN_225; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_227 = 7'h63 == index ? valid_0_99 : _GEN_226; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_228 = 7'h64 == index ? valid_0_100 : _GEN_227; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_229 = 7'h65 == index ? valid_0_101 : _GEN_228; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_230 = 7'h66 == index ? valid_0_102 : _GEN_229; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_231 = 7'h67 == index ? valid_0_103 : _GEN_230; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_232 = 7'h68 == index ? valid_0_104 : _GEN_231; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_233 = 7'h69 == index ? valid_0_105 : _GEN_232; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_234 = 7'h6a == index ? valid_0_106 : _GEN_233; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_235 = 7'h6b == index ? valid_0_107 : _GEN_234; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_236 = 7'h6c == index ? valid_0_108 : _GEN_235; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_237 = 7'h6d == index ? valid_0_109 : _GEN_236; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_238 = 7'h6e == index ? valid_0_110 : _GEN_237; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_239 = 7'h6f == index ? valid_0_111 : _GEN_238; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_240 = 7'h70 == index ? valid_0_112 : _GEN_239; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_241 = 7'h71 == index ? valid_0_113 : _GEN_240; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_242 = 7'h72 == index ? valid_0_114 : _GEN_241; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_243 = 7'h73 == index ? valid_0_115 : _GEN_242; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_244 = 7'h74 == index ? valid_0_116 : _GEN_243; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_245 = 7'h75 == index ? valid_0_117 : _GEN_244; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_246 = 7'h76 == index ? valid_0_118 : _GEN_245; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_247 = 7'h77 == index ? valid_0_119 : _GEN_246; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_248 = 7'h78 == index ? valid_0_120 : _GEN_247; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_249 = 7'h79 == index ? valid_0_121 : _GEN_248; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_250 = 7'h7a == index ? valid_0_122 : _GEN_249; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_251 = 7'h7b == index ? valid_0_123 : _GEN_250; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_252 = 7'h7c == index ? valid_0_124 : _GEN_251; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_253 = 7'h7d == index ? valid_0_125 : _GEN_252; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_254 = 7'h7e == index ? valid_0_126 : _GEN_253; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_255 = 7'h7f == index ? valid_0_127 : _GEN_254; // @[i_cache.scala 34:{50,50}]
  wire  _T_2 = _GEN_127 == _GEN_7706 & _GEN_255; // @[i_cache.scala 34:33]
  wire [31:0] _GEN_258 = 7'h1 == index ? tag_1_1 : tag_1_0; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_259 = 7'h2 == index ? tag_1_2 : _GEN_258; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_260 = 7'h3 == index ? tag_1_3 : _GEN_259; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_261 = 7'h4 == index ? tag_1_4 : _GEN_260; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_262 = 7'h5 == index ? tag_1_5 : _GEN_261; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_263 = 7'h6 == index ? tag_1_6 : _GEN_262; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_264 = 7'h7 == index ? tag_1_7 : _GEN_263; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_265 = 7'h8 == index ? tag_1_8 : _GEN_264; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_266 = 7'h9 == index ? tag_1_9 : _GEN_265; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_267 = 7'ha == index ? tag_1_10 : _GEN_266; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_268 = 7'hb == index ? tag_1_11 : _GEN_267; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_269 = 7'hc == index ? tag_1_12 : _GEN_268; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_270 = 7'hd == index ? tag_1_13 : _GEN_269; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_271 = 7'he == index ? tag_1_14 : _GEN_270; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_272 = 7'hf == index ? tag_1_15 : _GEN_271; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_273 = 7'h10 == index ? tag_1_16 : _GEN_272; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_274 = 7'h11 == index ? tag_1_17 : _GEN_273; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_275 = 7'h12 == index ? tag_1_18 : _GEN_274; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_276 = 7'h13 == index ? tag_1_19 : _GEN_275; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_277 = 7'h14 == index ? tag_1_20 : _GEN_276; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_278 = 7'h15 == index ? tag_1_21 : _GEN_277; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_279 = 7'h16 == index ? tag_1_22 : _GEN_278; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_280 = 7'h17 == index ? tag_1_23 : _GEN_279; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_281 = 7'h18 == index ? tag_1_24 : _GEN_280; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_282 = 7'h19 == index ? tag_1_25 : _GEN_281; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_283 = 7'h1a == index ? tag_1_26 : _GEN_282; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_284 = 7'h1b == index ? tag_1_27 : _GEN_283; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_285 = 7'h1c == index ? tag_1_28 : _GEN_284; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_286 = 7'h1d == index ? tag_1_29 : _GEN_285; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_287 = 7'h1e == index ? tag_1_30 : _GEN_286; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_288 = 7'h1f == index ? tag_1_31 : _GEN_287; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_289 = 7'h20 == index ? tag_1_32 : _GEN_288; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_290 = 7'h21 == index ? tag_1_33 : _GEN_289; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_291 = 7'h22 == index ? tag_1_34 : _GEN_290; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_292 = 7'h23 == index ? tag_1_35 : _GEN_291; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_293 = 7'h24 == index ? tag_1_36 : _GEN_292; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_294 = 7'h25 == index ? tag_1_37 : _GEN_293; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_295 = 7'h26 == index ? tag_1_38 : _GEN_294; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_296 = 7'h27 == index ? tag_1_39 : _GEN_295; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_297 = 7'h28 == index ? tag_1_40 : _GEN_296; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_298 = 7'h29 == index ? tag_1_41 : _GEN_297; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_299 = 7'h2a == index ? tag_1_42 : _GEN_298; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_300 = 7'h2b == index ? tag_1_43 : _GEN_299; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_301 = 7'h2c == index ? tag_1_44 : _GEN_300; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_302 = 7'h2d == index ? tag_1_45 : _GEN_301; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_303 = 7'h2e == index ? tag_1_46 : _GEN_302; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_304 = 7'h2f == index ? tag_1_47 : _GEN_303; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_305 = 7'h30 == index ? tag_1_48 : _GEN_304; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_306 = 7'h31 == index ? tag_1_49 : _GEN_305; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_307 = 7'h32 == index ? tag_1_50 : _GEN_306; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_308 = 7'h33 == index ? tag_1_51 : _GEN_307; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_309 = 7'h34 == index ? tag_1_52 : _GEN_308; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_310 = 7'h35 == index ? tag_1_53 : _GEN_309; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_311 = 7'h36 == index ? tag_1_54 : _GEN_310; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_312 = 7'h37 == index ? tag_1_55 : _GEN_311; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_313 = 7'h38 == index ? tag_1_56 : _GEN_312; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_314 = 7'h39 == index ? tag_1_57 : _GEN_313; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_315 = 7'h3a == index ? tag_1_58 : _GEN_314; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_316 = 7'h3b == index ? tag_1_59 : _GEN_315; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_317 = 7'h3c == index ? tag_1_60 : _GEN_316; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_318 = 7'h3d == index ? tag_1_61 : _GEN_317; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_319 = 7'h3e == index ? tag_1_62 : _GEN_318; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_320 = 7'h3f == index ? tag_1_63 : _GEN_319; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_321 = 7'h40 == index ? tag_1_64 : _GEN_320; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_322 = 7'h41 == index ? tag_1_65 : _GEN_321; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_323 = 7'h42 == index ? tag_1_66 : _GEN_322; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_324 = 7'h43 == index ? tag_1_67 : _GEN_323; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_325 = 7'h44 == index ? tag_1_68 : _GEN_324; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_326 = 7'h45 == index ? tag_1_69 : _GEN_325; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_327 = 7'h46 == index ? tag_1_70 : _GEN_326; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_328 = 7'h47 == index ? tag_1_71 : _GEN_327; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_329 = 7'h48 == index ? tag_1_72 : _GEN_328; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_330 = 7'h49 == index ? tag_1_73 : _GEN_329; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_331 = 7'h4a == index ? tag_1_74 : _GEN_330; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_332 = 7'h4b == index ? tag_1_75 : _GEN_331; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_333 = 7'h4c == index ? tag_1_76 : _GEN_332; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_334 = 7'h4d == index ? tag_1_77 : _GEN_333; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_335 = 7'h4e == index ? tag_1_78 : _GEN_334; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_336 = 7'h4f == index ? tag_1_79 : _GEN_335; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_337 = 7'h50 == index ? tag_1_80 : _GEN_336; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_338 = 7'h51 == index ? tag_1_81 : _GEN_337; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_339 = 7'h52 == index ? tag_1_82 : _GEN_338; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_340 = 7'h53 == index ? tag_1_83 : _GEN_339; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_341 = 7'h54 == index ? tag_1_84 : _GEN_340; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_342 = 7'h55 == index ? tag_1_85 : _GEN_341; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_343 = 7'h56 == index ? tag_1_86 : _GEN_342; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_344 = 7'h57 == index ? tag_1_87 : _GEN_343; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_345 = 7'h58 == index ? tag_1_88 : _GEN_344; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_346 = 7'h59 == index ? tag_1_89 : _GEN_345; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_347 = 7'h5a == index ? tag_1_90 : _GEN_346; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_348 = 7'h5b == index ? tag_1_91 : _GEN_347; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_349 = 7'h5c == index ? tag_1_92 : _GEN_348; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_350 = 7'h5d == index ? tag_1_93 : _GEN_349; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_351 = 7'h5e == index ? tag_1_94 : _GEN_350; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_352 = 7'h5f == index ? tag_1_95 : _GEN_351; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_353 = 7'h60 == index ? tag_1_96 : _GEN_352; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_354 = 7'h61 == index ? tag_1_97 : _GEN_353; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_355 = 7'h62 == index ? tag_1_98 : _GEN_354; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_356 = 7'h63 == index ? tag_1_99 : _GEN_355; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_357 = 7'h64 == index ? tag_1_100 : _GEN_356; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_358 = 7'h65 == index ? tag_1_101 : _GEN_357; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_359 = 7'h66 == index ? tag_1_102 : _GEN_358; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_360 = 7'h67 == index ? tag_1_103 : _GEN_359; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_361 = 7'h68 == index ? tag_1_104 : _GEN_360; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_362 = 7'h69 == index ? tag_1_105 : _GEN_361; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_363 = 7'h6a == index ? tag_1_106 : _GEN_362; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_364 = 7'h6b == index ? tag_1_107 : _GEN_363; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_365 = 7'h6c == index ? tag_1_108 : _GEN_364; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_366 = 7'h6d == index ? tag_1_109 : _GEN_365; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_367 = 7'h6e == index ? tag_1_110 : _GEN_366; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_368 = 7'h6f == index ? tag_1_111 : _GEN_367; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_369 = 7'h70 == index ? tag_1_112 : _GEN_368; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_370 = 7'h71 == index ? tag_1_113 : _GEN_369; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_371 = 7'h72 == index ? tag_1_114 : _GEN_370; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_372 = 7'h73 == index ? tag_1_115 : _GEN_371; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_373 = 7'h74 == index ? tag_1_116 : _GEN_372; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_374 = 7'h75 == index ? tag_1_117 : _GEN_373; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_375 = 7'h76 == index ? tag_1_118 : _GEN_374; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_376 = 7'h77 == index ? tag_1_119 : _GEN_375; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_377 = 7'h78 == index ? tag_1_120 : _GEN_376; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_378 = 7'h79 == index ? tag_1_121 : _GEN_377; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_379 = 7'h7a == index ? tag_1_122 : _GEN_378; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_380 = 7'h7b == index ? tag_1_123 : _GEN_379; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_381 = 7'h7c == index ? tag_1_124 : _GEN_380; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_382 = 7'h7d == index ? tag_1_125 : _GEN_381; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_383 = 7'h7e == index ? tag_1_126 : _GEN_382; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_384 = 7'h7f == index ? tag_1_127 : _GEN_383; // @[i_cache.scala 39:{24,24}]
  wire  _GEN_386 = 7'h1 == index ? valid_1_1 : valid_1_0; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_387 = 7'h2 == index ? valid_1_2 : _GEN_386; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_388 = 7'h3 == index ? valid_1_3 : _GEN_387; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_389 = 7'h4 == index ? valid_1_4 : _GEN_388; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_390 = 7'h5 == index ? valid_1_5 : _GEN_389; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_391 = 7'h6 == index ? valid_1_6 : _GEN_390; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_392 = 7'h7 == index ? valid_1_7 : _GEN_391; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_393 = 7'h8 == index ? valid_1_8 : _GEN_392; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_394 = 7'h9 == index ? valid_1_9 : _GEN_393; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_395 = 7'ha == index ? valid_1_10 : _GEN_394; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_396 = 7'hb == index ? valid_1_11 : _GEN_395; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_397 = 7'hc == index ? valid_1_12 : _GEN_396; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_398 = 7'hd == index ? valid_1_13 : _GEN_397; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_399 = 7'he == index ? valid_1_14 : _GEN_398; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_400 = 7'hf == index ? valid_1_15 : _GEN_399; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_401 = 7'h10 == index ? valid_1_16 : _GEN_400; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_402 = 7'h11 == index ? valid_1_17 : _GEN_401; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_403 = 7'h12 == index ? valid_1_18 : _GEN_402; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_404 = 7'h13 == index ? valid_1_19 : _GEN_403; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_405 = 7'h14 == index ? valid_1_20 : _GEN_404; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_406 = 7'h15 == index ? valid_1_21 : _GEN_405; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_407 = 7'h16 == index ? valid_1_22 : _GEN_406; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_408 = 7'h17 == index ? valid_1_23 : _GEN_407; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_409 = 7'h18 == index ? valid_1_24 : _GEN_408; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_410 = 7'h19 == index ? valid_1_25 : _GEN_409; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_411 = 7'h1a == index ? valid_1_26 : _GEN_410; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_412 = 7'h1b == index ? valid_1_27 : _GEN_411; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_413 = 7'h1c == index ? valid_1_28 : _GEN_412; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_414 = 7'h1d == index ? valid_1_29 : _GEN_413; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_415 = 7'h1e == index ? valid_1_30 : _GEN_414; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_416 = 7'h1f == index ? valid_1_31 : _GEN_415; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_417 = 7'h20 == index ? valid_1_32 : _GEN_416; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_418 = 7'h21 == index ? valid_1_33 : _GEN_417; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_419 = 7'h22 == index ? valid_1_34 : _GEN_418; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_420 = 7'h23 == index ? valid_1_35 : _GEN_419; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_421 = 7'h24 == index ? valid_1_36 : _GEN_420; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_422 = 7'h25 == index ? valid_1_37 : _GEN_421; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_423 = 7'h26 == index ? valid_1_38 : _GEN_422; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_424 = 7'h27 == index ? valid_1_39 : _GEN_423; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_425 = 7'h28 == index ? valid_1_40 : _GEN_424; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_426 = 7'h29 == index ? valid_1_41 : _GEN_425; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_427 = 7'h2a == index ? valid_1_42 : _GEN_426; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_428 = 7'h2b == index ? valid_1_43 : _GEN_427; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_429 = 7'h2c == index ? valid_1_44 : _GEN_428; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_430 = 7'h2d == index ? valid_1_45 : _GEN_429; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_431 = 7'h2e == index ? valid_1_46 : _GEN_430; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_432 = 7'h2f == index ? valid_1_47 : _GEN_431; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_433 = 7'h30 == index ? valid_1_48 : _GEN_432; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_434 = 7'h31 == index ? valid_1_49 : _GEN_433; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_435 = 7'h32 == index ? valid_1_50 : _GEN_434; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_436 = 7'h33 == index ? valid_1_51 : _GEN_435; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_437 = 7'h34 == index ? valid_1_52 : _GEN_436; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_438 = 7'h35 == index ? valid_1_53 : _GEN_437; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_439 = 7'h36 == index ? valid_1_54 : _GEN_438; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_440 = 7'h37 == index ? valid_1_55 : _GEN_439; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_441 = 7'h38 == index ? valid_1_56 : _GEN_440; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_442 = 7'h39 == index ? valid_1_57 : _GEN_441; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_443 = 7'h3a == index ? valid_1_58 : _GEN_442; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_444 = 7'h3b == index ? valid_1_59 : _GEN_443; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_445 = 7'h3c == index ? valid_1_60 : _GEN_444; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_446 = 7'h3d == index ? valid_1_61 : _GEN_445; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_447 = 7'h3e == index ? valid_1_62 : _GEN_446; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_448 = 7'h3f == index ? valid_1_63 : _GEN_447; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_449 = 7'h40 == index ? valid_1_64 : _GEN_448; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_450 = 7'h41 == index ? valid_1_65 : _GEN_449; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_451 = 7'h42 == index ? valid_1_66 : _GEN_450; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_452 = 7'h43 == index ? valid_1_67 : _GEN_451; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_453 = 7'h44 == index ? valid_1_68 : _GEN_452; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_454 = 7'h45 == index ? valid_1_69 : _GEN_453; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_455 = 7'h46 == index ? valid_1_70 : _GEN_454; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_456 = 7'h47 == index ? valid_1_71 : _GEN_455; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_457 = 7'h48 == index ? valid_1_72 : _GEN_456; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_458 = 7'h49 == index ? valid_1_73 : _GEN_457; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_459 = 7'h4a == index ? valid_1_74 : _GEN_458; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_460 = 7'h4b == index ? valid_1_75 : _GEN_459; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_461 = 7'h4c == index ? valid_1_76 : _GEN_460; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_462 = 7'h4d == index ? valid_1_77 : _GEN_461; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_463 = 7'h4e == index ? valid_1_78 : _GEN_462; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_464 = 7'h4f == index ? valid_1_79 : _GEN_463; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_465 = 7'h50 == index ? valid_1_80 : _GEN_464; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_466 = 7'h51 == index ? valid_1_81 : _GEN_465; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_467 = 7'h52 == index ? valid_1_82 : _GEN_466; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_468 = 7'h53 == index ? valid_1_83 : _GEN_467; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_469 = 7'h54 == index ? valid_1_84 : _GEN_468; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_470 = 7'h55 == index ? valid_1_85 : _GEN_469; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_471 = 7'h56 == index ? valid_1_86 : _GEN_470; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_472 = 7'h57 == index ? valid_1_87 : _GEN_471; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_473 = 7'h58 == index ? valid_1_88 : _GEN_472; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_474 = 7'h59 == index ? valid_1_89 : _GEN_473; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_475 = 7'h5a == index ? valid_1_90 : _GEN_474; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_476 = 7'h5b == index ? valid_1_91 : _GEN_475; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_477 = 7'h5c == index ? valid_1_92 : _GEN_476; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_478 = 7'h5d == index ? valid_1_93 : _GEN_477; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_479 = 7'h5e == index ? valid_1_94 : _GEN_478; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_480 = 7'h5f == index ? valid_1_95 : _GEN_479; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_481 = 7'h60 == index ? valid_1_96 : _GEN_480; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_482 = 7'h61 == index ? valid_1_97 : _GEN_481; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_483 = 7'h62 == index ? valid_1_98 : _GEN_482; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_484 = 7'h63 == index ? valid_1_99 : _GEN_483; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_485 = 7'h64 == index ? valid_1_100 : _GEN_484; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_486 = 7'h65 == index ? valid_1_101 : _GEN_485; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_487 = 7'h66 == index ? valid_1_102 : _GEN_486; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_488 = 7'h67 == index ? valid_1_103 : _GEN_487; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_489 = 7'h68 == index ? valid_1_104 : _GEN_488; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_490 = 7'h69 == index ? valid_1_105 : _GEN_489; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_491 = 7'h6a == index ? valid_1_106 : _GEN_490; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_492 = 7'h6b == index ? valid_1_107 : _GEN_491; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_493 = 7'h6c == index ? valid_1_108 : _GEN_492; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_494 = 7'h6d == index ? valid_1_109 : _GEN_493; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_495 = 7'h6e == index ? valid_1_110 : _GEN_494; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_496 = 7'h6f == index ? valid_1_111 : _GEN_495; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_497 = 7'h70 == index ? valid_1_112 : _GEN_496; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_498 = 7'h71 == index ? valid_1_113 : _GEN_497; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_499 = 7'h72 == index ? valid_1_114 : _GEN_498; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_500 = 7'h73 == index ? valid_1_115 : _GEN_499; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_501 = 7'h74 == index ? valid_1_116 : _GEN_500; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_502 = 7'h75 == index ? valid_1_117 : _GEN_501; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_503 = 7'h76 == index ? valid_1_118 : _GEN_502; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_504 = 7'h77 == index ? valid_1_119 : _GEN_503; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_505 = 7'h78 == index ? valid_1_120 : _GEN_504; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_506 = 7'h79 == index ? valid_1_121 : _GEN_505; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_507 = 7'h7a == index ? valid_1_122 : _GEN_506; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_508 = 7'h7b == index ? valid_1_123 : _GEN_507; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_509 = 7'h7c == index ? valid_1_124 : _GEN_508; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_510 = 7'h7d == index ? valid_1_125 : _GEN_509; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_511 = 7'h7e == index ? valid_1_126 : _GEN_510; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_512 = 7'h7f == index ? valid_1_127 : _GEN_511; // @[i_cache.scala 39:{50,50}]
  wire  _T_5 = _GEN_384 == _GEN_7706 & _GEN_512; // @[i_cache.scala 39:33]
  reg [2:0] state; // @[i_cache.scala 53:24]
  wire [2:0] _GEN_517 = io_from_ifu_rready ? 3'h0 : state; // @[i_cache.scala 53:24 64:41 65:27]
  wire [2:0] _GEN_518 = way1_hit ? _GEN_517 : 3'h2; // @[i_cache.scala 68:33 73:23]
  wire [2:0] _GEN_520 = io_from_axi_rvalid ? 3'h3 : state; // @[i_cache.scala 77:37 78:23 53:24]
  wire [63:0] _GEN_521 = io_from_axi_rvalid ? io_from_axi_rdata : receive_data; // @[i_cache.scala 80:37 81:30 27:31]
  wire [63:0] _GEN_522 = 7'h0 == index ? receive_data : ram_0_0; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_523 = 7'h1 == index ? receive_data : ram_0_1; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_524 = 7'h2 == index ? receive_data : ram_0_2; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_525 = 7'h3 == index ? receive_data : ram_0_3; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_526 = 7'h4 == index ? receive_data : ram_0_4; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_527 = 7'h5 == index ? receive_data : ram_0_5; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_528 = 7'h6 == index ? receive_data : ram_0_6; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_529 = 7'h7 == index ? receive_data : ram_0_7; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_530 = 7'h8 == index ? receive_data : ram_0_8; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_531 = 7'h9 == index ? receive_data : ram_0_9; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_532 = 7'ha == index ? receive_data : ram_0_10; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_533 = 7'hb == index ? receive_data : ram_0_11; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_534 = 7'hc == index ? receive_data : ram_0_12; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_535 = 7'hd == index ? receive_data : ram_0_13; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_536 = 7'he == index ? receive_data : ram_0_14; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_537 = 7'hf == index ? receive_data : ram_0_15; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_538 = 7'h10 == index ? receive_data : ram_0_16; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_539 = 7'h11 == index ? receive_data : ram_0_17; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_540 = 7'h12 == index ? receive_data : ram_0_18; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_541 = 7'h13 == index ? receive_data : ram_0_19; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_542 = 7'h14 == index ? receive_data : ram_0_20; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_543 = 7'h15 == index ? receive_data : ram_0_21; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_544 = 7'h16 == index ? receive_data : ram_0_22; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_545 = 7'h17 == index ? receive_data : ram_0_23; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_546 = 7'h18 == index ? receive_data : ram_0_24; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_547 = 7'h19 == index ? receive_data : ram_0_25; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_548 = 7'h1a == index ? receive_data : ram_0_26; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_549 = 7'h1b == index ? receive_data : ram_0_27; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_550 = 7'h1c == index ? receive_data : ram_0_28; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_551 = 7'h1d == index ? receive_data : ram_0_29; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_552 = 7'h1e == index ? receive_data : ram_0_30; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_553 = 7'h1f == index ? receive_data : ram_0_31; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_554 = 7'h20 == index ? receive_data : ram_0_32; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_555 = 7'h21 == index ? receive_data : ram_0_33; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_556 = 7'h22 == index ? receive_data : ram_0_34; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_557 = 7'h23 == index ? receive_data : ram_0_35; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_558 = 7'h24 == index ? receive_data : ram_0_36; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_559 = 7'h25 == index ? receive_data : ram_0_37; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_560 = 7'h26 == index ? receive_data : ram_0_38; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_561 = 7'h27 == index ? receive_data : ram_0_39; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_562 = 7'h28 == index ? receive_data : ram_0_40; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_563 = 7'h29 == index ? receive_data : ram_0_41; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_564 = 7'h2a == index ? receive_data : ram_0_42; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_565 = 7'h2b == index ? receive_data : ram_0_43; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_566 = 7'h2c == index ? receive_data : ram_0_44; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_567 = 7'h2d == index ? receive_data : ram_0_45; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_568 = 7'h2e == index ? receive_data : ram_0_46; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_569 = 7'h2f == index ? receive_data : ram_0_47; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_570 = 7'h30 == index ? receive_data : ram_0_48; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_571 = 7'h31 == index ? receive_data : ram_0_49; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_572 = 7'h32 == index ? receive_data : ram_0_50; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_573 = 7'h33 == index ? receive_data : ram_0_51; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_574 = 7'h34 == index ? receive_data : ram_0_52; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_575 = 7'h35 == index ? receive_data : ram_0_53; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_576 = 7'h36 == index ? receive_data : ram_0_54; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_577 = 7'h37 == index ? receive_data : ram_0_55; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_578 = 7'h38 == index ? receive_data : ram_0_56; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_579 = 7'h39 == index ? receive_data : ram_0_57; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_580 = 7'h3a == index ? receive_data : ram_0_58; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_581 = 7'h3b == index ? receive_data : ram_0_59; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_582 = 7'h3c == index ? receive_data : ram_0_60; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_583 = 7'h3d == index ? receive_data : ram_0_61; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_584 = 7'h3e == index ? receive_data : ram_0_62; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_585 = 7'h3f == index ? receive_data : ram_0_63; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_586 = 7'h40 == index ? receive_data : ram_0_64; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_587 = 7'h41 == index ? receive_data : ram_0_65; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_588 = 7'h42 == index ? receive_data : ram_0_66; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_589 = 7'h43 == index ? receive_data : ram_0_67; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_590 = 7'h44 == index ? receive_data : ram_0_68; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_591 = 7'h45 == index ? receive_data : ram_0_69; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_592 = 7'h46 == index ? receive_data : ram_0_70; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_593 = 7'h47 == index ? receive_data : ram_0_71; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_594 = 7'h48 == index ? receive_data : ram_0_72; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_595 = 7'h49 == index ? receive_data : ram_0_73; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_596 = 7'h4a == index ? receive_data : ram_0_74; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_597 = 7'h4b == index ? receive_data : ram_0_75; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_598 = 7'h4c == index ? receive_data : ram_0_76; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_599 = 7'h4d == index ? receive_data : ram_0_77; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_600 = 7'h4e == index ? receive_data : ram_0_78; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_601 = 7'h4f == index ? receive_data : ram_0_79; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_602 = 7'h50 == index ? receive_data : ram_0_80; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_603 = 7'h51 == index ? receive_data : ram_0_81; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_604 = 7'h52 == index ? receive_data : ram_0_82; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_605 = 7'h53 == index ? receive_data : ram_0_83; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_606 = 7'h54 == index ? receive_data : ram_0_84; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_607 = 7'h55 == index ? receive_data : ram_0_85; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_608 = 7'h56 == index ? receive_data : ram_0_86; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_609 = 7'h57 == index ? receive_data : ram_0_87; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_610 = 7'h58 == index ? receive_data : ram_0_88; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_611 = 7'h59 == index ? receive_data : ram_0_89; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_612 = 7'h5a == index ? receive_data : ram_0_90; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_613 = 7'h5b == index ? receive_data : ram_0_91; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_614 = 7'h5c == index ? receive_data : ram_0_92; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_615 = 7'h5d == index ? receive_data : ram_0_93; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_616 = 7'h5e == index ? receive_data : ram_0_94; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_617 = 7'h5f == index ? receive_data : ram_0_95; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_618 = 7'h60 == index ? receive_data : ram_0_96; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_619 = 7'h61 == index ? receive_data : ram_0_97; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_620 = 7'h62 == index ? receive_data : ram_0_98; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_621 = 7'h63 == index ? receive_data : ram_0_99; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_622 = 7'h64 == index ? receive_data : ram_0_100; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_623 = 7'h65 == index ? receive_data : ram_0_101; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_624 = 7'h66 == index ? receive_data : ram_0_102; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_625 = 7'h67 == index ? receive_data : ram_0_103; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_626 = 7'h68 == index ? receive_data : ram_0_104; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_627 = 7'h69 == index ? receive_data : ram_0_105; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_628 = 7'h6a == index ? receive_data : ram_0_106; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_629 = 7'h6b == index ? receive_data : ram_0_107; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_630 = 7'h6c == index ? receive_data : ram_0_108; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_631 = 7'h6d == index ? receive_data : ram_0_109; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_632 = 7'h6e == index ? receive_data : ram_0_110; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_633 = 7'h6f == index ? receive_data : ram_0_111; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_634 = 7'h70 == index ? receive_data : ram_0_112; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_635 = 7'h71 == index ? receive_data : ram_0_113; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_636 = 7'h72 == index ? receive_data : ram_0_114; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_637 = 7'h73 == index ? receive_data : ram_0_115; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_638 = 7'h74 == index ? receive_data : ram_0_116; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_639 = 7'h75 == index ? receive_data : ram_0_117; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_640 = 7'h76 == index ? receive_data : ram_0_118; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_641 = 7'h77 == index ? receive_data : ram_0_119; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_642 = 7'h78 == index ? receive_data : ram_0_120; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_643 = 7'h79 == index ? receive_data : ram_0_121; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_644 = 7'h7a == index ? receive_data : ram_0_122; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_645 = 7'h7b == index ? receive_data : ram_0_123; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_646 = 7'h7c == index ? receive_data : ram_0_124; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_647 = 7'h7d == index ? receive_data : ram_0_125; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_648 = 7'h7e == index ? receive_data : ram_0_126; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_649 = 7'h7f == index ? receive_data : ram_0_127; // @[i_cache.scala 17:24 87:{30,30}]
  wire [31:0] _GEN_650 = 7'h0 == index ? _GEN_7706 : tag_0_0; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_651 = 7'h1 == index ? _GEN_7706 : tag_0_1; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_652 = 7'h2 == index ? _GEN_7706 : tag_0_2; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_653 = 7'h3 == index ? _GEN_7706 : tag_0_3; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_654 = 7'h4 == index ? _GEN_7706 : tag_0_4; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_655 = 7'h5 == index ? _GEN_7706 : tag_0_5; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_656 = 7'h6 == index ? _GEN_7706 : tag_0_6; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_657 = 7'h7 == index ? _GEN_7706 : tag_0_7; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_658 = 7'h8 == index ? _GEN_7706 : tag_0_8; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_659 = 7'h9 == index ? _GEN_7706 : tag_0_9; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_660 = 7'ha == index ? _GEN_7706 : tag_0_10; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_661 = 7'hb == index ? _GEN_7706 : tag_0_11; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_662 = 7'hc == index ? _GEN_7706 : tag_0_12; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_663 = 7'hd == index ? _GEN_7706 : tag_0_13; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_664 = 7'he == index ? _GEN_7706 : tag_0_14; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_665 = 7'hf == index ? _GEN_7706 : tag_0_15; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_666 = 7'h10 == index ? _GEN_7706 : tag_0_16; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_667 = 7'h11 == index ? _GEN_7706 : tag_0_17; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_668 = 7'h12 == index ? _GEN_7706 : tag_0_18; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_669 = 7'h13 == index ? _GEN_7706 : tag_0_19; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_670 = 7'h14 == index ? _GEN_7706 : tag_0_20; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_671 = 7'h15 == index ? _GEN_7706 : tag_0_21; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_672 = 7'h16 == index ? _GEN_7706 : tag_0_22; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_673 = 7'h17 == index ? _GEN_7706 : tag_0_23; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_674 = 7'h18 == index ? _GEN_7706 : tag_0_24; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_675 = 7'h19 == index ? _GEN_7706 : tag_0_25; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_676 = 7'h1a == index ? _GEN_7706 : tag_0_26; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_677 = 7'h1b == index ? _GEN_7706 : tag_0_27; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_678 = 7'h1c == index ? _GEN_7706 : tag_0_28; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_679 = 7'h1d == index ? _GEN_7706 : tag_0_29; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_680 = 7'h1e == index ? _GEN_7706 : tag_0_30; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_681 = 7'h1f == index ? _GEN_7706 : tag_0_31; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_682 = 7'h20 == index ? _GEN_7706 : tag_0_32; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_683 = 7'h21 == index ? _GEN_7706 : tag_0_33; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_684 = 7'h22 == index ? _GEN_7706 : tag_0_34; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_685 = 7'h23 == index ? _GEN_7706 : tag_0_35; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_686 = 7'h24 == index ? _GEN_7706 : tag_0_36; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_687 = 7'h25 == index ? _GEN_7706 : tag_0_37; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_688 = 7'h26 == index ? _GEN_7706 : tag_0_38; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_689 = 7'h27 == index ? _GEN_7706 : tag_0_39; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_690 = 7'h28 == index ? _GEN_7706 : tag_0_40; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_691 = 7'h29 == index ? _GEN_7706 : tag_0_41; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_692 = 7'h2a == index ? _GEN_7706 : tag_0_42; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_693 = 7'h2b == index ? _GEN_7706 : tag_0_43; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_694 = 7'h2c == index ? _GEN_7706 : tag_0_44; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_695 = 7'h2d == index ? _GEN_7706 : tag_0_45; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_696 = 7'h2e == index ? _GEN_7706 : tag_0_46; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_697 = 7'h2f == index ? _GEN_7706 : tag_0_47; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_698 = 7'h30 == index ? _GEN_7706 : tag_0_48; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_699 = 7'h31 == index ? _GEN_7706 : tag_0_49; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_700 = 7'h32 == index ? _GEN_7706 : tag_0_50; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_701 = 7'h33 == index ? _GEN_7706 : tag_0_51; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_702 = 7'h34 == index ? _GEN_7706 : tag_0_52; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_703 = 7'h35 == index ? _GEN_7706 : tag_0_53; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_704 = 7'h36 == index ? _GEN_7706 : tag_0_54; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_705 = 7'h37 == index ? _GEN_7706 : tag_0_55; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_706 = 7'h38 == index ? _GEN_7706 : tag_0_56; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_707 = 7'h39 == index ? _GEN_7706 : tag_0_57; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_708 = 7'h3a == index ? _GEN_7706 : tag_0_58; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_709 = 7'h3b == index ? _GEN_7706 : tag_0_59; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_710 = 7'h3c == index ? _GEN_7706 : tag_0_60; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_711 = 7'h3d == index ? _GEN_7706 : tag_0_61; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_712 = 7'h3e == index ? _GEN_7706 : tag_0_62; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_713 = 7'h3f == index ? _GEN_7706 : tag_0_63; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_714 = 7'h40 == index ? _GEN_7706 : tag_0_64; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_715 = 7'h41 == index ? _GEN_7706 : tag_0_65; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_716 = 7'h42 == index ? _GEN_7706 : tag_0_66; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_717 = 7'h43 == index ? _GEN_7706 : tag_0_67; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_718 = 7'h44 == index ? _GEN_7706 : tag_0_68; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_719 = 7'h45 == index ? _GEN_7706 : tag_0_69; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_720 = 7'h46 == index ? _GEN_7706 : tag_0_70; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_721 = 7'h47 == index ? _GEN_7706 : tag_0_71; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_722 = 7'h48 == index ? _GEN_7706 : tag_0_72; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_723 = 7'h49 == index ? _GEN_7706 : tag_0_73; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_724 = 7'h4a == index ? _GEN_7706 : tag_0_74; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_725 = 7'h4b == index ? _GEN_7706 : tag_0_75; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_726 = 7'h4c == index ? _GEN_7706 : tag_0_76; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_727 = 7'h4d == index ? _GEN_7706 : tag_0_77; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_728 = 7'h4e == index ? _GEN_7706 : tag_0_78; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_729 = 7'h4f == index ? _GEN_7706 : tag_0_79; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_730 = 7'h50 == index ? _GEN_7706 : tag_0_80; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_731 = 7'h51 == index ? _GEN_7706 : tag_0_81; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_732 = 7'h52 == index ? _GEN_7706 : tag_0_82; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_733 = 7'h53 == index ? _GEN_7706 : tag_0_83; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_734 = 7'h54 == index ? _GEN_7706 : tag_0_84; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_735 = 7'h55 == index ? _GEN_7706 : tag_0_85; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_736 = 7'h56 == index ? _GEN_7706 : tag_0_86; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_737 = 7'h57 == index ? _GEN_7706 : tag_0_87; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_738 = 7'h58 == index ? _GEN_7706 : tag_0_88; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_739 = 7'h59 == index ? _GEN_7706 : tag_0_89; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_740 = 7'h5a == index ? _GEN_7706 : tag_0_90; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_741 = 7'h5b == index ? _GEN_7706 : tag_0_91; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_742 = 7'h5c == index ? _GEN_7706 : tag_0_92; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_743 = 7'h5d == index ? _GEN_7706 : tag_0_93; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_744 = 7'h5e == index ? _GEN_7706 : tag_0_94; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_745 = 7'h5f == index ? _GEN_7706 : tag_0_95; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_746 = 7'h60 == index ? _GEN_7706 : tag_0_96; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_747 = 7'h61 == index ? _GEN_7706 : tag_0_97; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_748 = 7'h62 == index ? _GEN_7706 : tag_0_98; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_749 = 7'h63 == index ? _GEN_7706 : tag_0_99; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_750 = 7'h64 == index ? _GEN_7706 : tag_0_100; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_751 = 7'h65 == index ? _GEN_7706 : tag_0_101; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_752 = 7'h66 == index ? _GEN_7706 : tag_0_102; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_753 = 7'h67 == index ? _GEN_7706 : tag_0_103; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_754 = 7'h68 == index ? _GEN_7706 : tag_0_104; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_755 = 7'h69 == index ? _GEN_7706 : tag_0_105; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_756 = 7'h6a == index ? _GEN_7706 : tag_0_106; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_757 = 7'h6b == index ? _GEN_7706 : tag_0_107; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_758 = 7'h6c == index ? _GEN_7706 : tag_0_108; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_759 = 7'h6d == index ? _GEN_7706 : tag_0_109; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_760 = 7'h6e == index ? _GEN_7706 : tag_0_110; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_761 = 7'h6f == index ? _GEN_7706 : tag_0_111; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_762 = 7'h70 == index ? _GEN_7706 : tag_0_112; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_763 = 7'h71 == index ? _GEN_7706 : tag_0_113; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_764 = 7'h72 == index ? _GEN_7706 : tag_0_114; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_765 = 7'h73 == index ? _GEN_7706 : tag_0_115; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_766 = 7'h74 == index ? _GEN_7706 : tag_0_116; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_767 = 7'h75 == index ? _GEN_7706 : tag_0_117; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_768 = 7'h76 == index ? _GEN_7706 : tag_0_118; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_769 = 7'h77 == index ? _GEN_7706 : tag_0_119; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_770 = 7'h78 == index ? _GEN_7706 : tag_0_120; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_771 = 7'h79 == index ? _GEN_7706 : tag_0_121; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_772 = 7'h7a == index ? _GEN_7706 : tag_0_122; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_773 = 7'h7b == index ? _GEN_7706 : tag_0_123; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_774 = 7'h7c == index ? _GEN_7706 : tag_0_124; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_775 = 7'h7d == index ? _GEN_7706 : tag_0_125; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_776 = 7'h7e == index ? _GEN_7706 : tag_0_126; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_777 = 7'h7f == index ? _GEN_7706 : tag_0_127; // @[i_cache.scala 19:24 88:{30,30}]
  wire  _GEN_7710 = 7'h0 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_778 = 7'h0 == index | valid_0_0; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7712 = 7'h1 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_779 = 7'h1 == index | valid_0_1; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7714 = 7'h2 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_780 = 7'h2 == index | valid_0_2; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7718 = 7'h3 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_781 = 7'h3 == index | valid_0_3; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7727 = 7'h4 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_782 = 7'h4 == index | valid_0_4; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7729 = 7'h5 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_783 = 7'h5 == index | valid_0_5; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7731 = 7'h6 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_784 = 7'h6 == index | valid_0_6; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7733 = 7'h7 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_785 = 7'h7 == index | valid_0_7; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7738 = 7'h8 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_786 = 7'h8 == index | valid_0_8; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7739 = 7'h9 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_787 = 7'h9 == index | valid_0_9; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7740 = 7'ha == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_788 = 7'ha == index | valid_0_10; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7741 = 7'hb == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_789 = 7'hb == index | valid_0_11; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7742 = 7'hc == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_790 = 7'hc == index | valid_0_12; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7743 = 7'hd == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_791 = 7'hd == index | valid_0_13; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7744 = 7'he == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_792 = 7'he == index | valid_0_14; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7745 = 7'hf == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_793 = 7'hf == index | valid_0_15; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7746 = 7'h10 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_794 = 7'h10 == index | valid_0_16; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7747 = 7'h11 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_795 = 7'h11 == index | valid_0_17; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7748 = 7'h12 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_796 = 7'h12 == index | valid_0_18; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7749 = 7'h13 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_797 = 7'h13 == index | valid_0_19; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7750 = 7'h14 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_798 = 7'h14 == index | valid_0_20; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7751 = 7'h15 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_799 = 7'h15 == index | valid_0_21; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7752 = 7'h16 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_800 = 7'h16 == index | valid_0_22; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7753 = 7'h17 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_801 = 7'h17 == index | valid_0_23; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7754 = 7'h18 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_802 = 7'h18 == index | valid_0_24; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7755 = 7'h19 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_803 = 7'h19 == index | valid_0_25; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7756 = 7'h1a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_804 = 7'h1a == index | valid_0_26; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7757 = 7'h1b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_805 = 7'h1b == index | valid_0_27; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7758 = 7'h1c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_806 = 7'h1c == index | valid_0_28; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7759 = 7'h1d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_807 = 7'h1d == index | valid_0_29; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7760 = 7'h1e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_808 = 7'h1e == index | valid_0_30; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7761 = 7'h1f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_809 = 7'h1f == index | valid_0_31; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7762 = 7'h20 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_810 = 7'h20 == index | valid_0_32; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7763 = 7'h21 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_811 = 7'h21 == index | valid_0_33; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7764 = 7'h22 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_812 = 7'h22 == index | valid_0_34; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7765 = 7'h23 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_813 = 7'h23 == index | valid_0_35; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7766 = 7'h24 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_814 = 7'h24 == index | valid_0_36; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7767 = 7'h25 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_815 = 7'h25 == index | valid_0_37; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7768 = 7'h26 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_816 = 7'h26 == index | valid_0_38; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7769 = 7'h27 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_817 = 7'h27 == index | valid_0_39; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7770 = 7'h28 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_818 = 7'h28 == index | valid_0_40; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7771 = 7'h29 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_819 = 7'h29 == index | valid_0_41; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7772 = 7'h2a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_820 = 7'h2a == index | valid_0_42; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7773 = 7'h2b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_821 = 7'h2b == index | valid_0_43; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7774 = 7'h2c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_822 = 7'h2c == index | valid_0_44; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7775 = 7'h2d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_823 = 7'h2d == index | valid_0_45; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7776 = 7'h2e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_824 = 7'h2e == index | valid_0_46; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7777 = 7'h2f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_825 = 7'h2f == index | valid_0_47; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7778 = 7'h30 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_826 = 7'h30 == index | valid_0_48; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7779 = 7'h31 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_827 = 7'h31 == index | valid_0_49; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7780 = 7'h32 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_828 = 7'h32 == index | valid_0_50; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7781 = 7'h33 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_829 = 7'h33 == index | valid_0_51; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7782 = 7'h34 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_830 = 7'h34 == index | valid_0_52; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7783 = 7'h35 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_831 = 7'h35 == index | valid_0_53; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7784 = 7'h36 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_832 = 7'h36 == index | valid_0_54; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7785 = 7'h37 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_833 = 7'h37 == index | valid_0_55; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7786 = 7'h38 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_834 = 7'h38 == index | valid_0_56; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7787 = 7'h39 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_835 = 7'h39 == index | valid_0_57; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7788 = 7'h3a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_836 = 7'h3a == index | valid_0_58; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7789 = 7'h3b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_837 = 7'h3b == index | valid_0_59; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7790 = 7'h3c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_838 = 7'h3c == index | valid_0_60; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7791 = 7'h3d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_839 = 7'h3d == index | valid_0_61; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7792 = 7'h3e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_840 = 7'h3e == index | valid_0_62; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7793 = 7'h3f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_841 = 7'h3f == index | valid_0_63; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7794 = 7'h40 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_842 = 7'h40 == index | valid_0_64; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7795 = 7'h41 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_843 = 7'h41 == index | valid_0_65; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7796 = 7'h42 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_844 = 7'h42 == index | valid_0_66; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7797 = 7'h43 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_845 = 7'h43 == index | valid_0_67; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7798 = 7'h44 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_846 = 7'h44 == index | valid_0_68; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7799 = 7'h45 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_847 = 7'h45 == index | valid_0_69; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7800 = 7'h46 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_848 = 7'h46 == index | valid_0_70; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7801 = 7'h47 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_849 = 7'h47 == index | valid_0_71; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7802 = 7'h48 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_850 = 7'h48 == index | valid_0_72; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7803 = 7'h49 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_851 = 7'h49 == index | valid_0_73; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7804 = 7'h4a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_852 = 7'h4a == index | valid_0_74; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7805 = 7'h4b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_853 = 7'h4b == index | valid_0_75; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7806 = 7'h4c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_854 = 7'h4c == index | valid_0_76; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7807 = 7'h4d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_855 = 7'h4d == index | valid_0_77; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7808 = 7'h4e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_856 = 7'h4e == index | valid_0_78; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7809 = 7'h4f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_857 = 7'h4f == index | valid_0_79; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7810 = 7'h50 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_858 = 7'h50 == index | valid_0_80; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7811 = 7'h51 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_859 = 7'h51 == index | valid_0_81; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7812 = 7'h52 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_860 = 7'h52 == index | valid_0_82; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7813 = 7'h53 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_861 = 7'h53 == index | valid_0_83; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7814 = 7'h54 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_862 = 7'h54 == index | valid_0_84; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7815 = 7'h55 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_863 = 7'h55 == index | valid_0_85; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7816 = 7'h56 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_864 = 7'h56 == index | valid_0_86; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7817 = 7'h57 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_865 = 7'h57 == index | valid_0_87; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7818 = 7'h58 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_866 = 7'h58 == index | valid_0_88; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7819 = 7'h59 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_867 = 7'h59 == index | valid_0_89; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7820 = 7'h5a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_868 = 7'h5a == index | valid_0_90; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7821 = 7'h5b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_869 = 7'h5b == index | valid_0_91; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7822 = 7'h5c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_870 = 7'h5c == index | valid_0_92; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7823 = 7'h5d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_871 = 7'h5d == index | valid_0_93; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7824 = 7'h5e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_872 = 7'h5e == index | valid_0_94; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7825 = 7'h5f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_873 = 7'h5f == index | valid_0_95; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7826 = 7'h60 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_874 = 7'h60 == index | valid_0_96; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7827 = 7'h61 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_875 = 7'h61 == index | valid_0_97; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7828 = 7'h62 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_876 = 7'h62 == index | valid_0_98; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7829 = 7'h63 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_877 = 7'h63 == index | valid_0_99; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7830 = 7'h64 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_878 = 7'h64 == index | valid_0_100; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7831 = 7'h65 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_879 = 7'h65 == index | valid_0_101; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7832 = 7'h66 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_880 = 7'h66 == index | valid_0_102; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7833 = 7'h67 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_881 = 7'h67 == index | valid_0_103; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7834 = 7'h68 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_882 = 7'h68 == index | valid_0_104; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7835 = 7'h69 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_883 = 7'h69 == index | valid_0_105; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7836 = 7'h6a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_884 = 7'h6a == index | valid_0_106; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7837 = 7'h6b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_885 = 7'h6b == index | valid_0_107; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7838 = 7'h6c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_886 = 7'h6c == index | valid_0_108; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7839 = 7'h6d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_887 = 7'h6d == index | valid_0_109; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7840 = 7'h6e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_888 = 7'h6e == index | valid_0_110; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7841 = 7'h6f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_889 = 7'h6f == index | valid_0_111; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7842 = 7'h70 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_890 = 7'h70 == index | valid_0_112; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7843 = 7'h71 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_891 = 7'h71 == index | valid_0_113; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7844 = 7'h72 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_892 = 7'h72 == index | valid_0_114; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7845 = 7'h73 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_893 = 7'h73 == index | valid_0_115; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7846 = 7'h74 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_894 = 7'h74 == index | valid_0_116; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7847 = 7'h75 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_895 = 7'h75 == index | valid_0_117; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7848 = 7'h76 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_896 = 7'h76 == index | valid_0_118; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7849 = 7'h77 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_897 = 7'h77 == index | valid_0_119; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7850 = 7'h78 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_898 = 7'h78 == index | valid_0_120; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7851 = 7'h79 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_899 = 7'h79 == index | valid_0_121; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7852 = 7'h7a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_900 = 7'h7a == index | valid_0_122; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7853 = 7'h7b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_901 = 7'h7b == index | valid_0_123; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7854 = 7'h7c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_902 = 7'h7c == index | valid_0_124; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7855 = 7'h7d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_903 = 7'h7d == index | valid_0_125; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7856 = 7'h7e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_904 = 7'h7e == index | valid_0_126; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7857 = 7'h7f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_905 = 7'h7f == index | valid_0_127; // @[i_cache.scala 21:26 89:{32,32}]
  wire [63:0] _GEN_906 = 7'h0 == index ? receive_data : ram_1_0; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_907 = 7'h1 == index ? receive_data : ram_1_1; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_908 = 7'h2 == index ? receive_data : ram_1_2; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_909 = 7'h3 == index ? receive_data : ram_1_3; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_910 = 7'h4 == index ? receive_data : ram_1_4; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_911 = 7'h5 == index ? receive_data : ram_1_5; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_912 = 7'h6 == index ? receive_data : ram_1_6; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_913 = 7'h7 == index ? receive_data : ram_1_7; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_914 = 7'h8 == index ? receive_data : ram_1_8; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_915 = 7'h9 == index ? receive_data : ram_1_9; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_916 = 7'ha == index ? receive_data : ram_1_10; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_917 = 7'hb == index ? receive_data : ram_1_11; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_918 = 7'hc == index ? receive_data : ram_1_12; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_919 = 7'hd == index ? receive_data : ram_1_13; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_920 = 7'he == index ? receive_data : ram_1_14; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_921 = 7'hf == index ? receive_data : ram_1_15; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_922 = 7'h10 == index ? receive_data : ram_1_16; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_923 = 7'h11 == index ? receive_data : ram_1_17; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_924 = 7'h12 == index ? receive_data : ram_1_18; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_925 = 7'h13 == index ? receive_data : ram_1_19; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_926 = 7'h14 == index ? receive_data : ram_1_20; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_927 = 7'h15 == index ? receive_data : ram_1_21; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_928 = 7'h16 == index ? receive_data : ram_1_22; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_929 = 7'h17 == index ? receive_data : ram_1_23; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_930 = 7'h18 == index ? receive_data : ram_1_24; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_931 = 7'h19 == index ? receive_data : ram_1_25; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_932 = 7'h1a == index ? receive_data : ram_1_26; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_933 = 7'h1b == index ? receive_data : ram_1_27; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_934 = 7'h1c == index ? receive_data : ram_1_28; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_935 = 7'h1d == index ? receive_data : ram_1_29; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_936 = 7'h1e == index ? receive_data : ram_1_30; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_937 = 7'h1f == index ? receive_data : ram_1_31; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_938 = 7'h20 == index ? receive_data : ram_1_32; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_939 = 7'h21 == index ? receive_data : ram_1_33; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_940 = 7'h22 == index ? receive_data : ram_1_34; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_941 = 7'h23 == index ? receive_data : ram_1_35; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_942 = 7'h24 == index ? receive_data : ram_1_36; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_943 = 7'h25 == index ? receive_data : ram_1_37; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_944 = 7'h26 == index ? receive_data : ram_1_38; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_945 = 7'h27 == index ? receive_data : ram_1_39; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_946 = 7'h28 == index ? receive_data : ram_1_40; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_947 = 7'h29 == index ? receive_data : ram_1_41; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_948 = 7'h2a == index ? receive_data : ram_1_42; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_949 = 7'h2b == index ? receive_data : ram_1_43; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_950 = 7'h2c == index ? receive_data : ram_1_44; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_951 = 7'h2d == index ? receive_data : ram_1_45; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_952 = 7'h2e == index ? receive_data : ram_1_46; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_953 = 7'h2f == index ? receive_data : ram_1_47; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_954 = 7'h30 == index ? receive_data : ram_1_48; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_955 = 7'h31 == index ? receive_data : ram_1_49; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_956 = 7'h32 == index ? receive_data : ram_1_50; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_957 = 7'h33 == index ? receive_data : ram_1_51; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_958 = 7'h34 == index ? receive_data : ram_1_52; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_959 = 7'h35 == index ? receive_data : ram_1_53; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_960 = 7'h36 == index ? receive_data : ram_1_54; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_961 = 7'h37 == index ? receive_data : ram_1_55; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_962 = 7'h38 == index ? receive_data : ram_1_56; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_963 = 7'h39 == index ? receive_data : ram_1_57; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_964 = 7'h3a == index ? receive_data : ram_1_58; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_965 = 7'h3b == index ? receive_data : ram_1_59; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_966 = 7'h3c == index ? receive_data : ram_1_60; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_967 = 7'h3d == index ? receive_data : ram_1_61; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_968 = 7'h3e == index ? receive_data : ram_1_62; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_969 = 7'h3f == index ? receive_data : ram_1_63; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_970 = 7'h40 == index ? receive_data : ram_1_64; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_971 = 7'h41 == index ? receive_data : ram_1_65; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_972 = 7'h42 == index ? receive_data : ram_1_66; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_973 = 7'h43 == index ? receive_data : ram_1_67; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_974 = 7'h44 == index ? receive_data : ram_1_68; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_975 = 7'h45 == index ? receive_data : ram_1_69; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_976 = 7'h46 == index ? receive_data : ram_1_70; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_977 = 7'h47 == index ? receive_data : ram_1_71; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_978 = 7'h48 == index ? receive_data : ram_1_72; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_979 = 7'h49 == index ? receive_data : ram_1_73; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_980 = 7'h4a == index ? receive_data : ram_1_74; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_981 = 7'h4b == index ? receive_data : ram_1_75; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_982 = 7'h4c == index ? receive_data : ram_1_76; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_983 = 7'h4d == index ? receive_data : ram_1_77; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_984 = 7'h4e == index ? receive_data : ram_1_78; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_985 = 7'h4f == index ? receive_data : ram_1_79; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_986 = 7'h50 == index ? receive_data : ram_1_80; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_987 = 7'h51 == index ? receive_data : ram_1_81; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_988 = 7'h52 == index ? receive_data : ram_1_82; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_989 = 7'h53 == index ? receive_data : ram_1_83; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_990 = 7'h54 == index ? receive_data : ram_1_84; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_991 = 7'h55 == index ? receive_data : ram_1_85; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_992 = 7'h56 == index ? receive_data : ram_1_86; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_993 = 7'h57 == index ? receive_data : ram_1_87; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_994 = 7'h58 == index ? receive_data : ram_1_88; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_995 = 7'h59 == index ? receive_data : ram_1_89; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_996 = 7'h5a == index ? receive_data : ram_1_90; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_997 = 7'h5b == index ? receive_data : ram_1_91; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_998 = 7'h5c == index ? receive_data : ram_1_92; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_999 = 7'h5d == index ? receive_data : ram_1_93; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1000 = 7'h5e == index ? receive_data : ram_1_94; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1001 = 7'h5f == index ? receive_data : ram_1_95; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1002 = 7'h60 == index ? receive_data : ram_1_96; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1003 = 7'h61 == index ? receive_data : ram_1_97; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1004 = 7'h62 == index ? receive_data : ram_1_98; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1005 = 7'h63 == index ? receive_data : ram_1_99; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1006 = 7'h64 == index ? receive_data : ram_1_100; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1007 = 7'h65 == index ? receive_data : ram_1_101; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1008 = 7'h66 == index ? receive_data : ram_1_102; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1009 = 7'h67 == index ? receive_data : ram_1_103; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1010 = 7'h68 == index ? receive_data : ram_1_104; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1011 = 7'h69 == index ? receive_data : ram_1_105; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1012 = 7'h6a == index ? receive_data : ram_1_106; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1013 = 7'h6b == index ? receive_data : ram_1_107; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1014 = 7'h6c == index ? receive_data : ram_1_108; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1015 = 7'h6d == index ? receive_data : ram_1_109; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1016 = 7'h6e == index ? receive_data : ram_1_110; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1017 = 7'h6f == index ? receive_data : ram_1_111; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1018 = 7'h70 == index ? receive_data : ram_1_112; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1019 = 7'h71 == index ? receive_data : ram_1_113; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1020 = 7'h72 == index ? receive_data : ram_1_114; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1021 = 7'h73 == index ? receive_data : ram_1_115; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1022 = 7'h74 == index ? receive_data : ram_1_116; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1023 = 7'h75 == index ? receive_data : ram_1_117; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1024 = 7'h76 == index ? receive_data : ram_1_118; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1025 = 7'h77 == index ? receive_data : ram_1_119; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1026 = 7'h78 == index ? receive_data : ram_1_120; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1027 = 7'h79 == index ? receive_data : ram_1_121; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1028 = 7'h7a == index ? receive_data : ram_1_122; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1029 = 7'h7b == index ? receive_data : ram_1_123; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1030 = 7'h7c == index ? receive_data : ram_1_124; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1031 = 7'h7d == index ? receive_data : ram_1_125; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1032 = 7'h7e == index ? receive_data : ram_1_126; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1033 = 7'h7f == index ? receive_data : ram_1_127; // @[i_cache.scala 18:24 92:{30,30}]
  wire [31:0] _GEN_1034 = 7'h0 == index ? _GEN_7706 : tag_1_0; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1035 = 7'h1 == index ? _GEN_7706 : tag_1_1; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1036 = 7'h2 == index ? _GEN_7706 : tag_1_2; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1037 = 7'h3 == index ? _GEN_7706 : tag_1_3; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1038 = 7'h4 == index ? _GEN_7706 : tag_1_4; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1039 = 7'h5 == index ? _GEN_7706 : tag_1_5; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1040 = 7'h6 == index ? _GEN_7706 : tag_1_6; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1041 = 7'h7 == index ? _GEN_7706 : tag_1_7; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1042 = 7'h8 == index ? _GEN_7706 : tag_1_8; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1043 = 7'h9 == index ? _GEN_7706 : tag_1_9; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1044 = 7'ha == index ? _GEN_7706 : tag_1_10; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1045 = 7'hb == index ? _GEN_7706 : tag_1_11; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1046 = 7'hc == index ? _GEN_7706 : tag_1_12; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1047 = 7'hd == index ? _GEN_7706 : tag_1_13; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1048 = 7'he == index ? _GEN_7706 : tag_1_14; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1049 = 7'hf == index ? _GEN_7706 : tag_1_15; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1050 = 7'h10 == index ? _GEN_7706 : tag_1_16; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1051 = 7'h11 == index ? _GEN_7706 : tag_1_17; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1052 = 7'h12 == index ? _GEN_7706 : tag_1_18; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1053 = 7'h13 == index ? _GEN_7706 : tag_1_19; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1054 = 7'h14 == index ? _GEN_7706 : tag_1_20; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1055 = 7'h15 == index ? _GEN_7706 : tag_1_21; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1056 = 7'h16 == index ? _GEN_7706 : tag_1_22; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1057 = 7'h17 == index ? _GEN_7706 : tag_1_23; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1058 = 7'h18 == index ? _GEN_7706 : tag_1_24; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1059 = 7'h19 == index ? _GEN_7706 : tag_1_25; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1060 = 7'h1a == index ? _GEN_7706 : tag_1_26; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1061 = 7'h1b == index ? _GEN_7706 : tag_1_27; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1062 = 7'h1c == index ? _GEN_7706 : tag_1_28; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1063 = 7'h1d == index ? _GEN_7706 : tag_1_29; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1064 = 7'h1e == index ? _GEN_7706 : tag_1_30; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1065 = 7'h1f == index ? _GEN_7706 : tag_1_31; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1066 = 7'h20 == index ? _GEN_7706 : tag_1_32; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1067 = 7'h21 == index ? _GEN_7706 : tag_1_33; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1068 = 7'h22 == index ? _GEN_7706 : tag_1_34; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1069 = 7'h23 == index ? _GEN_7706 : tag_1_35; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1070 = 7'h24 == index ? _GEN_7706 : tag_1_36; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1071 = 7'h25 == index ? _GEN_7706 : tag_1_37; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1072 = 7'h26 == index ? _GEN_7706 : tag_1_38; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1073 = 7'h27 == index ? _GEN_7706 : tag_1_39; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1074 = 7'h28 == index ? _GEN_7706 : tag_1_40; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1075 = 7'h29 == index ? _GEN_7706 : tag_1_41; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1076 = 7'h2a == index ? _GEN_7706 : tag_1_42; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1077 = 7'h2b == index ? _GEN_7706 : tag_1_43; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1078 = 7'h2c == index ? _GEN_7706 : tag_1_44; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1079 = 7'h2d == index ? _GEN_7706 : tag_1_45; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1080 = 7'h2e == index ? _GEN_7706 : tag_1_46; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1081 = 7'h2f == index ? _GEN_7706 : tag_1_47; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1082 = 7'h30 == index ? _GEN_7706 : tag_1_48; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1083 = 7'h31 == index ? _GEN_7706 : tag_1_49; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1084 = 7'h32 == index ? _GEN_7706 : tag_1_50; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1085 = 7'h33 == index ? _GEN_7706 : tag_1_51; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1086 = 7'h34 == index ? _GEN_7706 : tag_1_52; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1087 = 7'h35 == index ? _GEN_7706 : tag_1_53; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1088 = 7'h36 == index ? _GEN_7706 : tag_1_54; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1089 = 7'h37 == index ? _GEN_7706 : tag_1_55; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1090 = 7'h38 == index ? _GEN_7706 : tag_1_56; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1091 = 7'h39 == index ? _GEN_7706 : tag_1_57; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1092 = 7'h3a == index ? _GEN_7706 : tag_1_58; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1093 = 7'h3b == index ? _GEN_7706 : tag_1_59; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1094 = 7'h3c == index ? _GEN_7706 : tag_1_60; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1095 = 7'h3d == index ? _GEN_7706 : tag_1_61; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1096 = 7'h3e == index ? _GEN_7706 : tag_1_62; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1097 = 7'h3f == index ? _GEN_7706 : tag_1_63; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1098 = 7'h40 == index ? _GEN_7706 : tag_1_64; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1099 = 7'h41 == index ? _GEN_7706 : tag_1_65; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1100 = 7'h42 == index ? _GEN_7706 : tag_1_66; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1101 = 7'h43 == index ? _GEN_7706 : tag_1_67; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1102 = 7'h44 == index ? _GEN_7706 : tag_1_68; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1103 = 7'h45 == index ? _GEN_7706 : tag_1_69; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1104 = 7'h46 == index ? _GEN_7706 : tag_1_70; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1105 = 7'h47 == index ? _GEN_7706 : tag_1_71; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1106 = 7'h48 == index ? _GEN_7706 : tag_1_72; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1107 = 7'h49 == index ? _GEN_7706 : tag_1_73; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1108 = 7'h4a == index ? _GEN_7706 : tag_1_74; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1109 = 7'h4b == index ? _GEN_7706 : tag_1_75; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1110 = 7'h4c == index ? _GEN_7706 : tag_1_76; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1111 = 7'h4d == index ? _GEN_7706 : tag_1_77; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1112 = 7'h4e == index ? _GEN_7706 : tag_1_78; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1113 = 7'h4f == index ? _GEN_7706 : tag_1_79; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1114 = 7'h50 == index ? _GEN_7706 : tag_1_80; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1115 = 7'h51 == index ? _GEN_7706 : tag_1_81; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1116 = 7'h52 == index ? _GEN_7706 : tag_1_82; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1117 = 7'h53 == index ? _GEN_7706 : tag_1_83; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1118 = 7'h54 == index ? _GEN_7706 : tag_1_84; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1119 = 7'h55 == index ? _GEN_7706 : tag_1_85; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1120 = 7'h56 == index ? _GEN_7706 : tag_1_86; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1121 = 7'h57 == index ? _GEN_7706 : tag_1_87; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1122 = 7'h58 == index ? _GEN_7706 : tag_1_88; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1123 = 7'h59 == index ? _GEN_7706 : tag_1_89; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1124 = 7'h5a == index ? _GEN_7706 : tag_1_90; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1125 = 7'h5b == index ? _GEN_7706 : tag_1_91; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1126 = 7'h5c == index ? _GEN_7706 : tag_1_92; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1127 = 7'h5d == index ? _GEN_7706 : tag_1_93; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1128 = 7'h5e == index ? _GEN_7706 : tag_1_94; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1129 = 7'h5f == index ? _GEN_7706 : tag_1_95; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1130 = 7'h60 == index ? _GEN_7706 : tag_1_96; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1131 = 7'h61 == index ? _GEN_7706 : tag_1_97; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1132 = 7'h62 == index ? _GEN_7706 : tag_1_98; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1133 = 7'h63 == index ? _GEN_7706 : tag_1_99; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1134 = 7'h64 == index ? _GEN_7706 : tag_1_100; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1135 = 7'h65 == index ? _GEN_7706 : tag_1_101; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1136 = 7'h66 == index ? _GEN_7706 : tag_1_102; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1137 = 7'h67 == index ? _GEN_7706 : tag_1_103; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1138 = 7'h68 == index ? _GEN_7706 : tag_1_104; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1139 = 7'h69 == index ? _GEN_7706 : tag_1_105; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1140 = 7'h6a == index ? _GEN_7706 : tag_1_106; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1141 = 7'h6b == index ? _GEN_7706 : tag_1_107; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1142 = 7'h6c == index ? _GEN_7706 : tag_1_108; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1143 = 7'h6d == index ? _GEN_7706 : tag_1_109; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1144 = 7'h6e == index ? _GEN_7706 : tag_1_110; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1145 = 7'h6f == index ? _GEN_7706 : tag_1_111; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1146 = 7'h70 == index ? _GEN_7706 : tag_1_112; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1147 = 7'h71 == index ? _GEN_7706 : tag_1_113; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1148 = 7'h72 == index ? _GEN_7706 : tag_1_114; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1149 = 7'h73 == index ? _GEN_7706 : tag_1_115; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1150 = 7'h74 == index ? _GEN_7706 : tag_1_116; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1151 = 7'h75 == index ? _GEN_7706 : tag_1_117; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1152 = 7'h76 == index ? _GEN_7706 : tag_1_118; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1153 = 7'h77 == index ? _GEN_7706 : tag_1_119; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1154 = 7'h78 == index ? _GEN_7706 : tag_1_120; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1155 = 7'h79 == index ? _GEN_7706 : tag_1_121; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1156 = 7'h7a == index ? _GEN_7706 : tag_1_122; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1157 = 7'h7b == index ? _GEN_7706 : tag_1_123; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1158 = 7'h7c == index ? _GEN_7706 : tag_1_124; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1159 = 7'h7d == index ? _GEN_7706 : tag_1_125; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1160 = 7'h7e == index ? _GEN_7706 : tag_1_126; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1161 = 7'h7f == index ? _GEN_7706 : tag_1_127; // @[i_cache.scala 20:24 93:{30,30}]
  wire  _GEN_1162 = _GEN_7710 | valid_1_0; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1163 = _GEN_7712 | valid_1_1; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1164 = _GEN_7714 | valid_1_2; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1165 = _GEN_7718 | valid_1_3; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1166 = _GEN_7727 | valid_1_4; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1167 = _GEN_7729 | valid_1_5; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1168 = _GEN_7731 | valid_1_6; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1169 = _GEN_7733 | valid_1_7; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1170 = _GEN_7738 | valid_1_8; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1171 = _GEN_7739 | valid_1_9; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1172 = _GEN_7740 | valid_1_10; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1173 = _GEN_7741 | valid_1_11; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1174 = _GEN_7742 | valid_1_12; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1175 = _GEN_7743 | valid_1_13; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1176 = _GEN_7744 | valid_1_14; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1177 = _GEN_7745 | valid_1_15; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1178 = _GEN_7746 | valid_1_16; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1179 = _GEN_7747 | valid_1_17; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1180 = _GEN_7748 | valid_1_18; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1181 = _GEN_7749 | valid_1_19; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1182 = _GEN_7750 | valid_1_20; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1183 = _GEN_7751 | valid_1_21; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1184 = _GEN_7752 | valid_1_22; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1185 = _GEN_7753 | valid_1_23; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1186 = _GEN_7754 | valid_1_24; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1187 = _GEN_7755 | valid_1_25; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1188 = _GEN_7756 | valid_1_26; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1189 = _GEN_7757 | valid_1_27; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1190 = _GEN_7758 | valid_1_28; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1191 = _GEN_7759 | valid_1_29; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1192 = _GEN_7760 | valid_1_30; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1193 = _GEN_7761 | valid_1_31; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1194 = _GEN_7762 | valid_1_32; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1195 = _GEN_7763 | valid_1_33; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1196 = _GEN_7764 | valid_1_34; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1197 = _GEN_7765 | valid_1_35; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1198 = _GEN_7766 | valid_1_36; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1199 = _GEN_7767 | valid_1_37; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1200 = _GEN_7768 | valid_1_38; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1201 = _GEN_7769 | valid_1_39; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1202 = _GEN_7770 | valid_1_40; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1203 = _GEN_7771 | valid_1_41; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1204 = _GEN_7772 | valid_1_42; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1205 = _GEN_7773 | valid_1_43; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1206 = _GEN_7774 | valid_1_44; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1207 = _GEN_7775 | valid_1_45; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1208 = _GEN_7776 | valid_1_46; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1209 = _GEN_7777 | valid_1_47; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1210 = _GEN_7778 | valid_1_48; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1211 = _GEN_7779 | valid_1_49; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1212 = _GEN_7780 | valid_1_50; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1213 = _GEN_7781 | valid_1_51; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1214 = _GEN_7782 | valid_1_52; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1215 = _GEN_7783 | valid_1_53; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1216 = _GEN_7784 | valid_1_54; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1217 = _GEN_7785 | valid_1_55; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1218 = _GEN_7786 | valid_1_56; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1219 = _GEN_7787 | valid_1_57; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1220 = _GEN_7788 | valid_1_58; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1221 = _GEN_7789 | valid_1_59; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1222 = _GEN_7790 | valid_1_60; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1223 = _GEN_7791 | valid_1_61; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1224 = _GEN_7792 | valid_1_62; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1225 = _GEN_7793 | valid_1_63; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1226 = _GEN_7794 | valid_1_64; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1227 = _GEN_7795 | valid_1_65; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1228 = _GEN_7796 | valid_1_66; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1229 = _GEN_7797 | valid_1_67; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1230 = _GEN_7798 | valid_1_68; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1231 = _GEN_7799 | valid_1_69; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1232 = _GEN_7800 | valid_1_70; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1233 = _GEN_7801 | valid_1_71; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1234 = _GEN_7802 | valid_1_72; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1235 = _GEN_7803 | valid_1_73; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1236 = _GEN_7804 | valid_1_74; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1237 = _GEN_7805 | valid_1_75; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1238 = _GEN_7806 | valid_1_76; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1239 = _GEN_7807 | valid_1_77; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1240 = _GEN_7808 | valid_1_78; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1241 = _GEN_7809 | valid_1_79; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1242 = _GEN_7810 | valid_1_80; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1243 = _GEN_7811 | valid_1_81; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1244 = _GEN_7812 | valid_1_82; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1245 = _GEN_7813 | valid_1_83; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1246 = _GEN_7814 | valid_1_84; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1247 = _GEN_7815 | valid_1_85; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1248 = _GEN_7816 | valid_1_86; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1249 = _GEN_7817 | valid_1_87; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1250 = _GEN_7818 | valid_1_88; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1251 = _GEN_7819 | valid_1_89; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1252 = _GEN_7820 | valid_1_90; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1253 = _GEN_7821 | valid_1_91; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1254 = _GEN_7822 | valid_1_92; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1255 = _GEN_7823 | valid_1_93; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1256 = _GEN_7824 | valid_1_94; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1257 = _GEN_7825 | valid_1_95; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1258 = _GEN_7826 | valid_1_96; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1259 = _GEN_7827 | valid_1_97; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1260 = _GEN_7828 | valid_1_98; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1261 = _GEN_7829 | valid_1_99; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1262 = _GEN_7830 | valid_1_100; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1263 = _GEN_7831 | valid_1_101; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1264 = _GEN_7832 | valid_1_102; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1265 = _GEN_7833 | valid_1_103; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1266 = _GEN_7834 | valid_1_104; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1267 = _GEN_7835 | valid_1_105; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1268 = _GEN_7836 | valid_1_106; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1269 = _GEN_7837 | valid_1_107; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1270 = _GEN_7838 | valid_1_108; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1271 = _GEN_7839 | valid_1_109; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1272 = _GEN_7840 | valid_1_110; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1273 = _GEN_7841 | valid_1_111; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1274 = _GEN_7842 | valid_1_112; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1275 = _GEN_7843 | valid_1_113; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1276 = _GEN_7844 | valid_1_114; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1277 = _GEN_7845 | valid_1_115; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1278 = _GEN_7846 | valid_1_116; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1279 = _GEN_7847 | valid_1_117; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1280 = _GEN_7848 | valid_1_118; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1281 = _GEN_7849 | valid_1_119; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1282 = _GEN_7850 | valid_1_120; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1283 = _GEN_7851 | valid_1_121; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1284 = _GEN_7852 | valid_1_122; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1285 = _GEN_7853 | valid_1_123; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1286 = _GEN_7854 | valid_1_124; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1287 = _GEN_7855 | valid_1_125; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1288 = _GEN_7856 | valid_1_126; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1289 = _GEN_7857 | valid_1_127; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _T_14 = ~quene; // @[i_cache.scala 97:27]
  wire [63:0] _GEN_2058 = ~quene ? _GEN_522 : ram_0_0; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2059 = ~quene ? _GEN_523 : ram_0_1; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2060 = ~quene ? _GEN_524 : ram_0_2; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2061 = ~quene ? _GEN_525 : ram_0_3; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2062 = ~quene ? _GEN_526 : ram_0_4; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2063 = ~quene ? _GEN_527 : ram_0_5; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2064 = ~quene ? _GEN_528 : ram_0_6; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2065 = ~quene ? _GEN_529 : ram_0_7; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2066 = ~quene ? _GEN_530 : ram_0_8; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2067 = ~quene ? _GEN_531 : ram_0_9; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2068 = ~quene ? _GEN_532 : ram_0_10; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2069 = ~quene ? _GEN_533 : ram_0_11; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2070 = ~quene ? _GEN_534 : ram_0_12; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2071 = ~quene ? _GEN_535 : ram_0_13; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2072 = ~quene ? _GEN_536 : ram_0_14; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2073 = ~quene ? _GEN_537 : ram_0_15; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2074 = ~quene ? _GEN_538 : ram_0_16; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2075 = ~quene ? _GEN_539 : ram_0_17; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2076 = ~quene ? _GEN_540 : ram_0_18; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2077 = ~quene ? _GEN_541 : ram_0_19; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2078 = ~quene ? _GEN_542 : ram_0_20; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2079 = ~quene ? _GEN_543 : ram_0_21; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2080 = ~quene ? _GEN_544 : ram_0_22; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2081 = ~quene ? _GEN_545 : ram_0_23; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2082 = ~quene ? _GEN_546 : ram_0_24; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2083 = ~quene ? _GEN_547 : ram_0_25; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2084 = ~quene ? _GEN_548 : ram_0_26; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2085 = ~quene ? _GEN_549 : ram_0_27; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2086 = ~quene ? _GEN_550 : ram_0_28; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2087 = ~quene ? _GEN_551 : ram_0_29; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2088 = ~quene ? _GEN_552 : ram_0_30; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2089 = ~quene ? _GEN_553 : ram_0_31; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2090 = ~quene ? _GEN_554 : ram_0_32; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2091 = ~quene ? _GEN_555 : ram_0_33; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2092 = ~quene ? _GEN_556 : ram_0_34; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2093 = ~quene ? _GEN_557 : ram_0_35; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2094 = ~quene ? _GEN_558 : ram_0_36; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2095 = ~quene ? _GEN_559 : ram_0_37; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2096 = ~quene ? _GEN_560 : ram_0_38; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2097 = ~quene ? _GEN_561 : ram_0_39; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2098 = ~quene ? _GEN_562 : ram_0_40; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2099 = ~quene ? _GEN_563 : ram_0_41; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2100 = ~quene ? _GEN_564 : ram_0_42; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2101 = ~quene ? _GEN_565 : ram_0_43; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2102 = ~quene ? _GEN_566 : ram_0_44; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2103 = ~quene ? _GEN_567 : ram_0_45; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2104 = ~quene ? _GEN_568 : ram_0_46; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2105 = ~quene ? _GEN_569 : ram_0_47; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2106 = ~quene ? _GEN_570 : ram_0_48; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2107 = ~quene ? _GEN_571 : ram_0_49; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2108 = ~quene ? _GEN_572 : ram_0_50; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2109 = ~quene ? _GEN_573 : ram_0_51; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2110 = ~quene ? _GEN_574 : ram_0_52; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2111 = ~quene ? _GEN_575 : ram_0_53; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2112 = ~quene ? _GEN_576 : ram_0_54; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2113 = ~quene ? _GEN_577 : ram_0_55; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2114 = ~quene ? _GEN_578 : ram_0_56; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2115 = ~quene ? _GEN_579 : ram_0_57; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2116 = ~quene ? _GEN_580 : ram_0_58; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2117 = ~quene ? _GEN_581 : ram_0_59; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2118 = ~quene ? _GEN_582 : ram_0_60; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2119 = ~quene ? _GEN_583 : ram_0_61; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2120 = ~quene ? _GEN_584 : ram_0_62; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2121 = ~quene ? _GEN_585 : ram_0_63; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2122 = ~quene ? _GEN_586 : ram_0_64; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2123 = ~quene ? _GEN_587 : ram_0_65; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2124 = ~quene ? _GEN_588 : ram_0_66; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2125 = ~quene ? _GEN_589 : ram_0_67; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2126 = ~quene ? _GEN_590 : ram_0_68; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2127 = ~quene ? _GEN_591 : ram_0_69; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2128 = ~quene ? _GEN_592 : ram_0_70; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2129 = ~quene ? _GEN_593 : ram_0_71; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2130 = ~quene ? _GEN_594 : ram_0_72; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2131 = ~quene ? _GEN_595 : ram_0_73; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2132 = ~quene ? _GEN_596 : ram_0_74; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2133 = ~quene ? _GEN_597 : ram_0_75; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2134 = ~quene ? _GEN_598 : ram_0_76; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2135 = ~quene ? _GEN_599 : ram_0_77; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2136 = ~quene ? _GEN_600 : ram_0_78; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2137 = ~quene ? _GEN_601 : ram_0_79; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2138 = ~quene ? _GEN_602 : ram_0_80; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2139 = ~quene ? _GEN_603 : ram_0_81; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2140 = ~quene ? _GEN_604 : ram_0_82; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2141 = ~quene ? _GEN_605 : ram_0_83; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2142 = ~quene ? _GEN_606 : ram_0_84; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2143 = ~quene ? _GEN_607 : ram_0_85; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2144 = ~quene ? _GEN_608 : ram_0_86; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2145 = ~quene ? _GEN_609 : ram_0_87; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2146 = ~quene ? _GEN_610 : ram_0_88; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2147 = ~quene ? _GEN_611 : ram_0_89; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2148 = ~quene ? _GEN_612 : ram_0_90; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2149 = ~quene ? _GEN_613 : ram_0_91; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2150 = ~quene ? _GEN_614 : ram_0_92; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2151 = ~quene ? _GEN_615 : ram_0_93; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2152 = ~quene ? _GEN_616 : ram_0_94; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2153 = ~quene ? _GEN_617 : ram_0_95; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2154 = ~quene ? _GEN_618 : ram_0_96; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2155 = ~quene ? _GEN_619 : ram_0_97; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2156 = ~quene ? _GEN_620 : ram_0_98; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2157 = ~quene ? _GEN_621 : ram_0_99; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2158 = ~quene ? _GEN_622 : ram_0_100; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2159 = ~quene ? _GEN_623 : ram_0_101; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2160 = ~quene ? _GEN_624 : ram_0_102; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2161 = ~quene ? _GEN_625 : ram_0_103; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2162 = ~quene ? _GEN_626 : ram_0_104; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2163 = ~quene ? _GEN_627 : ram_0_105; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2164 = ~quene ? _GEN_628 : ram_0_106; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2165 = ~quene ? _GEN_629 : ram_0_107; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2166 = ~quene ? _GEN_630 : ram_0_108; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2167 = ~quene ? _GEN_631 : ram_0_109; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2168 = ~quene ? _GEN_632 : ram_0_110; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2169 = ~quene ? _GEN_633 : ram_0_111; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2170 = ~quene ? _GEN_634 : ram_0_112; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2171 = ~quene ? _GEN_635 : ram_0_113; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2172 = ~quene ? _GEN_636 : ram_0_114; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2173 = ~quene ? _GEN_637 : ram_0_115; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2174 = ~quene ? _GEN_638 : ram_0_116; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2175 = ~quene ? _GEN_639 : ram_0_117; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2176 = ~quene ? _GEN_640 : ram_0_118; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2177 = ~quene ? _GEN_641 : ram_0_119; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2178 = ~quene ? _GEN_642 : ram_0_120; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2179 = ~quene ? _GEN_643 : ram_0_121; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2180 = ~quene ? _GEN_644 : ram_0_122; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2181 = ~quene ? _GEN_645 : ram_0_123; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2182 = ~quene ? _GEN_646 : ram_0_124; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2183 = ~quene ? _GEN_647 : ram_0_125; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2184 = ~quene ? _GEN_648 : ram_0_126; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2185 = ~quene ? _GEN_649 : ram_0_127; // @[i_cache.scala 17:24 97:34]
  wire [31:0] _GEN_2186 = ~quene ? _GEN_650 : tag_0_0; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2187 = ~quene ? _GEN_651 : tag_0_1; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2188 = ~quene ? _GEN_652 : tag_0_2; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2189 = ~quene ? _GEN_653 : tag_0_3; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2190 = ~quene ? _GEN_654 : tag_0_4; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2191 = ~quene ? _GEN_655 : tag_0_5; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2192 = ~quene ? _GEN_656 : tag_0_6; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2193 = ~quene ? _GEN_657 : tag_0_7; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2194 = ~quene ? _GEN_658 : tag_0_8; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2195 = ~quene ? _GEN_659 : tag_0_9; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2196 = ~quene ? _GEN_660 : tag_0_10; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2197 = ~quene ? _GEN_661 : tag_0_11; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2198 = ~quene ? _GEN_662 : tag_0_12; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2199 = ~quene ? _GEN_663 : tag_0_13; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2200 = ~quene ? _GEN_664 : tag_0_14; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2201 = ~quene ? _GEN_665 : tag_0_15; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2202 = ~quene ? _GEN_666 : tag_0_16; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2203 = ~quene ? _GEN_667 : tag_0_17; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2204 = ~quene ? _GEN_668 : tag_0_18; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2205 = ~quene ? _GEN_669 : tag_0_19; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2206 = ~quene ? _GEN_670 : tag_0_20; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2207 = ~quene ? _GEN_671 : tag_0_21; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2208 = ~quene ? _GEN_672 : tag_0_22; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2209 = ~quene ? _GEN_673 : tag_0_23; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2210 = ~quene ? _GEN_674 : tag_0_24; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2211 = ~quene ? _GEN_675 : tag_0_25; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2212 = ~quene ? _GEN_676 : tag_0_26; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2213 = ~quene ? _GEN_677 : tag_0_27; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2214 = ~quene ? _GEN_678 : tag_0_28; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2215 = ~quene ? _GEN_679 : tag_0_29; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2216 = ~quene ? _GEN_680 : tag_0_30; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2217 = ~quene ? _GEN_681 : tag_0_31; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2218 = ~quene ? _GEN_682 : tag_0_32; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2219 = ~quene ? _GEN_683 : tag_0_33; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2220 = ~quene ? _GEN_684 : tag_0_34; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2221 = ~quene ? _GEN_685 : tag_0_35; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2222 = ~quene ? _GEN_686 : tag_0_36; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2223 = ~quene ? _GEN_687 : tag_0_37; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2224 = ~quene ? _GEN_688 : tag_0_38; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2225 = ~quene ? _GEN_689 : tag_0_39; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2226 = ~quene ? _GEN_690 : tag_0_40; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2227 = ~quene ? _GEN_691 : tag_0_41; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2228 = ~quene ? _GEN_692 : tag_0_42; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2229 = ~quene ? _GEN_693 : tag_0_43; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2230 = ~quene ? _GEN_694 : tag_0_44; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2231 = ~quene ? _GEN_695 : tag_0_45; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2232 = ~quene ? _GEN_696 : tag_0_46; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2233 = ~quene ? _GEN_697 : tag_0_47; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2234 = ~quene ? _GEN_698 : tag_0_48; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2235 = ~quene ? _GEN_699 : tag_0_49; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2236 = ~quene ? _GEN_700 : tag_0_50; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2237 = ~quene ? _GEN_701 : tag_0_51; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2238 = ~quene ? _GEN_702 : tag_0_52; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2239 = ~quene ? _GEN_703 : tag_0_53; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2240 = ~quene ? _GEN_704 : tag_0_54; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2241 = ~quene ? _GEN_705 : tag_0_55; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2242 = ~quene ? _GEN_706 : tag_0_56; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2243 = ~quene ? _GEN_707 : tag_0_57; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2244 = ~quene ? _GEN_708 : tag_0_58; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2245 = ~quene ? _GEN_709 : tag_0_59; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2246 = ~quene ? _GEN_710 : tag_0_60; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2247 = ~quene ? _GEN_711 : tag_0_61; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2248 = ~quene ? _GEN_712 : tag_0_62; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2249 = ~quene ? _GEN_713 : tag_0_63; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2250 = ~quene ? _GEN_714 : tag_0_64; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2251 = ~quene ? _GEN_715 : tag_0_65; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2252 = ~quene ? _GEN_716 : tag_0_66; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2253 = ~quene ? _GEN_717 : tag_0_67; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2254 = ~quene ? _GEN_718 : tag_0_68; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2255 = ~quene ? _GEN_719 : tag_0_69; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2256 = ~quene ? _GEN_720 : tag_0_70; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2257 = ~quene ? _GEN_721 : tag_0_71; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2258 = ~quene ? _GEN_722 : tag_0_72; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2259 = ~quene ? _GEN_723 : tag_0_73; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2260 = ~quene ? _GEN_724 : tag_0_74; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2261 = ~quene ? _GEN_725 : tag_0_75; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2262 = ~quene ? _GEN_726 : tag_0_76; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2263 = ~quene ? _GEN_727 : tag_0_77; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2264 = ~quene ? _GEN_728 : tag_0_78; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2265 = ~quene ? _GEN_729 : tag_0_79; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2266 = ~quene ? _GEN_730 : tag_0_80; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2267 = ~quene ? _GEN_731 : tag_0_81; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2268 = ~quene ? _GEN_732 : tag_0_82; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2269 = ~quene ? _GEN_733 : tag_0_83; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2270 = ~quene ? _GEN_734 : tag_0_84; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2271 = ~quene ? _GEN_735 : tag_0_85; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2272 = ~quene ? _GEN_736 : tag_0_86; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2273 = ~quene ? _GEN_737 : tag_0_87; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2274 = ~quene ? _GEN_738 : tag_0_88; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2275 = ~quene ? _GEN_739 : tag_0_89; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2276 = ~quene ? _GEN_740 : tag_0_90; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2277 = ~quene ? _GEN_741 : tag_0_91; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2278 = ~quene ? _GEN_742 : tag_0_92; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2279 = ~quene ? _GEN_743 : tag_0_93; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2280 = ~quene ? _GEN_744 : tag_0_94; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2281 = ~quene ? _GEN_745 : tag_0_95; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2282 = ~quene ? _GEN_746 : tag_0_96; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2283 = ~quene ? _GEN_747 : tag_0_97; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2284 = ~quene ? _GEN_748 : tag_0_98; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2285 = ~quene ? _GEN_749 : tag_0_99; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2286 = ~quene ? _GEN_750 : tag_0_100; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2287 = ~quene ? _GEN_751 : tag_0_101; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2288 = ~quene ? _GEN_752 : tag_0_102; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2289 = ~quene ? _GEN_753 : tag_0_103; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2290 = ~quene ? _GEN_754 : tag_0_104; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2291 = ~quene ? _GEN_755 : tag_0_105; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2292 = ~quene ? _GEN_756 : tag_0_106; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2293 = ~quene ? _GEN_757 : tag_0_107; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2294 = ~quene ? _GEN_758 : tag_0_108; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2295 = ~quene ? _GEN_759 : tag_0_109; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2296 = ~quene ? _GEN_760 : tag_0_110; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2297 = ~quene ? _GEN_761 : tag_0_111; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2298 = ~quene ? _GEN_762 : tag_0_112; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2299 = ~quene ? _GEN_763 : tag_0_113; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2300 = ~quene ? _GEN_764 : tag_0_114; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2301 = ~quene ? _GEN_765 : tag_0_115; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2302 = ~quene ? _GEN_766 : tag_0_116; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2303 = ~quene ? _GEN_767 : tag_0_117; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2304 = ~quene ? _GEN_768 : tag_0_118; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2305 = ~quene ? _GEN_769 : tag_0_119; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2306 = ~quene ? _GEN_770 : tag_0_120; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2307 = ~quene ? _GEN_771 : tag_0_121; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2308 = ~quene ? _GEN_772 : tag_0_122; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2309 = ~quene ? _GEN_773 : tag_0_123; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2310 = ~quene ? _GEN_774 : tag_0_124; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2311 = ~quene ? _GEN_775 : tag_0_125; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2312 = ~quene ? _GEN_776 : tag_0_126; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2313 = ~quene ? _GEN_777 : tag_0_127; // @[i_cache.scala 19:24 97:34]
  wire  _GEN_2314 = ~quene ? _GEN_778 : valid_0_0; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2315 = ~quene ? _GEN_779 : valid_0_1; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2316 = ~quene ? _GEN_780 : valid_0_2; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2317 = ~quene ? _GEN_781 : valid_0_3; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2318 = ~quene ? _GEN_782 : valid_0_4; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2319 = ~quene ? _GEN_783 : valid_0_5; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2320 = ~quene ? _GEN_784 : valid_0_6; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2321 = ~quene ? _GEN_785 : valid_0_7; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2322 = ~quene ? _GEN_786 : valid_0_8; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2323 = ~quene ? _GEN_787 : valid_0_9; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2324 = ~quene ? _GEN_788 : valid_0_10; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2325 = ~quene ? _GEN_789 : valid_0_11; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2326 = ~quene ? _GEN_790 : valid_0_12; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2327 = ~quene ? _GEN_791 : valid_0_13; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2328 = ~quene ? _GEN_792 : valid_0_14; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2329 = ~quene ? _GEN_793 : valid_0_15; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2330 = ~quene ? _GEN_794 : valid_0_16; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2331 = ~quene ? _GEN_795 : valid_0_17; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2332 = ~quene ? _GEN_796 : valid_0_18; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2333 = ~quene ? _GEN_797 : valid_0_19; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2334 = ~quene ? _GEN_798 : valid_0_20; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2335 = ~quene ? _GEN_799 : valid_0_21; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2336 = ~quene ? _GEN_800 : valid_0_22; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2337 = ~quene ? _GEN_801 : valid_0_23; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2338 = ~quene ? _GEN_802 : valid_0_24; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2339 = ~quene ? _GEN_803 : valid_0_25; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2340 = ~quene ? _GEN_804 : valid_0_26; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2341 = ~quene ? _GEN_805 : valid_0_27; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2342 = ~quene ? _GEN_806 : valid_0_28; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2343 = ~quene ? _GEN_807 : valid_0_29; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2344 = ~quene ? _GEN_808 : valid_0_30; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2345 = ~quene ? _GEN_809 : valid_0_31; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2346 = ~quene ? _GEN_810 : valid_0_32; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2347 = ~quene ? _GEN_811 : valid_0_33; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2348 = ~quene ? _GEN_812 : valid_0_34; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2349 = ~quene ? _GEN_813 : valid_0_35; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2350 = ~quene ? _GEN_814 : valid_0_36; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2351 = ~quene ? _GEN_815 : valid_0_37; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2352 = ~quene ? _GEN_816 : valid_0_38; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2353 = ~quene ? _GEN_817 : valid_0_39; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2354 = ~quene ? _GEN_818 : valid_0_40; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2355 = ~quene ? _GEN_819 : valid_0_41; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2356 = ~quene ? _GEN_820 : valid_0_42; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2357 = ~quene ? _GEN_821 : valid_0_43; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2358 = ~quene ? _GEN_822 : valid_0_44; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2359 = ~quene ? _GEN_823 : valid_0_45; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2360 = ~quene ? _GEN_824 : valid_0_46; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2361 = ~quene ? _GEN_825 : valid_0_47; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2362 = ~quene ? _GEN_826 : valid_0_48; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2363 = ~quene ? _GEN_827 : valid_0_49; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2364 = ~quene ? _GEN_828 : valid_0_50; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2365 = ~quene ? _GEN_829 : valid_0_51; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2366 = ~quene ? _GEN_830 : valid_0_52; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2367 = ~quene ? _GEN_831 : valid_0_53; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2368 = ~quene ? _GEN_832 : valid_0_54; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2369 = ~quene ? _GEN_833 : valid_0_55; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2370 = ~quene ? _GEN_834 : valid_0_56; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2371 = ~quene ? _GEN_835 : valid_0_57; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2372 = ~quene ? _GEN_836 : valid_0_58; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2373 = ~quene ? _GEN_837 : valid_0_59; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2374 = ~quene ? _GEN_838 : valid_0_60; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2375 = ~quene ? _GEN_839 : valid_0_61; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2376 = ~quene ? _GEN_840 : valid_0_62; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2377 = ~quene ? _GEN_841 : valid_0_63; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2378 = ~quene ? _GEN_842 : valid_0_64; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2379 = ~quene ? _GEN_843 : valid_0_65; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2380 = ~quene ? _GEN_844 : valid_0_66; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2381 = ~quene ? _GEN_845 : valid_0_67; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2382 = ~quene ? _GEN_846 : valid_0_68; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2383 = ~quene ? _GEN_847 : valid_0_69; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2384 = ~quene ? _GEN_848 : valid_0_70; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2385 = ~quene ? _GEN_849 : valid_0_71; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2386 = ~quene ? _GEN_850 : valid_0_72; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2387 = ~quene ? _GEN_851 : valid_0_73; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2388 = ~quene ? _GEN_852 : valid_0_74; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2389 = ~quene ? _GEN_853 : valid_0_75; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2390 = ~quene ? _GEN_854 : valid_0_76; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2391 = ~quene ? _GEN_855 : valid_0_77; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2392 = ~quene ? _GEN_856 : valid_0_78; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2393 = ~quene ? _GEN_857 : valid_0_79; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2394 = ~quene ? _GEN_858 : valid_0_80; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2395 = ~quene ? _GEN_859 : valid_0_81; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2396 = ~quene ? _GEN_860 : valid_0_82; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2397 = ~quene ? _GEN_861 : valid_0_83; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2398 = ~quene ? _GEN_862 : valid_0_84; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2399 = ~quene ? _GEN_863 : valid_0_85; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2400 = ~quene ? _GEN_864 : valid_0_86; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2401 = ~quene ? _GEN_865 : valid_0_87; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2402 = ~quene ? _GEN_866 : valid_0_88; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2403 = ~quene ? _GEN_867 : valid_0_89; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2404 = ~quene ? _GEN_868 : valid_0_90; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2405 = ~quene ? _GEN_869 : valid_0_91; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2406 = ~quene ? _GEN_870 : valid_0_92; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2407 = ~quene ? _GEN_871 : valid_0_93; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2408 = ~quene ? _GEN_872 : valid_0_94; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2409 = ~quene ? _GEN_873 : valid_0_95; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2410 = ~quene ? _GEN_874 : valid_0_96; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2411 = ~quene ? _GEN_875 : valid_0_97; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2412 = ~quene ? _GEN_876 : valid_0_98; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2413 = ~quene ? _GEN_877 : valid_0_99; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2414 = ~quene ? _GEN_878 : valid_0_100; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2415 = ~quene ? _GEN_879 : valid_0_101; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2416 = ~quene ? _GEN_880 : valid_0_102; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2417 = ~quene ? _GEN_881 : valid_0_103; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2418 = ~quene ? _GEN_882 : valid_0_104; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2419 = ~quene ? _GEN_883 : valid_0_105; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2420 = ~quene ? _GEN_884 : valid_0_106; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2421 = ~quene ? _GEN_885 : valid_0_107; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2422 = ~quene ? _GEN_886 : valid_0_108; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2423 = ~quene ? _GEN_887 : valid_0_109; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2424 = ~quene ? _GEN_888 : valid_0_110; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2425 = ~quene ? _GEN_889 : valid_0_111; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2426 = ~quene ? _GEN_890 : valid_0_112; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2427 = ~quene ? _GEN_891 : valid_0_113; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2428 = ~quene ? _GEN_892 : valid_0_114; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2429 = ~quene ? _GEN_893 : valid_0_115; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2430 = ~quene ? _GEN_894 : valid_0_116; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2431 = ~quene ? _GEN_895 : valid_0_117; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2432 = ~quene ? _GEN_896 : valid_0_118; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2433 = ~quene ? _GEN_897 : valid_0_119; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2434 = ~quene ? _GEN_898 : valid_0_120; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2435 = ~quene ? _GEN_899 : valid_0_121; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2436 = ~quene ? _GEN_900 : valid_0_122; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2437 = ~quene ? _GEN_901 : valid_0_123; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2438 = ~quene ? _GEN_902 : valid_0_124; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2439 = ~quene ? _GEN_903 : valid_0_125; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2440 = ~quene ? _GEN_904 : valid_0_126; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2441 = ~quene ? _GEN_905 : valid_0_127; // @[i_cache.scala 21:26 97:34]
  wire [63:0] _GEN_2443 = ~quene ? ram_1_0 : _GEN_906; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2444 = ~quene ? ram_1_1 : _GEN_907; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2445 = ~quene ? ram_1_2 : _GEN_908; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2446 = ~quene ? ram_1_3 : _GEN_909; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2447 = ~quene ? ram_1_4 : _GEN_910; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2448 = ~quene ? ram_1_5 : _GEN_911; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2449 = ~quene ? ram_1_6 : _GEN_912; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2450 = ~quene ? ram_1_7 : _GEN_913; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2451 = ~quene ? ram_1_8 : _GEN_914; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2452 = ~quene ? ram_1_9 : _GEN_915; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2453 = ~quene ? ram_1_10 : _GEN_916; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2454 = ~quene ? ram_1_11 : _GEN_917; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2455 = ~quene ? ram_1_12 : _GEN_918; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2456 = ~quene ? ram_1_13 : _GEN_919; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2457 = ~quene ? ram_1_14 : _GEN_920; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2458 = ~quene ? ram_1_15 : _GEN_921; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2459 = ~quene ? ram_1_16 : _GEN_922; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2460 = ~quene ? ram_1_17 : _GEN_923; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2461 = ~quene ? ram_1_18 : _GEN_924; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2462 = ~quene ? ram_1_19 : _GEN_925; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2463 = ~quene ? ram_1_20 : _GEN_926; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2464 = ~quene ? ram_1_21 : _GEN_927; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2465 = ~quene ? ram_1_22 : _GEN_928; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2466 = ~quene ? ram_1_23 : _GEN_929; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2467 = ~quene ? ram_1_24 : _GEN_930; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2468 = ~quene ? ram_1_25 : _GEN_931; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2469 = ~quene ? ram_1_26 : _GEN_932; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2470 = ~quene ? ram_1_27 : _GEN_933; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2471 = ~quene ? ram_1_28 : _GEN_934; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2472 = ~quene ? ram_1_29 : _GEN_935; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2473 = ~quene ? ram_1_30 : _GEN_936; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2474 = ~quene ? ram_1_31 : _GEN_937; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2475 = ~quene ? ram_1_32 : _GEN_938; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2476 = ~quene ? ram_1_33 : _GEN_939; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2477 = ~quene ? ram_1_34 : _GEN_940; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2478 = ~quene ? ram_1_35 : _GEN_941; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2479 = ~quene ? ram_1_36 : _GEN_942; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2480 = ~quene ? ram_1_37 : _GEN_943; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2481 = ~quene ? ram_1_38 : _GEN_944; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2482 = ~quene ? ram_1_39 : _GEN_945; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2483 = ~quene ? ram_1_40 : _GEN_946; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2484 = ~quene ? ram_1_41 : _GEN_947; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2485 = ~quene ? ram_1_42 : _GEN_948; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2486 = ~quene ? ram_1_43 : _GEN_949; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2487 = ~quene ? ram_1_44 : _GEN_950; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2488 = ~quene ? ram_1_45 : _GEN_951; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2489 = ~quene ? ram_1_46 : _GEN_952; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2490 = ~quene ? ram_1_47 : _GEN_953; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2491 = ~quene ? ram_1_48 : _GEN_954; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2492 = ~quene ? ram_1_49 : _GEN_955; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2493 = ~quene ? ram_1_50 : _GEN_956; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2494 = ~quene ? ram_1_51 : _GEN_957; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2495 = ~quene ? ram_1_52 : _GEN_958; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2496 = ~quene ? ram_1_53 : _GEN_959; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2497 = ~quene ? ram_1_54 : _GEN_960; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2498 = ~quene ? ram_1_55 : _GEN_961; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2499 = ~quene ? ram_1_56 : _GEN_962; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2500 = ~quene ? ram_1_57 : _GEN_963; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2501 = ~quene ? ram_1_58 : _GEN_964; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2502 = ~quene ? ram_1_59 : _GEN_965; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2503 = ~quene ? ram_1_60 : _GEN_966; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2504 = ~quene ? ram_1_61 : _GEN_967; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2505 = ~quene ? ram_1_62 : _GEN_968; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2506 = ~quene ? ram_1_63 : _GEN_969; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2507 = ~quene ? ram_1_64 : _GEN_970; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2508 = ~quene ? ram_1_65 : _GEN_971; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2509 = ~quene ? ram_1_66 : _GEN_972; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2510 = ~quene ? ram_1_67 : _GEN_973; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2511 = ~quene ? ram_1_68 : _GEN_974; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2512 = ~quene ? ram_1_69 : _GEN_975; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2513 = ~quene ? ram_1_70 : _GEN_976; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2514 = ~quene ? ram_1_71 : _GEN_977; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2515 = ~quene ? ram_1_72 : _GEN_978; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2516 = ~quene ? ram_1_73 : _GEN_979; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2517 = ~quene ? ram_1_74 : _GEN_980; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2518 = ~quene ? ram_1_75 : _GEN_981; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2519 = ~quene ? ram_1_76 : _GEN_982; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2520 = ~quene ? ram_1_77 : _GEN_983; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2521 = ~quene ? ram_1_78 : _GEN_984; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2522 = ~quene ? ram_1_79 : _GEN_985; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2523 = ~quene ? ram_1_80 : _GEN_986; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2524 = ~quene ? ram_1_81 : _GEN_987; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2525 = ~quene ? ram_1_82 : _GEN_988; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2526 = ~quene ? ram_1_83 : _GEN_989; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2527 = ~quene ? ram_1_84 : _GEN_990; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2528 = ~quene ? ram_1_85 : _GEN_991; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2529 = ~quene ? ram_1_86 : _GEN_992; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2530 = ~quene ? ram_1_87 : _GEN_993; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2531 = ~quene ? ram_1_88 : _GEN_994; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2532 = ~quene ? ram_1_89 : _GEN_995; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2533 = ~quene ? ram_1_90 : _GEN_996; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2534 = ~quene ? ram_1_91 : _GEN_997; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2535 = ~quene ? ram_1_92 : _GEN_998; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2536 = ~quene ? ram_1_93 : _GEN_999; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2537 = ~quene ? ram_1_94 : _GEN_1000; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2538 = ~quene ? ram_1_95 : _GEN_1001; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2539 = ~quene ? ram_1_96 : _GEN_1002; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2540 = ~quene ? ram_1_97 : _GEN_1003; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2541 = ~quene ? ram_1_98 : _GEN_1004; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2542 = ~quene ? ram_1_99 : _GEN_1005; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2543 = ~quene ? ram_1_100 : _GEN_1006; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2544 = ~quene ? ram_1_101 : _GEN_1007; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2545 = ~quene ? ram_1_102 : _GEN_1008; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2546 = ~quene ? ram_1_103 : _GEN_1009; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2547 = ~quene ? ram_1_104 : _GEN_1010; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2548 = ~quene ? ram_1_105 : _GEN_1011; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2549 = ~quene ? ram_1_106 : _GEN_1012; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2550 = ~quene ? ram_1_107 : _GEN_1013; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2551 = ~quene ? ram_1_108 : _GEN_1014; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2552 = ~quene ? ram_1_109 : _GEN_1015; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2553 = ~quene ? ram_1_110 : _GEN_1016; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2554 = ~quene ? ram_1_111 : _GEN_1017; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2555 = ~quene ? ram_1_112 : _GEN_1018; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2556 = ~quene ? ram_1_113 : _GEN_1019; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2557 = ~quene ? ram_1_114 : _GEN_1020; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2558 = ~quene ? ram_1_115 : _GEN_1021; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2559 = ~quene ? ram_1_116 : _GEN_1022; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2560 = ~quene ? ram_1_117 : _GEN_1023; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2561 = ~quene ? ram_1_118 : _GEN_1024; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2562 = ~quene ? ram_1_119 : _GEN_1025; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2563 = ~quene ? ram_1_120 : _GEN_1026; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2564 = ~quene ? ram_1_121 : _GEN_1027; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2565 = ~quene ? ram_1_122 : _GEN_1028; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2566 = ~quene ? ram_1_123 : _GEN_1029; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2567 = ~quene ? ram_1_124 : _GEN_1030; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2568 = ~quene ? ram_1_125 : _GEN_1031; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2569 = ~quene ? ram_1_126 : _GEN_1032; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2570 = ~quene ? ram_1_127 : _GEN_1033; // @[i_cache.scala 18:24 97:34]
  wire [31:0] _GEN_2571 = ~quene ? tag_1_0 : _GEN_1034; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2572 = ~quene ? tag_1_1 : _GEN_1035; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2573 = ~quene ? tag_1_2 : _GEN_1036; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2574 = ~quene ? tag_1_3 : _GEN_1037; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2575 = ~quene ? tag_1_4 : _GEN_1038; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2576 = ~quene ? tag_1_5 : _GEN_1039; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2577 = ~quene ? tag_1_6 : _GEN_1040; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2578 = ~quene ? tag_1_7 : _GEN_1041; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2579 = ~quene ? tag_1_8 : _GEN_1042; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2580 = ~quene ? tag_1_9 : _GEN_1043; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2581 = ~quene ? tag_1_10 : _GEN_1044; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2582 = ~quene ? tag_1_11 : _GEN_1045; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2583 = ~quene ? tag_1_12 : _GEN_1046; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2584 = ~quene ? tag_1_13 : _GEN_1047; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2585 = ~quene ? tag_1_14 : _GEN_1048; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2586 = ~quene ? tag_1_15 : _GEN_1049; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2587 = ~quene ? tag_1_16 : _GEN_1050; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2588 = ~quene ? tag_1_17 : _GEN_1051; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2589 = ~quene ? tag_1_18 : _GEN_1052; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2590 = ~quene ? tag_1_19 : _GEN_1053; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2591 = ~quene ? tag_1_20 : _GEN_1054; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2592 = ~quene ? tag_1_21 : _GEN_1055; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2593 = ~quene ? tag_1_22 : _GEN_1056; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2594 = ~quene ? tag_1_23 : _GEN_1057; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2595 = ~quene ? tag_1_24 : _GEN_1058; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2596 = ~quene ? tag_1_25 : _GEN_1059; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2597 = ~quene ? tag_1_26 : _GEN_1060; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2598 = ~quene ? tag_1_27 : _GEN_1061; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2599 = ~quene ? tag_1_28 : _GEN_1062; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2600 = ~quene ? tag_1_29 : _GEN_1063; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2601 = ~quene ? tag_1_30 : _GEN_1064; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2602 = ~quene ? tag_1_31 : _GEN_1065; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2603 = ~quene ? tag_1_32 : _GEN_1066; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2604 = ~quene ? tag_1_33 : _GEN_1067; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2605 = ~quene ? tag_1_34 : _GEN_1068; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2606 = ~quene ? tag_1_35 : _GEN_1069; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2607 = ~quene ? tag_1_36 : _GEN_1070; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2608 = ~quene ? tag_1_37 : _GEN_1071; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2609 = ~quene ? tag_1_38 : _GEN_1072; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2610 = ~quene ? tag_1_39 : _GEN_1073; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2611 = ~quene ? tag_1_40 : _GEN_1074; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2612 = ~quene ? tag_1_41 : _GEN_1075; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2613 = ~quene ? tag_1_42 : _GEN_1076; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2614 = ~quene ? tag_1_43 : _GEN_1077; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2615 = ~quene ? tag_1_44 : _GEN_1078; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2616 = ~quene ? tag_1_45 : _GEN_1079; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2617 = ~quene ? tag_1_46 : _GEN_1080; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2618 = ~quene ? tag_1_47 : _GEN_1081; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2619 = ~quene ? tag_1_48 : _GEN_1082; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2620 = ~quene ? tag_1_49 : _GEN_1083; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2621 = ~quene ? tag_1_50 : _GEN_1084; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2622 = ~quene ? tag_1_51 : _GEN_1085; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2623 = ~quene ? tag_1_52 : _GEN_1086; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2624 = ~quene ? tag_1_53 : _GEN_1087; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2625 = ~quene ? tag_1_54 : _GEN_1088; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2626 = ~quene ? tag_1_55 : _GEN_1089; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2627 = ~quene ? tag_1_56 : _GEN_1090; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2628 = ~quene ? tag_1_57 : _GEN_1091; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2629 = ~quene ? tag_1_58 : _GEN_1092; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2630 = ~quene ? tag_1_59 : _GEN_1093; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2631 = ~quene ? tag_1_60 : _GEN_1094; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2632 = ~quene ? tag_1_61 : _GEN_1095; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2633 = ~quene ? tag_1_62 : _GEN_1096; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2634 = ~quene ? tag_1_63 : _GEN_1097; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2635 = ~quene ? tag_1_64 : _GEN_1098; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2636 = ~quene ? tag_1_65 : _GEN_1099; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2637 = ~quene ? tag_1_66 : _GEN_1100; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2638 = ~quene ? tag_1_67 : _GEN_1101; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2639 = ~quene ? tag_1_68 : _GEN_1102; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2640 = ~quene ? tag_1_69 : _GEN_1103; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2641 = ~quene ? tag_1_70 : _GEN_1104; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2642 = ~quene ? tag_1_71 : _GEN_1105; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2643 = ~quene ? tag_1_72 : _GEN_1106; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2644 = ~quene ? tag_1_73 : _GEN_1107; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2645 = ~quene ? tag_1_74 : _GEN_1108; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2646 = ~quene ? tag_1_75 : _GEN_1109; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2647 = ~quene ? tag_1_76 : _GEN_1110; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2648 = ~quene ? tag_1_77 : _GEN_1111; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2649 = ~quene ? tag_1_78 : _GEN_1112; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2650 = ~quene ? tag_1_79 : _GEN_1113; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2651 = ~quene ? tag_1_80 : _GEN_1114; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2652 = ~quene ? tag_1_81 : _GEN_1115; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2653 = ~quene ? tag_1_82 : _GEN_1116; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2654 = ~quene ? tag_1_83 : _GEN_1117; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2655 = ~quene ? tag_1_84 : _GEN_1118; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2656 = ~quene ? tag_1_85 : _GEN_1119; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2657 = ~quene ? tag_1_86 : _GEN_1120; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2658 = ~quene ? tag_1_87 : _GEN_1121; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2659 = ~quene ? tag_1_88 : _GEN_1122; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2660 = ~quene ? tag_1_89 : _GEN_1123; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2661 = ~quene ? tag_1_90 : _GEN_1124; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2662 = ~quene ? tag_1_91 : _GEN_1125; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2663 = ~quene ? tag_1_92 : _GEN_1126; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2664 = ~quene ? tag_1_93 : _GEN_1127; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2665 = ~quene ? tag_1_94 : _GEN_1128; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2666 = ~quene ? tag_1_95 : _GEN_1129; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2667 = ~quene ? tag_1_96 : _GEN_1130; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2668 = ~quene ? tag_1_97 : _GEN_1131; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2669 = ~quene ? tag_1_98 : _GEN_1132; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2670 = ~quene ? tag_1_99 : _GEN_1133; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2671 = ~quene ? tag_1_100 : _GEN_1134; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2672 = ~quene ? tag_1_101 : _GEN_1135; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2673 = ~quene ? tag_1_102 : _GEN_1136; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2674 = ~quene ? tag_1_103 : _GEN_1137; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2675 = ~quene ? tag_1_104 : _GEN_1138; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2676 = ~quene ? tag_1_105 : _GEN_1139; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2677 = ~quene ? tag_1_106 : _GEN_1140; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2678 = ~quene ? tag_1_107 : _GEN_1141; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2679 = ~quene ? tag_1_108 : _GEN_1142; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2680 = ~quene ? tag_1_109 : _GEN_1143; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2681 = ~quene ? tag_1_110 : _GEN_1144; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2682 = ~quene ? tag_1_111 : _GEN_1145; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2683 = ~quene ? tag_1_112 : _GEN_1146; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2684 = ~quene ? tag_1_113 : _GEN_1147; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2685 = ~quene ? tag_1_114 : _GEN_1148; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2686 = ~quene ? tag_1_115 : _GEN_1149; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2687 = ~quene ? tag_1_116 : _GEN_1150; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2688 = ~quene ? tag_1_117 : _GEN_1151; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2689 = ~quene ? tag_1_118 : _GEN_1152; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2690 = ~quene ? tag_1_119 : _GEN_1153; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2691 = ~quene ? tag_1_120 : _GEN_1154; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2692 = ~quene ? tag_1_121 : _GEN_1155; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2693 = ~quene ? tag_1_122 : _GEN_1156; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2694 = ~quene ? tag_1_123 : _GEN_1157; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2695 = ~quene ? tag_1_124 : _GEN_1158; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2696 = ~quene ? tag_1_125 : _GEN_1159; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2697 = ~quene ? tag_1_126 : _GEN_1160; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2698 = ~quene ? tag_1_127 : _GEN_1161; // @[i_cache.scala 20:24 97:34]
  wire  _GEN_2699 = ~quene ? valid_1_0 : _GEN_1162; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2700 = ~quene ? valid_1_1 : _GEN_1163; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2701 = ~quene ? valid_1_2 : _GEN_1164; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2702 = ~quene ? valid_1_3 : _GEN_1165; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2703 = ~quene ? valid_1_4 : _GEN_1166; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2704 = ~quene ? valid_1_5 : _GEN_1167; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2705 = ~quene ? valid_1_6 : _GEN_1168; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2706 = ~quene ? valid_1_7 : _GEN_1169; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2707 = ~quene ? valid_1_8 : _GEN_1170; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2708 = ~quene ? valid_1_9 : _GEN_1171; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2709 = ~quene ? valid_1_10 : _GEN_1172; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2710 = ~quene ? valid_1_11 : _GEN_1173; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2711 = ~quene ? valid_1_12 : _GEN_1174; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2712 = ~quene ? valid_1_13 : _GEN_1175; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2713 = ~quene ? valid_1_14 : _GEN_1176; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2714 = ~quene ? valid_1_15 : _GEN_1177; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2715 = ~quene ? valid_1_16 : _GEN_1178; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2716 = ~quene ? valid_1_17 : _GEN_1179; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2717 = ~quene ? valid_1_18 : _GEN_1180; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2718 = ~quene ? valid_1_19 : _GEN_1181; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2719 = ~quene ? valid_1_20 : _GEN_1182; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2720 = ~quene ? valid_1_21 : _GEN_1183; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2721 = ~quene ? valid_1_22 : _GEN_1184; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2722 = ~quene ? valid_1_23 : _GEN_1185; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2723 = ~quene ? valid_1_24 : _GEN_1186; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2724 = ~quene ? valid_1_25 : _GEN_1187; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2725 = ~quene ? valid_1_26 : _GEN_1188; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2726 = ~quene ? valid_1_27 : _GEN_1189; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2727 = ~quene ? valid_1_28 : _GEN_1190; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2728 = ~quene ? valid_1_29 : _GEN_1191; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2729 = ~quene ? valid_1_30 : _GEN_1192; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2730 = ~quene ? valid_1_31 : _GEN_1193; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2731 = ~quene ? valid_1_32 : _GEN_1194; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2732 = ~quene ? valid_1_33 : _GEN_1195; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2733 = ~quene ? valid_1_34 : _GEN_1196; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2734 = ~quene ? valid_1_35 : _GEN_1197; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2735 = ~quene ? valid_1_36 : _GEN_1198; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2736 = ~quene ? valid_1_37 : _GEN_1199; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2737 = ~quene ? valid_1_38 : _GEN_1200; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2738 = ~quene ? valid_1_39 : _GEN_1201; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2739 = ~quene ? valid_1_40 : _GEN_1202; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2740 = ~quene ? valid_1_41 : _GEN_1203; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2741 = ~quene ? valid_1_42 : _GEN_1204; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2742 = ~quene ? valid_1_43 : _GEN_1205; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2743 = ~quene ? valid_1_44 : _GEN_1206; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2744 = ~quene ? valid_1_45 : _GEN_1207; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2745 = ~quene ? valid_1_46 : _GEN_1208; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2746 = ~quene ? valid_1_47 : _GEN_1209; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2747 = ~quene ? valid_1_48 : _GEN_1210; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2748 = ~quene ? valid_1_49 : _GEN_1211; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2749 = ~quene ? valid_1_50 : _GEN_1212; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2750 = ~quene ? valid_1_51 : _GEN_1213; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2751 = ~quene ? valid_1_52 : _GEN_1214; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2752 = ~quene ? valid_1_53 : _GEN_1215; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2753 = ~quene ? valid_1_54 : _GEN_1216; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2754 = ~quene ? valid_1_55 : _GEN_1217; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2755 = ~quene ? valid_1_56 : _GEN_1218; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2756 = ~quene ? valid_1_57 : _GEN_1219; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2757 = ~quene ? valid_1_58 : _GEN_1220; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2758 = ~quene ? valid_1_59 : _GEN_1221; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2759 = ~quene ? valid_1_60 : _GEN_1222; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2760 = ~quene ? valid_1_61 : _GEN_1223; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2761 = ~quene ? valid_1_62 : _GEN_1224; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2762 = ~quene ? valid_1_63 : _GEN_1225; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2763 = ~quene ? valid_1_64 : _GEN_1226; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2764 = ~quene ? valid_1_65 : _GEN_1227; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2765 = ~quene ? valid_1_66 : _GEN_1228; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2766 = ~quene ? valid_1_67 : _GEN_1229; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2767 = ~quene ? valid_1_68 : _GEN_1230; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2768 = ~quene ? valid_1_69 : _GEN_1231; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2769 = ~quene ? valid_1_70 : _GEN_1232; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2770 = ~quene ? valid_1_71 : _GEN_1233; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2771 = ~quene ? valid_1_72 : _GEN_1234; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2772 = ~quene ? valid_1_73 : _GEN_1235; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2773 = ~quene ? valid_1_74 : _GEN_1236; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2774 = ~quene ? valid_1_75 : _GEN_1237; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2775 = ~quene ? valid_1_76 : _GEN_1238; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2776 = ~quene ? valid_1_77 : _GEN_1239; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2777 = ~quene ? valid_1_78 : _GEN_1240; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2778 = ~quene ? valid_1_79 : _GEN_1241; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2779 = ~quene ? valid_1_80 : _GEN_1242; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2780 = ~quene ? valid_1_81 : _GEN_1243; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2781 = ~quene ? valid_1_82 : _GEN_1244; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2782 = ~quene ? valid_1_83 : _GEN_1245; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2783 = ~quene ? valid_1_84 : _GEN_1246; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2784 = ~quene ? valid_1_85 : _GEN_1247; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2785 = ~quene ? valid_1_86 : _GEN_1248; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2786 = ~quene ? valid_1_87 : _GEN_1249; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2787 = ~quene ? valid_1_88 : _GEN_1250; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2788 = ~quene ? valid_1_89 : _GEN_1251; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2789 = ~quene ? valid_1_90 : _GEN_1252; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2790 = ~quene ? valid_1_91 : _GEN_1253; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2791 = ~quene ? valid_1_92 : _GEN_1254; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2792 = ~quene ? valid_1_93 : _GEN_1255; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2793 = ~quene ? valid_1_94 : _GEN_1256; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2794 = ~quene ? valid_1_95 : _GEN_1257; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2795 = ~quene ? valid_1_96 : _GEN_1258; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2796 = ~quene ? valid_1_97 : _GEN_1259; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2797 = ~quene ? valid_1_98 : _GEN_1260; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2798 = ~quene ? valid_1_99 : _GEN_1261; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2799 = ~quene ? valid_1_100 : _GEN_1262; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2800 = ~quene ? valid_1_101 : _GEN_1263; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2801 = ~quene ? valid_1_102 : _GEN_1264; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2802 = ~quene ? valid_1_103 : _GEN_1265; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2803 = ~quene ? valid_1_104 : _GEN_1266; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2804 = ~quene ? valid_1_105 : _GEN_1267; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2805 = ~quene ? valid_1_106 : _GEN_1268; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2806 = ~quene ? valid_1_107 : _GEN_1269; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2807 = ~quene ? valid_1_108 : _GEN_1270; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2808 = ~quene ? valid_1_109 : _GEN_1271; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2809 = ~quene ? valid_1_110 : _GEN_1272; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2810 = ~quene ? valid_1_111 : _GEN_1273; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2811 = ~quene ? valid_1_112 : _GEN_1274; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2812 = ~quene ? valid_1_113 : _GEN_1275; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2813 = ~quene ? valid_1_114 : _GEN_1276; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2814 = ~quene ? valid_1_115 : _GEN_1277; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2815 = ~quene ? valid_1_116 : _GEN_1278; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2816 = ~quene ? valid_1_117 : _GEN_1279; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2817 = ~quene ? valid_1_118 : _GEN_1280; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2818 = ~quene ? valid_1_119 : _GEN_1281; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2819 = ~quene ? valid_1_120 : _GEN_1282; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2820 = ~quene ? valid_1_121 : _GEN_1283; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2821 = ~quene ? valid_1_122 : _GEN_1284; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2822 = ~quene ? valid_1_123 : _GEN_1285; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2823 = ~quene ? valid_1_124 : _GEN_1286; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2824 = ~quene ? valid_1_125 : _GEN_1287; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2825 = ~quene ? valid_1_126 : _GEN_1288; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2826 = ~quene ? valid_1_127 : _GEN_1289; // @[i_cache.scala 22:26 97:34]
  wire [63:0] _GEN_2827 = unuse_way == 2'h2 ? _GEN_906 : _GEN_2443; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2828 = unuse_way == 2'h2 ? _GEN_907 : _GEN_2444; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2829 = unuse_way == 2'h2 ? _GEN_908 : _GEN_2445; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2830 = unuse_way == 2'h2 ? _GEN_909 : _GEN_2446; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2831 = unuse_way == 2'h2 ? _GEN_910 : _GEN_2447; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2832 = unuse_way == 2'h2 ? _GEN_911 : _GEN_2448; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2833 = unuse_way == 2'h2 ? _GEN_912 : _GEN_2449; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2834 = unuse_way == 2'h2 ? _GEN_913 : _GEN_2450; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2835 = unuse_way == 2'h2 ? _GEN_914 : _GEN_2451; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2836 = unuse_way == 2'h2 ? _GEN_915 : _GEN_2452; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2837 = unuse_way == 2'h2 ? _GEN_916 : _GEN_2453; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2838 = unuse_way == 2'h2 ? _GEN_917 : _GEN_2454; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2839 = unuse_way == 2'h2 ? _GEN_918 : _GEN_2455; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2840 = unuse_way == 2'h2 ? _GEN_919 : _GEN_2456; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2841 = unuse_way == 2'h2 ? _GEN_920 : _GEN_2457; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2842 = unuse_way == 2'h2 ? _GEN_921 : _GEN_2458; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2843 = unuse_way == 2'h2 ? _GEN_922 : _GEN_2459; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2844 = unuse_way == 2'h2 ? _GEN_923 : _GEN_2460; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2845 = unuse_way == 2'h2 ? _GEN_924 : _GEN_2461; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2846 = unuse_way == 2'h2 ? _GEN_925 : _GEN_2462; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2847 = unuse_way == 2'h2 ? _GEN_926 : _GEN_2463; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2848 = unuse_way == 2'h2 ? _GEN_927 : _GEN_2464; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2849 = unuse_way == 2'h2 ? _GEN_928 : _GEN_2465; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2850 = unuse_way == 2'h2 ? _GEN_929 : _GEN_2466; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2851 = unuse_way == 2'h2 ? _GEN_930 : _GEN_2467; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2852 = unuse_way == 2'h2 ? _GEN_931 : _GEN_2468; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2853 = unuse_way == 2'h2 ? _GEN_932 : _GEN_2469; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2854 = unuse_way == 2'h2 ? _GEN_933 : _GEN_2470; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2855 = unuse_way == 2'h2 ? _GEN_934 : _GEN_2471; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2856 = unuse_way == 2'h2 ? _GEN_935 : _GEN_2472; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2857 = unuse_way == 2'h2 ? _GEN_936 : _GEN_2473; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2858 = unuse_way == 2'h2 ? _GEN_937 : _GEN_2474; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2859 = unuse_way == 2'h2 ? _GEN_938 : _GEN_2475; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2860 = unuse_way == 2'h2 ? _GEN_939 : _GEN_2476; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2861 = unuse_way == 2'h2 ? _GEN_940 : _GEN_2477; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2862 = unuse_way == 2'h2 ? _GEN_941 : _GEN_2478; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2863 = unuse_way == 2'h2 ? _GEN_942 : _GEN_2479; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2864 = unuse_way == 2'h2 ? _GEN_943 : _GEN_2480; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2865 = unuse_way == 2'h2 ? _GEN_944 : _GEN_2481; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2866 = unuse_way == 2'h2 ? _GEN_945 : _GEN_2482; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2867 = unuse_way == 2'h2 ? _GEN_946 : _GEN_2483; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2868 = unuse_way == 2'h2 ? _GEN_947 : _GEN_2484; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2869 = unuse_way == 2'h2 ? _GEN_948 : _GEN_2485; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2870 = unuse_way == 2'h2 ? _GEN_949 : _GEN_2486; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2871 = unuse_way == 2'h2 ? _GEN_950 : _GEN_2487; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2872 = unuse_way == 2'h2 ? _GEN_951 : _GEN_2488; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2873 = unuse_way == 2'h2 ? _GEN_952 : _GEN_2489; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2874 = unuse_way == 2'h2 ? _GEN_953 : _GEN_2490; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2875 = unuse_way == 2'h2 ? _GEN_954 : _GEN_2491; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2876 = unuse_way == 2'h2 ? _GEN_955 : _GEN_2492; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2877 = unuse_way == 2'h2 ? _GEN_956 : _GEN_2493; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2878 = unuse_way == 2'h2 ? _GEN_957 : _GEN_2494; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2879 = unuse_way == 2'h2 ? _GEN_958 : _GEN_2495; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2880 = unuse_way == 2'h2 ? _GEN_959 : _GEN_2496; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2881 = unuse_way == 2'h2 ? _GEN_960 : _GEN_2497; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2882 = unuse_way == 2'h2 ? _GEN_961 : _GEN_2498; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2883 = unuse_way == 2'h2 ? _GEN_962 : _GEN_2499; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2884 = unuse_way == 2'h2 ? _GEN_963 : _GEN_2500; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2885 = unuse_way == 2'h2 ? _GEN_964 : _GEN_2501; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2886 = unuse_way == 2'h2 ? _GEN_965 : _GEN_2502; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2887 = unuse_way == 2'h2 ? _GEN_966 : _GEN_2503; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2888 = unuse_way == 2'h2 ? _GEN_967 : _GEN_2504; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2889 = unuse_way == 2'h2 ? _GEN_968 : _GEN_2505; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2890 = unuse_way == 2'h2 ? _GEN_969 : _GEN_2506; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2891 = unuse_way == 2'h2 ? _GEN_970 : _GEN_2507; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2892 = unuse_way == 2'h2 ? _GEN_971 : _GEN_2508; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2893 = unuse_way == 2'h2 ? _GEN_972 : _GEN_2509; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2894 = unuse_way == 2'h2 ? _GEN_973 : _GEN_2510; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2895 = unuse_way == 2'h2 ? _GEN_974 : _GEN_2511; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2896 = unuse_way == 2'h2 ? _GEN_975 : _GEN_2512; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2897 = unuse_way == 2'h2 ? _GEN_976 : _GEN_2513; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2898 = unuse_way == 2'h2 ? _GEN_977 : _GEN_2514; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2899 = unuse_way == 2'h2 ? _GEN_978 : _GEN_2515; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2900 = unuse_way == 2'h2 ? _GEN_979 : _GEN_2516; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2901 = unuse_way == 2'h2 ? _GEN_980 : _GEN_2517; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2902 = unuse_way == 2'h2 ? _GEN_981 : _GEN_2518; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2903 = unuse_way == 2'h2 ? _GEN_982 : _GEN_2519; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2904 = unuse_way == 2'h2 ? _GEN_983 : _GEN_2520; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2905 = unuse_way == 2'h2 ? _GEN_984 : _GEN_2521; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2906 = unuse_way == 2'h2 ? _GEN_985 : _GEN_2522; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2907 = unuse_way == 2'h2 ? _GEN_986 : _GEN_2523; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2908 = unuse_way == 2'h2 ? _GEN_987 : _GEN_2524; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2909 = unuse_way == 2'h2 ? _GEN_988 : _GEN_2525; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2910 = unuse_way == 2'h2 ? _GEN_989 : _GEN_2526; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2911 = unuse_way == 2'h2 ? _GEN_990 : _GEN_2527; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2912 = unuse_way == 2'h2 ? _GEN_991 : _GEN_2528; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2913 = unuse_way == 2'h2 ? _GEN_992 : _GEN_2529; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2914 = unuse_way == 2'h2 ? _GEN_993 : _GEN_2530; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2915 = unuse_way == 2'h2 ? _GEN_994 : _GEN_2531; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2916 = unuse_way == 2'h2 ? _GEN_995 : _GEN_2532; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2917 = unuse_way == 2'h2 ? _GEN_996 : _GEN_2533; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2918 = unuse_way == 2'h2 ? _GEN_997 : _GEN_2534; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2919 = unuse_way == 2'h2 ? _GEN_998 : _GEN_2535; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2920 = unuse_way == 2'h2 ? _GEN_999 : _GEN_2536; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2921 = unuse_way == 2'h2 ? _GEN_1000 : _GEN_2537; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2922 = unuse_way == 2'h2 ? _GEN_1001 : _GEN_2538; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2923 = unuse_way == 2'h2 ? _GEN_1002 : _GEN_2539; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2924 = unuse_way == 2'h2 ? _GEN_1003 : _GEN_2540; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2925 = unuse_way == 2'h2 ? _GEN_1004 : _GEN_2541; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2926 = unuse_way == 2'h2 ? _GEN_1005 : _GEN_2542; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2927 = unuse_way == 2'h2 ? _GEN_1006 : _GEN_2543; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2928 = unuse_way == 2'h2 ? _GEN_1007 : _GEN_2544; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2929 = unuse_way == 2'h2 ? _GEN_1008 : _GEN_2545; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2930 = unuse_way == 2'h2 ? _GEN_1009 : _GEN_2546; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2931 = unuse_way == 2'h2 ? _GEN_1010 : _GEN_2547; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2932 = unuse_way == 2'h2 ? _GEN_1011 : _GEN_2548; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2933 = unuse_way == 2'h2 ? _GEN_1012 : _GEN_2549; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2934 = unuse_way == 2'h2 ? _GEN_1013 : _GEN_2550; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2935 = unuse_way == 2'h2 ? _GEN_1014 : _GEN_2551; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2936 = unuse_way == 2'h2 ? _GEN_1015 : _GEN_2552; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2937 = unuse_way == 2'h2 ? _GEN_1016 : _GEN_2553; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2938 = unuse_way == 2'h2 ? _GEN_1017 : _GEN_2554; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2939 = unuse_way == 2'h2 ? _GEN_1018 : _GEN_2555; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2940 = unuse_way == 2'h2 ? _GEN_1019 : _GEN_2556; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2941 = unuse_way == 2'h2 ? _GEN_1020 : _GEN_2557; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2942 = unuse_way == 2'h2 ? _GEN_1021 : _GEN_2558; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2943 = unuse_way == 2'h2 ? _GEN_1022 : _GEN_2559; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2944 = unuse_way == 2'h2 ? _GEN_1023 : _GEN_2560; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2945 = unuse_way == 2'h2 ? _GEN_1024 : _GEN_2561; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2946 = unuse_way == 2'h2 ? _GEN_1025 : _GEN_2562; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2947 = unuse_way == 2'h2 ? _GEN_1026 : _GEN_2563; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2948 = unuse_way == 2'h2 ? _GEN_1027 : _GEN_2564; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2949 = unuse_way == 2'h2 ? _GEN_1028 : _GEN_2565; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2950 = unuse_way == 2'h2 ? _GEN_1029 : _GEN_2566; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2951 = unuse_way == 2'h2 ? _GEN_1030 : _GEN_2567; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2952 = unuse_way == 2'h2 ? _GEN_1031 : _GEN_2568; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2953 = unuse_way == 2'h2 ? _GEN_1032 : _GEN_2569; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2954 = unuse_way == 2'h2 ? _GEN_1033 : _GEN_2570; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2955 = unuse_way == 2'h2 ? _GEN_1034 : _GEN_2571; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2956 = unuse_way == 2'h2 ? _GEN_1035 : _GEN_2572; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2957 = unuse_way == 2'h2 ? _GEN_1036 : _GEN_2573; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2958 = unuse_way == 2'h2 ? _GEN_1037 : _GEN_2574; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2959 = unuse_way == 2'h2 ? _GEN_1038 : _GEN_2575; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2960 = unuse_way == 2'h2 ? _GEN_1039 : _GEN_2576; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2961 = unuse_way == 2'h2 ? _GEN_1040 : _GEN_2577; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2962 = unuse_way == 2'h2 ? _GEN_1041 : _GEN_2578; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2963 = unuse_way == 2'h2 ? _GEN_1042 : _GEN_2579; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2964 = unuse_way == 2'h2 ? _GEN_1043 : _GEN_2580; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2965 = unuse_way == 2'h2 ? _GEN_1044 : _GEN_2581; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2966 = unuse_way == 2'h2 ? _GEN_1045 : _GEN_2582; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2967 = unuse_way == 2'h2 ? _GEN_1046 : _GEN_2583; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2968 = unuse_way == 2'h2 ? _GEN_1047 : _GEN_2584; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2969 = unuse_way == 2'h2 ? _GEN_1048 : _GEN_2585; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2970 = unuse_way == 2'h2 ? _GEN_1049 : _GEN_2586; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2971 = unuse_way == 2'h2 ? _GEN_1050 : _GEN_2587; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2972 = unuse_way == 2'h2 ? _GEN_1051 : _GEN_2588; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2973 = unuse_way == 2'h2 ? _GEN_1052 : _GEN_2589; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2974 = unuse_way == 2'h2 ? _GEN_1053 : _GEN_2590; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2975 = unuse_way == 2'h2 ? _GEN_1054 : _GEN_2591; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2976 = unuse_way == 2'h2 ? _GEN_1055 : _GEN_2592; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2977 = unuse_way == 2'h2 ? _GEN_1056 : _GEN_2593; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2978 = unuse_way == 2'h2 ? _GEN_1057 : _GEN_2594; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2979 = unuse_way == 2'h2 ? _GEN_1058 : _GEN_2595; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2980 = unuse_way == 2'h2 ? _GEN_1059 : _GEN_2596; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2981 = unuse_way == 2'h2 ? _GEN_1060 : _GEN_2597; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2982 = unuse_way == 2'h2 ? _GEN_1061 : _GEN_2598; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2983 = unuse_way == 2'h2 ? _GEN_1062 : _GEN_2599; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2984 = unuse_way == 2'h2 ? _GEN_1063 : _GEN_2600; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2985 = unuse_way == 2'h2 ? _GEN_1064 : _GEN_2601; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2986 = unuse_way == 2'h2 ? _GEN_1065 : _GEN_2602; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2987 = unuse_way == 2'h2 ? _GEN_1066 : _GEN_2603; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2988 = unuse_way == 2'h2 ? _GEN_1067 : _GEN_2604; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2989 = unuse_way == 2'h2 ? _GEN_1068 : _GEN_2605; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2990 = unuse_way == 2'h2 ? _GEN_1069 : _GEN_2606; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2991 = unuse_way == 2'h2 ? _GEN_1070 : _GEN_2607; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2992 = unuse_way == 2'h2 ? _GEN_1071 : _GEN_2608; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2993 = unuse_way == 2'h2 ? _GEN_1072 : _GEN_2609; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2994 = unuse_way == 2'h2 ? _GEN_1073 : _GEN_2610; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2995 = unuse_way == 2'h2 ? _GEN_1074 : _GEN_2611; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2996 = unuse_way == 2'h2 ? _GEN_1075 : _GEN_2612; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2997 = unuse_way == 2'h2 ? _GEN_1076 : _GEN_2613; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2998 = unuse_way == 2'h2 ? _GEN_1077 : _GEN_2614; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2999 = unuse_way == 2'h2 ? _GEN_1078 : _GEN_2615; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3000 = unuse_way == 2'h2 ? _GEN_1079 : _GEN_2616; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3001 = unuse_way == 2'h2 ? _GEN_1080 : _GEN_2617; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3002 = unuse_way == 2'h2 ? _GEN_1081 : _GEN_2618; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3003 = unuse_way == 2'h2 ? _GEN_1082 : _GEN_2619; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3004 = unuse_way == 2'h2 ? _GEN_1083 : _GEN_2620; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3005 = unuse_way == 2'h2 ? _GEN_1084 : _GEN_2621; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3006 = unuse_way == 2'h2 ? _GEN_1085 : _GEN_2622; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3007 = unuse_way == 2'h2 ? _GEN_1086 : _GEN_2623; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3008 = unuse_way == 2'h2 ? _GEN_1087 : _GEN_2624; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3009 = unuse_way == 2'h2 ? _GEN_1088 : _GEN_2625; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3010 = unuse_way == 2'h2 ? _GEN_1089 : _GEN_2626; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3011 = unuse_way == 2'h2 ? _GEN_1090 : _GEN_2627; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3012 = unuse_way == 2'h2 ? _GEN_1091 : _GEN_2628; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3013 = unuse_way == 2'h2 ? _GEN_1092 : _GEN_2629; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3014 = unuse_way == 2'h2 ? _GEN_1093 : _GEN_2630; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3015 = unuse_way == 2'h2 ? _GEN_1094 : _GEN_2631; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3016 = unuse_way == 2'h2 ? _GEN_1095 : _GEN_2632; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3017 = unuse_way == 2'h2 ? _GEN_1096 : _GEN_2633; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3018 = unuse_way == 2'h2 ? _GEN_1097 : _GEN_2634; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3019 = unuse_way == 2'h2 ? _GEN_1098 : _GEN_2635; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3020 = unuse_way == 2'h2 ? _GEN_1099 : _GEN_2636; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3021 = unuse_way == 2'h2 ? _GEN_1100 : _GEN_2637; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3022 = unuse_way == 2'h2 ? _GEN_1101 : _GEN_2638; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3023 = unuse_way == 2'h2 ? _GEN_1102 : _GEN_2639; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3024 = unuse_way == 2'h2 ? _GEN_1103 : _GEN_2640; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3025 = unuse_way == 2'h2 ? _GEN_1104 : _GEN_2641; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3026 = unuse_way == 2'h2 ? _GEN_1105 : _GEN_2642; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3027 = unuse_way == 2'h2 ? _GEN_1106 : _GEN_2643; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3028 = unuse_way == 2'h2 ? _GEN_1107 : _GEN_2644; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3029 = unuse_way == 2'h2 ? _GEN_1108 : _GEN_2645; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3030 = unuse_way == 2'h2 ? _GEN_1109 : _GEN_2646; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3031 = unuse_way == 2'h2 ? _GEN_1110 : _GEN_2647; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3032 = unuse_way == 2'h2 ? _GEN_1111 : _GEN_2648; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3033 = unuse_way == 2'h2 ? _GEN_1112 : _GEN_2649; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3034 = unuse_way == 2'h2 ? _GEN_1113 : _GEN_2650; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3035 = unuse_way == 2'h2 ? _GEN_1114 : _GEN_2651; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3036 = unuse_way == 2'h2 ? _GEN_1115 : _GEN_2652; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3037 = unuse_way == 2'h2 ? _GEN_1116 : _GEN_2653; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3038 = unuse_way == 2'h2 ? _GEN_1117 : _GEN_2654; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3039 = unuse_way == 2'h2 ? _GEN_1118 : _GEN_2655; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3040 = unuse_way == 2'h2 ? _GEN_1119 : _GEN_2656; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3041 = unuse_way == 2'h2 ? _GEN_1120 : _GEN_2657; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3042 = unuse_way == 2'h2 ? _GEN_1121 : _GEN_2658; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3043 = unuse_way == 2'h2 ? _GEN_1122 : _GEN_2659; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3044 = unuse_way == 2'h2 ? _GEN_1123 : _GEN_2660; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3045 = unuse_way == 2'h2 ? _GEN_1124 : _GEN_2661; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3046 = unuse_way == 2'h2 ? _GEN_1125 : _GEN_2662; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3047 = unuse_way == 2'h2 ? _GEN_1126 : _GEN_2663; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3048 = unuse_way == 2'h2 ? _GEN_1127 : _GEN_2664; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3049 = unuse_way == 2'h2 ? _GEN_1128 : _GEN_2665; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3050 = unuse_way == 2'h2 ? _GEN_1129 : _GEN_2666; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3051 = unuse_way == 2'h2 ? _GEN_1130 : _GEN_2667; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3052 = unuse_way == 2'h2 ? _GEN_1131 : _GEN_2668; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3053 = unuse_way == 2'h2 ? _GEN_1132 : _GEN_2669; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3054 = unuse_way == 2'h2 ? _GEN_1133 : _GEN_2670; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3055 = unuse_way == 2'h2 ? _GEN_1134 : _GEN_2671; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3056 = unuse_way == 2'h2 ? _GEN_1135 : _GEN_2672; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3057 = unuse_way == 2'h2 ? _GEN_1136 : _GEN_2673; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3058 = unuse_way == 2'h2 ? _GEN_1137 : _GEN_2674; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3059 = unuse_way == 2'h2 ? _GEN_1138 : _GEN_2675; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3060 = unuse_way == 2'h2 ? _GEN_1139 : _GEN_2676; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3061 = unuse_way == 2'h2 ? _GEN_1140 : _GEN_2677; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3062 = unuse_way == 2'h2 ? _GEN_1141 : _GEN_2678; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3063 = unuse_way == 2'h2 ? _GEN_1142 : _GEN_2679; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3064 = unuse_way == 2'h2 ? _GEN_1143 : _GEN_2680; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3065 = unuse_way == 2'h2 ? _GEN_1144 : _GEN_2681; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3066 = unuse_way == 2'h2 ? _GEN_1145 : _GEN_2682; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3067 = unuse_way == 2'h2 ? _GEN_1146 : _GEN_2683; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3068 = unuse_way == 2'h2 ? _GEN_1147 : _GEN_2684; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3069 = unuse_way == 2'h2 ? _GEN_1148 : _GEN_2685; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3070 = unuse_way == 2'h2 ? _GEN_1149 : _GEN_2686; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3071 = unuse_way == 2'h2 ? _GEN_1150 : _GEN_2687; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3072 = unuse_way == 2'h2 ? _GEN_1151 : _GEN_2688; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3073 = unuse_way == 2'h2 ? _GEN_1152 : _GEN_2689; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3074 = unuse_way == 2'h2 ? _GEN_1153 : _GEN_2690; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3075 = unuse_way == 2'h2 ? _GEN_1154 : _GEN_2691; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3076 = unuse_way == 2'h2 ? _GEN_1155 : _GEN_2692; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3077 = unuse_way == 2'h2 ? _GEN_1156 : _GEN_2693; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3078 = unuse_way == 2'h2 ? _GEN_1157 : _GEN_2694; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3079 = unuse_way == 2'h2 ? _GEN_1158 : _GEN_2695; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3080 = unuse_way == 2'h2 ? _GEN_1159 : _GEN_2696; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3081 = unuse_way == 2'h2 ? _GEN_1160 : _GEN_2697; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3082 = unuse_way == 2'h2 ? _GEN_1161 : _GEN_2698; // @[i_cache.scala 91:40]
  wire  _GEN_3083 = unuse_way == 2'h2 ? _GEN_1162 : _GEN_2699; // @[i_cache.scala 91:40]
  wire  _GEN_3084 = unuse_way == 2'h2 ? _GEN_1163 : _GEN_2700; // @[i_cache.scala 91:40]
  wire  _GEN_3085 = unuse_way == 2'h2 ? _GEN_1164 : _GEN_2701; // @[i_cache.scala 91:40]
  wire  _GEN_3086 = unuse_way == 2'h2 ? _GEN_1165 : _GEN_2702; // @[i_cache.scala 91:40]
  wire  _GEN_3087 = unuse_way == 2'h2 ? _GEN_1166 : _GEN_2703; // @[i_cache.scala 91:40]
  wire  _GEN_3088 = unuse_way == 2'h2 ? _GEN_1167 : _GEN_2704; // @[i_cache.scala 91:40]
  wire  _GEN_3089 = unuse_way == 2'h2 ? _GEN_1168 : _GEN_2705; // @[i_cache.scala 91:40]
  wire  _GEN_3090 = unuse_way == 2'h2 ? _GEN_1169 : _GEN_2706; // @[i_cache.scala 91:40]
  wire  _GEN_3091 = unuse_way == 2'h2 ? _GEN_1170 : _GEN_2707; // @[i_cache.scala 91:40]
  wire  _GEN_3092 = unuse_way == 2'h2 ? _GEN_1171 : _GEN_2708; // @[i_cache.scala 91:40]
  wire  _GEN_3093 = unuse_way == 2'h2 ? _GEN_1172 : _GEN_2709; // @[i_cache.scala 91:40]
  wire  _GEN_3094 = unuse_way == 2'h2 ? _GEN_1173 : _GEN_2710; // @[i_cache.scala 91:40]
  wire  _GEN_3095 = unuse_way == 2'h2 ? _GEN_1174 : _GEN_2711; // @[i_cache.scala 91:40]
  wire  _GEN_3096 = unuse_way == 2'h2 ? _GEN_1175 : _GEN_2712; // @[i_cache.scala 91:40]
  wire  _GEN_3097 = unuse_way == 2'h2 ? _GEN_1176 : _GEN_2713; // @[i_cache.scala 91:40]
  wire  _GEN_3098 = unuse_way == 2'h2 ? _GEN_1177 : _GEN_2714; // @[i_cache.scala 91:40]
  wire  _GEN_3099 = unuse_way == 2'h2 ? _GEN_1178 : _GEN_2715; // @[i_cache.scala 91:40]
  wire  _GEN_3100 = unuse_way == 2'h2 ? _GEN_1179 : _GEN_2716; // @[i_cache.scala 91:40]
  wire  _GEN_3101 = unuse_way == 2'h2 ? _GEN_1180 : _GEN_2717; // @[i_cache.scala 91:40]
  wire  _GEN_3102 = unuse_way == 2'h2 ? _GEN_1181 : _GEN_2718; // @[i_cache.scala 91:40]
  wire  _GEN_3103 = unuse_way == 2'h2 ? _GEN_1182 : _GEN_2719; // @[i_cache.scala 91:40]
  wire  _GEN_3104 = unuse_way == 2'h2 ? _GEN_1183 : _GEN_2720; // @[i_cache.scala 91:40]
  wire  _GEN_3105 = unuse_way == 2'h2 ? _GEN_1184 : _GEN_2721; // @[i_cache.scala 91:40]
  wire  _GEN_3106 = unuse_way == 2'h2 ? _GEN_1185 : _GEN_2722; // @[i_cache.scala 91:40]
  wire  _GEN_3107 = unuse_way == 2'h2 ? _GEN_1186 : _GEN_2723; // @[i_cache.scala 91:40]
  wire  _GEN_3108 = unuse_way == 2'h2 ? _GEN_1187 : _GEN_2724; // @[i_cache.scala 91:40]
  wire  _GEN_3109 = unuse_way == 2'h2 ? _GEN_1188 : _GEN_2725; // @[i_cache.scala 91:40]
  wire  _GEN_3110 = unuse_way == 2'h2 ? _GEN_1189 : _GEN_2726; // @[i_cache.scala 91:40]
  wire  _GEN_3111 = unuse_way == 2'h2 ? _GEN_1190 : _GEN_2727; // @[i_cache.scala 91:40]
  wire  _GEN_3112 = unuse_way == 2'h2 ? _GEN_1191 : _GEN_2728; // @[i_cache.scala 91:40]
  wire  _GEN_3113 = unuse_way == 2'h2 ? _GEN_1192 : _GEN_2729; // @[i_cache.scala 91:40]
  wire  _GEN_3114 = unuse_way == 2'h2 ? _GEN_1193 : _GEN_2730; // @[i_cache.scala 91:40]
  wire  _GEN_3115 = unuse_way == 2'h2 ? _GEN_1194 : _GEN_2731; // @[i_cache.scala 91:40]
  wire  _GEN_3116 = unuse_way == 2'h2 ? _GEN_1195 : _GEN_2732; // @[i_cache.scala 91:40]
  wire  _GEN_3117 = unuse_way == 2'h2 ? _GEN_1196 : _GEN_2733; // @[i_cache.scala 91:40]
  wire  _GEN_3118 = unuse_way == 2'h2 ? _GEN_1197 : _GEN_2734; // @[i_cache.scala 91:40]
  wire  _GEN_3119 = unuse_way == 2'h2 ? _GEN_1198 : _GEN_2735; // @[i_cache.scala 91:40]
  wire  _GEN_3120 = unuse_way == 2'h2 ? _GEN_1199 : _GEN_2736; // @[i_cache.scala 91:40]
  wire  _GEN_3121 = unuse_way == 2'h2 ? _GEN_1200 : _GEN_2737; // @[i_cache.scala 91:40]
  wire  _GEN_3122 = unuse_way == 2'h2 ? _GEN_1201 : _GEN_2738; // @[i_cache.scala 91:40]
  wire  _GEN_3123 = unuse_way == 2'h2 ? _GEN_1202 : _GEN_2739; // @[i_cache.scala 91:40]
  wire  _GEN_3124 = unuse_way == 2'h2 ? _GEN_1203 : _GEN_2740; // @[i_cache.scala 91:40]
  wire  _GEN_3125 = unuse_way == 2'h2 ? _GEN_1204 : _GEN_2741; // @[i_cache.scala 91:40]
  wire  _GEN_3126 = unuse_way == 2'h2 ? _GEN_1205 : _GEN_2742; // @[i_cache.scala 91:40]
  wire  _GEN_3127 = unuse_way == 2'h2 ? _GEN_1206 : _GEN_2743; // @[i_cache.scala 91:40]
  wire  _GEN_3128 = unuse_way == 2'h2 ? _GEN_1207 : _GEN_2744; // @[i_cache.scala 91:40]
  wire  _GEN_3129 = unuse_way == 2'h2 ? _GEN_1208 : _GEN_2745; // @[i_cache.scala 91:40]
  wire  _GEN_3130 = unuse_way == 2'h2 ? _GEN_1209 : _GEN_2746; // @[i_cache.scala 91:40]
  wire  _GEN_3131 = unuse_way == 2'h2 ? _GEN_1210 : _GEN_2747; // @[i_cache.scala 91:40]
  wire  _GEN_3132 = unuse_way == 2'h2 ? _GEN_1211 : _GEN_2748; // @[i_cache.scala 91:40]
  wire  _GEN_3133 = unuse_way == 2'h2 ? _GEN_1212 : _GEN_2749; // @[i_cache.scala 91:40]
  wire  _GEN_3134 = unuse_way == 2'h2 ? _GEN_1213 : _GEN_2750; // @[i_cache.scala 91:40]
  wire  _GEN_3135 = unuse_way == 2'h2 ? _GEN_1214 : _GEN_2751; // @[i_cache.scala 91:40]
  wire  _GEN_3136 = unuse_way == 2'h2 ? _GEN_1215 : _GEN_2752; // @[i_cache.scala 91:40]
  wire  _GEN_3137 = unuse_way == 2'h2 ? _GEN_1216 : _GEN_2753; // @[i_cache.scala 91:40]
  wire  _GEN_3138 = unuse_way == 2'h2 ? _GEN_1217 : _GEN_2754; // @[i_cache.scala 91:40]
  wire  _GEN_3139 = unuse_way == 2'h2 ? _GEN_1218 : _GEN_2755; // @[i_cache.scala 91:40]
  wire  _GEN_3140 = unuse_way == 2'h2 ? _GEN_1219 : _GEN_2756; // @[i_cache.scala 91:40]
  wire  _GEN_3141 = unuse_way == 2'h2 ? _GEN_1220 : _GEN_2757; // @[i_cache.scala 91:40]
  wire  _GEN_3142 = unuse_way == 2'h2 ? _GEN_1221 : _GEN_2758; // @[i_cache.scala 91:40]
  wire  _GEN_3143 = unuse_way == 2'h2 ? _GEN_1222 : _GEN_2759; // @[i_cache.scala 91:40]
  wire  _GEN_3144 = unuse_way == 2'h2 ? _GEN_1223 : _GEN_2760; // @[i_cache.scala 91:40]
  wire  _GEN_3145 = unuse_way == 2'h2 ? _GEN_1224 : _GEN_2761; // @[i_cache.scala 91:40]
  wire  _GEN_3146 = unuse_way == 2'h2 ? _GEN_1225 : _GEN_2762; // @[i_cache.scala 91:40]
  wire  _GEN_3147 = unuse_way == 2'h2 ? _GEN_1226 : _GEN_2763; // @[i_cache.scala 91:40]
  wire  _GEN_3148 = unuse_way == 2'h2 ? _GEN_1227 : _GEN_2764; // @[i_cache.scala 91:40]
  wire  _GEN_3149 = unuse_way == 2'h2 ? _GEN_1228 : _GEN_2765; // @[i_cache.scala 91:40]
  wire  _GEN_3150 = unuse_way == 2'h2 ? _GEN_1229 : _GEN_2766; // @[i_cache.scala 91:40]
  wire  _GEN_3151 = unuse_way == 2'h2 ? _GEN_1230 : _GEN_2767; // @[i_cache.scala 91:40]
  wire  _GEN_3152 = unuse_way == 2'h2 ? _GEN_1231 : _GEN_2768; // @[i_cache.scala 91:40]
  wire  _GEN_3153 = unuse_way == 2'h2 ? _GEN_1232 : _GEN_2769; // @[i_cache.scala 91:40]
  wire  _GEN_3154 = unuse_way == 2'h2 ? _GEN_1233 : _GEN_2770; // @[i_cache.scala 91:40]
  wire  _GEN_3155 = unuse_way == 2'h2 ? _GEN_1234 : _GEN_2771; // @[i_cache.scala 91:40]
  wire  _GEN_3156 = unuse_way == 2'h2 ? _GEN_1235 : _GEN_2772; // @[i_cache.scala 91:40]
  wire  _GEN_3157 = unuse_way == 2'h2 ? _GEN_1236 : _GEN_2773; // @[i_cache.scala 91:40]
  wire  _GEN_3158 = unuse_way == 2'h2 ? _GEN_1237 : _GEN_2774; // @[i_cache.scala 91:40]
  wire  _GEN_3159 = unuse_way == 2'h2 ? _GEN_1238 : _GEN_2775; // @[i_cache.scala 91:40]
  wire  _GEN_3160 = unuse_way == 2'h2 ? _GEN_1239 : _GEN_2776; // @[i_cache.scala 91:40]
  wire  _GEN_3161 = unuse_way == 2'h2 ? _GEN_1240 : _GEN_2777; // @[i_cache.scala 91:40]
  wire  _GEN_3162 = unuse_way == 2'h2 ? _GEN_1241 : _GEN_2778; // @[i_cache.scala 91:40]
  wire  _GEN_3163 = unuse_way == 2'h2 ? _GEN_1242 : _GEN_2779; // @[i_cache.scala 91:40]
  wire  _GEN_3164 = unuse_way == 2'h2 ? _GEN_1243 : _GEN_2780; // @[i_cache.scala 91:40]
  wire  _GEN_3165 = unuse_way == 2'h2 ? _GEN_1244 : _GEN_2781; // @[i_cache.scala 91:40]
  wire  _GEN_3166 = unuse_way == 2'h2 ? _GEN_1245 : _GEN_2782; // @[i_cache.scala 91:40]
  wire  _GEN_3167 = unuse_way == 2'h2 ? _GEN_1246 : _GEN_2783; // @[i_cache.scala 91:40]
  wire  _GEN_3168 = unuse_way == 2'h2 ? _GEN_1247 : _GEN_2784; // @[i_cache.scala 91:40]
  wire  _GEN_3169 = unuse_way == 2'h2 ? _GEN_1248 : _GEN_2785; // @[i_cache.scala 91:40]
  wire  _GEN_3170 = unuse_way == 2'h2 ? _GEN_1249 : _GEN_2786; // @[i_cache.scala 91:40]
  wire  _GEN_3171 = unuse_way == 2'h2 ? _GEN_1250 : _GEN_2787; // @[i_cache.scala 91:40]
  wire  _GEN_3172 = unuse_way == 2'h2 ? _GEN_1251 : _GEN_2788; // @[i_cache.scala 91:40]
  wire  _GEN_3173 = unuse_way == 2'h2 ? _GEN_1252 : _GEN_2789; // @[i_cache.scala 91:40]
  wire  _GEN_3174 = unuse_way == 2'h2 ? _GEN_1253 : _GEN_2790; // @[i_cache.scala 91:40]
  wire  _GEN_3175 = unuse_way == 2'h2 ? _GEN_1254 : _GEN_2791; // @[i_cache.scala 91:40]
  wire  _GEN_3176 = unuse_way == 2'h2 ? _GEN_1255 : _GEN_2792; // @[i_cache.scala 91:40]
  wire  _GEN_3177 = unuse_way == 2'h2 ? _GEN_1256 : _GEN_2793; // @[i_cache.scala 91:40]
  wire  _GEN_3178 = unuse_way == 2'h2 ? _GEN_1257 : _GEN_2794; // @[i_cache.scala 91:40]
  wire  _GEN_3179 = unuse_way == 2'h2 ? _GEN_1258 : _GEN_2795; // @[i_cache.scala 91:40]
  wire  _GEN_3180 = unuse_way == 2'h2 ? _GEN_1259 : _GEN_2796; // @[i_cache.scala 91:40]
  wire  _GEN_3181 = unuse_way == 2'h2 ? _GEN_1260 : _GEN_2797; // @[i_cache.scala 91:40]
  wire  _GEN_3182 = unuse_way == 2'h2 ? _GEN_1261 : _GEN_2798; // @[i_cache.scala 91:40]
  wire  _GEN_3183 = unuse_way == 2'h2 ? _GEN_1262 : _GEN_2799; // @[i_cache.scala 91:40]
  wire  _GEN_3184 = unuse_way == 2'h2 ? _GEN_1263 : _GEN_2800; // @[i_cache.scala 91:40]
  wire  _GEN_3185 = unuse_way == 2'h2 ? _GEN_1264 : _GEN_2801; // @[i_cache.scala 91:40]
  wire  _GEN_3186 = unuse_way == 2'h2 ? _GEN_1265 : _GEN_2802; // @[i_cache.scala 91:40]
  wire  _GEN_3187 = unuse_way == 2'h2 ? _GEN_1266 : _GEN_2803; // @[i_cache.scala 91:40]
  wire  _GEN_3188 = unuse_way == 2'h2 ? _GEN_1267 : _GEN_2804; // @[i_cache.scala 91:40]
  wire  _GEN_3189 = unuse_way == 2'h2 ? _GEN_1268 : _GEN_2805; // @[i_cache.scala 91:40]
  wire  _GEN_3190 = unuse_way == 2'h2 ? _GEN_1269 : _GEN_2806; // @[i_cache.scala 91:40]
  wire  _GEN_3191 = unuse_way == 2'h2 ? _GEN_1270 : _GEN_2807; // @[i_cache.scala 91:40]
  wire  _GEN_3192 = unuse_way == 2'h2 ? _GEN_1271 : _GEN_2808; // @[i_cache.scala 91:40]
  wire  _GEN_3193 = unuse_way == 2'h2 ? _GEN_1272 : _GEN_2809; // @[i_cache.scala 91:40]
  wire  _GEN_3194 = unuse_way == 2'h2 ? _GEN_1273 : _GEN_2810; // @[i_cache.scala 91:40]
  wire  _GEN_3195 = unuse_way == 2'h2 ? _GEN_1274 : _GEN_2811; // @[i_cache.scala 91:40]
  wire  _GEN_3196 = unuse_way == 2'h2 ? _GEN_1275 : _GEN_2812; // @[i_cache.scala 91:40]
  wire  _GEN_3197 = unuse_way == 2'h2 ? _GEN_1276 : _GEN_2813; // @[i_cache.scala 91:40]
  wire  _GEN_3198 = unuse_way == 2'h2 ? _GEN_1277 : _GEN_2814; // @[i_cache.scala 91:40]
  wire  _GEN_3199 = unuse_way == 2'h2 ? _GEN_1278 : _GEN_2815; // @[i_cache.scala 91:40]
  wire  _GEN_3200 = unuse_way == 2'h2 ? _GEN_1279 : _GEN_2816; // @[i_cache.scala 91:40]
  wire  _GEN_3201 = unuse_way == 2'h2 ? _GEN_1280 : _GEN_2817; // @[i_cache.scala 91:40]
  wire  _GEN_3202 = unuse_way == 2'h2 ? _GEN_1281 : _GEN_2818; // @[i_cache.scala 91:40]
  wire  _GEN_3203 = unuse_way == 2'h2 ? _GEN_1282 : _GEN_2819; // @[i_cache.scala 91:40]
  wire  _GEN_3204 = unuse_way == 2'h2 ? _GEN_1283 : _GEN_2820; // @[i_cache.scala 91:40]
  wire  _GEN_3205 = unuse_way == 2'h2 ? _GEN_1284 : _GEN_2821; // @[i_cache.scala 91:40]
  wire  _GEN_3206 = unuse_way == 2'h2 ? _GEN_1285 : _GEN_2822; // @[i_cache.scala 91:40]
  wire  _GEN_3207 = unuse_way == 2'h2 ? _GEN_1286 : _GEN_2823; // @[i_cache.scala 91:40]
  wire  _GEN_3208 = unuse_way == 2'h2 ? _GEN_1287 : _GEN_2824; // @[i_cache.scala 91:40]
  wire  _GEN_3209 = unuse_way == 2'h2 ? _GEN_1288 : _GEN_2825; // @[i_cache.scala 91:40]
  wire  _GEN_3210 = unuse_way == 2'h2 ? _GEN_1289 : _GEN_2826; // @[i_cache.scala 91:40]
  wire  _GEN_3211 = unuse_way == 2'h2 ? 1'h0 : _T_14; // @[i_cache.scala 91:40 95:23]
  wire [63:0] _GEN_3212 = unuse_way == 2'h2 ? ram_0_0 : _GEN_2058; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3213 = unuse_way == 2'h2 ? ram_0_1 : _GEN_2059; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3214 = unuse_way == 2'h2 ? ram_0_2 : _GEN_2060; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3215 = unuse_way == 2'h2 ? ram_0_3 : _GEN_2061; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3216 = unuse_way == 2'h2 ? ram_0_4 : _GEN_2062; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3217 = unuse_way == 2'h2 ? ram_0_5 : _GEN_2063; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3218 = unuse_way == 2'h2 ? ram_0_6 : _GEN_2064; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3219 = unuse_way == 2'h2 ? ram_0_7 : _GEN_2065; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3220 = unuse_way == 2'h2 ? ram_0_8 : _GEN_2066; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3221 = unuse_way == 2'h2 ? ram_0_9 : _GEN_2067; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3222 = unuse_way == 2'h2 ? ram_0_10 : _GEN_2068; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3223 = unuse_way == 2'h2 ? ram_0_11 : _GEN_2069; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3224 = unuse_way == 2'h2 ? ram_0_12 : _GEN_2070; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3225 = unuse_way == 2'h2 ? ram_0_13 : _GEN_2071; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3226 = unuse_way == 2'h2 ? ram_0_14 : _GEN_2072; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3227 = unuse_way == 2'h2 ? ram_0_15 : _GEN_2073; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3228 = unuse_way == 2'h2 ? ram_0_16 : _GEN_2074; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3229 = unuse_way == 2'h2 ? ram_0_17 : _GEN_2075; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3230 = unuse_way == 2'h2 ? ram_0_18 : _GEN_2076; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3231 = unuse_way == 2'h2 ? ram_0_19 : _GEN_2077; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3232 = unuse_way == 2'h2 ? ram_0_20 : _GEN_2078; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3233 = unuse_way == 2'h2 ? ram_0_21 : _GEN_2079; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3234 = unuse_way == 2'h2 ? ram_0_22 : _GEN_2080; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3235 = unuse_way == 2'h2 ? ram_0_23 : _GEN_2081; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3236 = unuse_way == 2'h2 ? ram_0_24 : _GEN_2082; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3237 = unuse_way == 2'h2 ? ram_0_25 : _GEN_2083; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3238 = unuse_way == 2'h2 ? ram_0_26 : _GEN_2084; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3239 = unuse_way == 2'h2 ? ram_0_27 : _GEN_2085; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3240 = unuse_way == 2'h2 ? ram_0_28 : _GEN_2086; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3241 = unuse_way == 2'h2 ? ram_0_29 : _GEN_2087; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3242 = unuse_way == 2'h2 ? ram_0_30 : _GEN_2088; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3243 = unuse_way == 2'h2 ? ram_0_31 : _GEN_2089; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3244 = unuse_way == 2'h2 ? ram_0_32 : _GEN_2090; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3245 = unuse_way == 2'h2 ? ram_0_33 : _GEN_2091; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3246 = unuse_way == 2'h2 ? ram_0_34 : _GEN_2092; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3247 = unuse_way == 2'h2 ? ram_0_35 : _GEN_2093; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3248 = unuse_way == 2'h2 ? ram_0_36 : _GEN_2094; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3249 = unuse_way == 2'h2 ? ram_0_37 : _GEN_2095; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3250 = unuse_way == 2'h2 ? ram_0_38 : _GEN_2096; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3251 = unuse_way == 2'h2 ? ram_0_39 : _GEN_2097; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3252 = unuse_way == 2'h2 ? ram_0_40 : _GEN_2098; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3253 = unuse_way == 2'h2 ? ram_0_41 : _GEN_2099; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3254 = unuse_way == 2'h2 ? ram_0_42 : _GEN_2100; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3255 = unuse_way == 2'h2 ? ram_0_43 : _GEN_2101; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3256 = unuse_way == 2'h2 ? ram_0_44 : _GEN_2102; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3257 = unuse_way == 2'h2 ? ram_0_45 : _GEN_2103; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3258 = unuse_way == 2'h2 ? ram_0_46 : _GEN_2104; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3259 = unuse_way == 2'h2 ? ram_0_47 : _GEN_2105; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3260 = unuse_way == 2'h2 ? ram_0_48 : _GEN_2106; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3261 = unuse_way == 2'h2 ? ram_0_49 : _GEN_2107; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3262 = unuse_way == 2'h2 ? ram_0_50 : _GEN_2108; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3263 = unuse_way == 2'h2 ? ram_0_51 : _GEN_2109; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3264 = unuse_way == 2'h2 ? ram_0_52 : _GEN_2110; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3265 = unuse_way == 2'h2 ? ram_0_53 : _GEN_2111; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3266 = unuse_way == 2'h2 ? ram_0_54 : _GEN_2112; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3267 = unuse_way == 2'h2 ? ram_0_55 : _GEN_2113; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3268 = unuse_way == 2'h2 ? ram_0_56 : _GEN_2114; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3269 = unuse_way == 2'h2 ? ram_0_57 : _GEN_2115; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3270 = unuse_way == 2'h2 ? ram_0_58 : _GEN_2116; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3271 = unuse_way == 2'h2 ? ram_0_59 : _GEN_2117; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3272 = unuse_way == 2'h2 ? ram_0_60 : _GEN_2118; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3273 = unuse_way == 2'h2 ? ram_0_61 : _GEN_2119; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3274 = unuse_way == 2'h2 ? ram_0_62 : _GEN_2120; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3275 = unuse_way == 2'h2 ? ram_0_63 : _GEN_2121; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3276 = unuse_way == 2'h2 ? ram_0_64 : _GEN_2122; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3277 = unuse_way == 2'h2 ? ram_0_65 : _GEN_2123; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3278 = unuse_way == 2'h2 ? ram_0_66 : _GEN_2124; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3279 = unuse_way == 2'h2 ? ram_0_67 : _GEN_2125; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3280 = unuse_way == 2'h2 ? ram_0_68 : _GEN_2126; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3281 = unuse_way == 2'h2 ? ram_0_69 : _GEN_2127; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3282 = unuse_way == 2'h2 ? ram_0_70 : _GEN_2128; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3283 = unuse_way == 2'h2 ? ram_0_71 : _GEN_2129; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3284 = unuse_way == 2'h2 ? ram_0_72 : _GEN_2130; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3285 = unuse_way == 2'h2 ? ram_0_73 : _GEN_2131; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3286 = unuse_way == 2'h2 ? ram_0_74 : _GEN_2132; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3287 = unuse_way == 2'h2 ? ram_0_75 : _GEN_2133; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3288 = unuse_way == 2'h2 ? ram_0_76 : _GEN_2134; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3289 = unuse_way == 2'h2 ? ram_0_77 : _GEN_2135; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3290 = unuse_way == 2'h2 ? ram_0_78 : _GEN_2136; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3291 = unuse_way == 2'h2 ? ram_0_79 : _GEN_2137; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3292 = unuse_way == 2'h2 ? ram_0_80 : _GEN_2138; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3293 = unuse_way == 2'h2 ? ram_0_81 : _GEN_2139; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3294 = unuse_way == 2'h2 ? ram_0_82 : _GEN_2140; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3295 = unuse_way == 2'h2 ? ram_0_83 : _GEN_2141; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3296 = unuse_way == 2'h2 ? ram_0_84 : _GEN_2142; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3297 = unuse_way == 2'h2 ? ram_0_85 : _GEN_2143; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3298 = unuse_way == 2'h2 ? ram_0_86 : _GEN_2144; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3299 = unuse_way == 2'h2 ? ram_0_87 : _GEN_2145; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3300 = unuse_way == 2'h2 ? ram_0_88 : _GEN_2146; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3301 = unuse_way == 2'h2 ? ram_0_89 : _GEN_2147; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3302 = unuse_way == 2'h2 ? ram_0_90 : _GEN_2148; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3303 = unuse_way == 2'h2 ? ram_0_91 : _GEN_2149; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3304 = unuse_way == 2'h2 ? ram_0_92 : _GEN_2150; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3305 = unuse_way == 2'h2 ? ram_0_93 : _GEN_2151; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3306 = unuse_way == 2'h2 ? ram_0_94 : _GEN_2152; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3307 = unuse_way == 2'h2 ? ram_0_95 : _GEN_2153; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3308 = unuse_way == 2'h2 ? ram_0_96 : _GEN_2154; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3309 = unuse_way == 2'h2 ? ram_0_97 : _GEN_2155; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3310 = unuse_way == 2'h2 ? ram_0_98 : _GEN_2156; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3311 = unuse_way == 2'h2 ? ram_0_99 : _GEN_2157; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3312 = unuse_way == 2'h2 ? ram_0_100 : _GEN_2158; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3313 = unuse_way == 2'h2 ? ram_0_101 : _GEN_2159; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3314 = unuse_way == 2'h2 ? ram_0_102 : _GEN_2160; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3315 = unuse_way == 2'h2 ? ram_0_103 : _GEN_2161; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3316 = unuse_way == 2'h2 ? ram_0_104 : _GEN_2162; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3317 = unuse_way == 2'h2 ? ram_0_105 : _GEN_2163; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3318 = unuse_way == 2'h2 ? ram_0_106 : _GEN_2164; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3319 = unuse_way == 2'h2 ? ram_0_107 : _GEN_2165; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3320 = unuse_way == 2'h2 ? ram_0_108 : _GEN_2166; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3321 = unuse_way == 2'h2 ? ram_0_109 : _GEN_2167; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3322 = unuse_way == 2'h2 ? ram_0_110 : _GEN_2168; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3323 = unuse_way == 2'h2 ? ram_0_111 : _GEN_2169; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3324 = unuse_way == 2'h2 ? ram_0_112 : _GEN_2170; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3325 = unuse_way == 2'h2 ? ram_0_113 : _GEN_2171; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3326 = unuse_way == 2'h2 ? ram_0_114 : _GEN_2172; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3327 = unuse_way == 2'h2 ? ram_0_115 : _GEN_2173; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3328 = unuse_way == 2'h2 ? ram_0_116 : _GEN_2174; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3329 = unuse_way == 2'h2 ? ram_0_117 : _GEN_2175; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3330 = unuse_way == 2'h2 ? ram_0_118 : _GEN_2176; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3331 = unuse_way == 2'h2 ? ram_0_119 : _GEN_2177; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3332 = unuse_way == 2'h2 ? ram_0_120 : _GEN_2178; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3333 = unuse_way == 2'h2 ? ram_0_121 : _GEN_2179; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3334 = unuse_way == 2'h2 ? ram_0_122 : _GEN_2180; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3335 = unuse_way == 2'h2 ? ram_0_123 : _GEN_2181; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3336 = unuse_way == 2'h2 ? ram_0_124 : _GEN_2182; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3337 = unuse_way == 2'h2 ? ram_0_125 : _GEN_2183; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3338 = unuse_way == 2'h2 ? ram_0_126 : _GEN_2184; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3339 = unuse_way == 2'h2 ? ram_0_127 : _GEN_2185; // @[i_cache.scala 17:24 91:40]
  wire [31:0] _GEN_3340 = unuse_way == 2'h2 ? tag_0_0 : _GEN_2186; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3341 = unuse_way == 2'h2 ? tag_0_1 : _GEN_2187; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3342 = unuse_way == 2'h2 ? tag_0_2 : _GEN_2188; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3343 = unuse_way == 2'h2 ? tag_0_3 : _GEN_2189; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3344 = unuse_way == 2'h2 ? tag_0_4 : _GEN_2190; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3345 = unuse_way == 2'h2 ? tag_0_5 : _GEN_2191; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3346 = unuse_way == 2'h2 ? tag_0_6 : _GEN_2192; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3347 = unuse_way == 2'h2 ? tag_0_7 : _GEN_2193; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3348 = unuse_way == 2'h2 ? tag_0_8 : _GEN_2194; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3349 = unuse_way == 2'h2 ? tag_0_9 : _GEN_2195; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3350 = unuse_way == 2'h2 ? tag_0_10 : _GEN_2196; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3351 = unuse_way == 2'h2 ? tag_0_11 : _GEN_2197; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3352 = unuse_way == 2'h2 ? tag_0_12 : _GEN_2198; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3353 = unuse_way == 2'h2 ? tag_0_13 : _GEN_2199; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3354 = unuse_way == 2'h2 ? tag_0_14 : _GEN_2200; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3355 = unuse_way == 2'h2 ? tag_0_15 : _GEN_2201; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3356 = unuse_way == 2'h2 ? tag_0_16 : _GEN_2202; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3357 = unuse_way == 2'h2 ? tag_0_17 : _GEN_2203; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3358 = unuse_way == 2'h2 ? tag_0_18 : _GEN_2204; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3359 = unuse_way == 2'h2 ? tag_0_19 : _GEN_2205; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3360 = unuse_way == 2'h2 ? tag_0_20 : _GEN_2206; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3361 = unuse_way == 2'h2 ? tag_0_21 : _GEN_2207; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3362 = unuse_way == 2'h2 ? tag_0_22 : _GEN_2208; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3363 = unuse_way == 2'h2 ? tag_0_23 : _GEN_2209; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3364 = unuse_way == 2'h2 ? tag_0_24 : _GEN_2210; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3365 = unuse_way == 2'h2 ? tag_0_25 : _GEN_2211; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3366 = unuse_way == 2'h2 ? tag_0_26 : _GEN_2212; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3367 = unuse_way == 2'h2 ? tag_0_27 : _GEN_2213; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3368 = unuse_way == 2'h2 ? tag_0_28 : _GEN_2214; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3369 = unuse_way == 2'h2 ? tag_0_29 : _GEN_2215; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3370 = unuse_way == 2'h2 ? tag_0_30 : _GEN_2216; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3371 = unuse_way == 2'h2 ? tag_0_31 : _GEN_2217; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3372 = unuse_way == 2'h2 ? tag_0_32 : _GEN_2218; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3373 = unuse_way == 2'h2 ? tag_0_33 : _GEN_2219; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3374 = unuse_way == 2'h2 ? tag_0_34 : _GEN_2220; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3375 = unuse_way == 2'h2 ? tag_0_35 : _GEN_2221; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3376 = unuse_way == 2'h2 ? tag_0_36 : _GEN_2222; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3377 = unuse_way == 2'h2 ? tag_0_37 : _GEN_2223; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3378 = unuse_way == 2'h2 ? tag_0_38 : _GEN_2224; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3379 = unuse_way == 2'h2 ? tag_0_39 : _GEN_2225; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3380 = unuse_way == 2'h2 ? tag_0_40 : _GEN_2226; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3381 = unuse_way == 2'h2 ? tag_0_41 : _GEN_2227; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3382 = unuse_way == 2'h2 ? tag_0_42 : _GEN_2228; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3383 = unuse_way == 2'h2 ? tag_0_43 : _GEN_2229; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3384 = unuse_way == 2'h2 ? tag_0_44 : _GEN_2230; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3385 = unuse_way == 2'h2 ? tag_0_45 : _GEN_2231; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3386 = unuse_way == 2'h2 ? tag_0_46 : _GEN_2232; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3387 = unuse_way == 2'h2 ? tag_0_47 : _GEN_2233; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3388 = unuse_way == 2'h2 ? tag_0_48 : _GEN_2234; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3389 = unuse_way == 2'h2 ? tag_0_49 : _GEN_2235; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3390 = unuse_way == 2'h2 ? tag_0_50 : _GEN_2236; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3391 = unuse_way == 2'h2 ? tag_0_51 : _GEN_2237; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3392 = unuse_way == 2'h2 ? tag_0_52 : _GEN_2238; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3393 = unuse_way == 2'h2 ? tag_0_53 : _GEN_2239; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3394 = unuse_way == 2'h2 ? tag_0_54 : _GEN_2240; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3395 = unuse_way == 2'h2 ? tag_0_55 : _GEN_2241; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3396 = unuse_way == 2'h2 ? tag_0_56 : _GEN_2242; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3397 = unuse_way == 2'h2 ? tag_0_57 : _GEN_2243; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3398 = unuse_way == 2'h2 ? tag_0_58 : _GEN_2244; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3399 = unuse_way == 2'h2 ? tag_0_59 : _GEN_2245; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3400 = unuse_way == 2'h2 ? tag_0_60 : _GEN_2246; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3401 = unuse_way == 2'h2 ? tag_0_61 : _GEN_2247; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3402 = unuse_way == 2'h2 ? tag_0_62 : _GEN_2248; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3403 = unuse_way == 2'h2 ? tag_0_63 : _GEN_2249; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3404 = unuse_way == 2'h2 ? tag_0_64 : _GEN_2250; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3405 = unuse_way == 2'h2 ? tag_0_65 : _GEN_2251; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3406 = unuse_way == 2'h2 ? tag_0_66 : _GEN_2252; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3407 = unuse_way == 2'h2 ? tag_0_67 : _GEN_2253; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3408 = unuse_way == 2'h2 ? tag_0_68 : _GEN_2254; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3409 = unuse_way == 2'h2 ? tag_0_69 : _GEN_2255; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3410 = unuse_way == 2'h2 ? tag_0_70 : _GEN_2256; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3411 = unuse_way == 2'h2 ? tag_0_71 : _GEN_2257; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3412 = unuse_way == 2'h2 ? tag_0_72 : _GEN_2258; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3413 = unuse_way == 2'h2 ? tag_0_73 : _GEN_2259; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3414 = unuse_way == 2'h2 ? tag_0_74 : _GEN_2260; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3415 = unuse_way == 2'h2 ? tag_0_75 : _GEN_2261; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3416 = unuse_way == 2'h2 ? tag_0_76 : _GEN_2262; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3417 = unuse_way == 2'h2 ? tag_0_77 : _GEN_2263; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3418 = unuse_way == 2'h2 ? tag_0_78 : _GEN_2264; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3419 = unuse_way == 2'h2 ? tag_0_79 : _GEN_2265; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3420 = unuse_way == 2'h2 ? tag_0_80 : _GEN_2266; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3421 = unuse_way == 2'h2 ? tag_0_81 : _GEN_2267; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3422 = unuse_way == 2'h2 ? tag_0_82 : _GEN_2268; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3423 = unuse_way == 2'h2 ? tag_0_83 : _GEN_2269; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3424 = unuse_way == 2'h2 ? tag_0_84 : _GEN_2270; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3425 = unuse_way == 2'h2 ? tag_0_85 : _GEN_2271; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3426 = unuse_way == 2'h2 ? tag_0_86 : _GEN_2272; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3427 = unuse_way == 2'h2 ? tag_0_87 : _GEN_2273; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3428 = unuse_way == 2'h2 ? tag_0_88 : _GEN_2274; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3429 = unuse_way == 2'h2 ? tag_0_89 : _GEN_2275; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3430 = unuse_way == 2'h2 ? tag_0_90 : _GEN_2276; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3431 = unuse_way == 2'h2 ? tag_0_91 : _GEN_2277; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3432 = unuse_way == 2'h2 ? tag_0_92 : _GEN_2278; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3433 = unuse_way == 2'h2 ? tag_0_93 : _GEN_2279; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3434 = unuse_way == 2'h2 ? tag_0_94 : _GEN_2280; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3435 = unuse_way == 2'h2 ? tag_0_95 : _GEN_2281; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3436 = unuse_way == 2'h2 ? tag_0_96 : _GEN_2282; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3437 = unuse_way == 2'h2 ? tag_0_97 : _GEN_2283; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3438 = unuse_way == 2'h2 ? tag_0_98 : _GEN_2284; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3439 = unuse_way == 2'h2 ? tag_0_99 : _GEN_2285; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3440 = unuse_way == 2'h2 ? tag_0_100 : _GEN_2286; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3441 = unuse_way == 2'h2 ? tag_0_101 : _GEN_2287; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3442 = unuse_way == 2'h2 ? tag_0_102 : _GEN_2288; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3443 = unuse_way == 2'h2 ? tag_0_103 : _GEN_2289; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3444 = unuse_way == 2'h2 ? tag_0_104 : _GEN_2290; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3445 = unuse_way == 2'h2 ? tag_0_105 : _GEN_2291; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3446 = unuse_way == 2'h2 ? tag_0_106 : _GEN_2292; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3447 = unuse_way == 2'h2 ? tag_0_107 : _GEN_2293; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3448 = unuse_way == 2'h2 ? tag_0_108 : _GEN_2294; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3449 = unuse_way == 2'h2 ? tag_0_109 : _GEN_2295; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3450 = unuse_way == 2'h2 ? tag_0_110 : _GEN_2296; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3451 = unuse_way == 2'h2 ? tag_0_111 : _GEN_2297; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3452 = unuse_way == 2'h2 ? tag_0_112 : _GEN_2298; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3453 = unuse_way == 2'h2 ? tag_0_113 : _GEN_2299; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3454 = unuse_way == 2'h2 ? tag_0_114 : _GEN_2300; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3455 = unuse_way == 2'h2 ? tag_0_115 : _GEN_2301; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3456 = unuse_way == 2'h2 ? tag_0_116 : _GEN_2302; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3457 = unuse_way == 2'h2 ? tag_0_117 : _GEN_2303; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3458 = unuse_way == 2'h2 ? tag_0_118 : _GEN_2304; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3459 = unuse_way == 2'h2 ? tag_0_119 : _GEN_2305; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3460 = unuse_way == 2'h2 ? tag_0_120 : _GEN_2306; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3461 = unuse_way == 2'h2 ? tag_0_121 : _GEN_2307; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3462 = unuse_way == 2'h2 ? tag_0_122 : _GEN_2308; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3463 = unuse_way == 2'h2 ? tag_0_123 : _GEN_2309; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3464 = unuse_way == 2'h2 ? tag_0_124 : _GEN_2310; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3465 = unuse_way == 2'h2 ? tag_0_125 : _GEN_2311; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3466 = unuse_way == 2'h2 ? tag_0_126 : _GEN_2312; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3467 = unuse_way == 2'h2 ? tag_0_127 : _GEN_2313; // @[i_cache.scala 19:24 91:40]
  wire  _GEN_3468 = unuse_way == 2'h2 ? valid_0_0 : _GEN_2314; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3469 = unuse_way == 2'h2 ? valid_0_1 : _GEN_2315; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3470 = unuse_way == 2'h2 ? valid_0_2 : _GEN_2316; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3471 = unuse_way == 2'h2 ? valid_0_3 : _GEN_2317; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3472 = unuse_way == 2'h2 ? valid_0_4 : _GEN_2318; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3473 = unuse_way == 2'h2 ? valid_0_5 : _GEN_2319; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3474 = unuse_way == 2'h2 ? valid_0_6 : _GEN_2320; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3475 = unuse_way == 2'h2 ? valid_0_7 : _GEN_2321; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3476 = unuse_way == 2'h2 ? valid_0_8 : _GEN_2322; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3477 = unuse_way == 2'h2 ? valid_0_9 : _GEN_2323; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3478 = unuse_way == 2'h2 ? valid_0_10 : _GEN_2324; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3479 = unuse_way == 2'h2 ? valid_0_11 : _GEN_2325; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3480 = unuse_way == 2'h2 ? valid_0_12 : _GEN_2326; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3481 = unuse_way == 2'h2 ? valid_0_13 : _GEN_2327; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3482 = unuse_way == 2'h2 ? valid_0_14 : _GEN_2328; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3483 = unuse_way == 2'h2 ? valid_0_15 : _GEN_2329; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3484 = unuse_way == 2'h2 ? valid_0_16 : _GEN_2330; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3485 = unuse_way == 2'h2 ? valid_0_17 : _GEN_2331; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3486 = unuse_way == 2'h2 ? valid_0_18 : _GEN_2332; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3487 = unuse_way == 2'h2 ? valid_0_19 : _GEN_2333; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3488 = unuse_way == 2'h2 ? valid_0_20 : _GEN_2334; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3489 = unuse_way == 2'h2 ? valid_0_21 : _GEN_2335; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3490 = unuse_way == 2'h2 ? valid_0_22 : _GEN_2336; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3491 = unuse_way == 2'h2 ? valid_0_23 : _GEN_2337; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3492 = unuse_way == 2'h2 ? valid_0_24 : _GEN_2338; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3493 = unuse_way == 2'h2 ? valid_0_25 : _GEN_2339; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3494 = unuse_way == 2'h2 ? valid_0_26 : _GEN_2340; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3495 = unuse_way == 2'h2 ? valid_0_27 : _GEN_2341; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3496 = unuse_way == 2'h2 ? valid_0_28 : _GEN_2342; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3497 = unuse_way == 2'h2 ? valid_0_29 : _GEN_2343; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3498 = unuse_way == 2'h2 ? valid_0_30 : _GEN_2344; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3499 = unuse_way == 2'h2 ? valid_0_31 : _GEN_2345; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3500 = unuse_way == 2'h2 ? valid_0_32 : _GEN_2346; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3501 = unuse_way == 2'h2 ? valid_0_33 : _GEN_2347; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3502 = unuse_way == 2'h2 ? valid_0_34 : _GEN_2348; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3503 = unuse_way == 2'h2 ? valid_0_35 : _GEN_2349; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3504 = unuse_way == 2'h2 ? valid_0_36 : _GEN_2350; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3505 = unuse_way == 2'h2 ? valid_0_37 : _GEN_2351; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3506 = unuse_way == 2'h2 ? valid_0_38 : _GEN_2352; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3507 = unuse_way == 2'h2 ? valid_0_39 : _GEN_2353; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3508 = unuse_way == 2'h2 ? valid_0_40 : _GEN_2354; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3509 = unuse_way == 2'h2 ? valid_0_41 : _GEN_2355; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3510 = unuse_way == 2'h2 ? valid_0_42 : _GEN_2356; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3511 = unuse_way == 2'h2 ? valid_0_43 : _GEN_2357; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3512 = unuse_way == 2'h2 ? valid_0_44 : _GEN_2358; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3513 = unuse_way == 2'h2 ? valid_0_45 : _GEN_2359; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3514 = unuse_way == 2'h2 ? valid_0_46 : _GEN_2360; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3515 = unuse_way == 2'h2 ? valid_0_47 : _GEN_2361; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3516 = unuse_way == 2'h2 ? valid_0_48 : _GEN_2362; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3517 = unuse_way == 2'h2 ? valid_0_49 : _GEN_2363; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3518 = unuse_way == 2'h2 ? valid_0_50 : _GEN_2364; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3519 = unuse_way == 2'h2 ? valid_0_51 : _GEN_2365; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3520 = unuse_way == 2'h2 ? valid_0_52 : _GEN_2366; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3521 = unuse_way == 2'h2 ? valid_0_53 : _GEN_2367; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3522 = unuse_way == 2'h2 ? valid_0_54 : _GEN_2368; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3523 = unuse_way == 2'h2 ? valid_0_55 : _GEN_2369; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3524 = unuse_way == 2'h2 ? valid_0_56 : _GEN_2370; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3525 = unuse_way == 2'h2 ? valid_0_57 : _GEN_2371; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3526 = unuse_way == 2'h2 ? valid_0_58 : _GEN_2372; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3527 = unuse_way == 2'h2 ? valid_0_59 : _GEN_2373; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3528 = unuse_way == 2'h2 ? valid_0_60 : _GEN_2374; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3529 = unuse_way == 2'h2 ? valid_0_61 : _GEN_2375; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3530 = unuse_way == 2'h2 ? valid_0_62 : _GEN_2376; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3531 = unuse_way == 2'h2 ? valid_0_63 : _GEN_2377; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3532 = unuse_way == 2'h2 ? valid_0_64 : _GEN_2378; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3533 = unuse_way == 2'h2 ? valid_0_65 : _GEN_2379; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3534 = unuse_way == 2'h2 ? valid_0_66 : _GEN_2380; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3535 = unuse_way == 2'h2 ? valid_0_67 : _GEN_2381; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3536 = unuse_way == 2'h2 ? valid_0_68 : _GEN_2382; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3537 = unuse_way == 2'h2 ? valid_0_69 : _GEN_2383; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3538 = unuse_way == 2'h2 ? valid_0_70 : _GEN_2384; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3539 = unuse_way == 2'h2 ? valid_0_71 : _GEN_2385; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3540 = unuse_way == 2'h2 ? valid_0_72 : _GEN_2386; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3541 = unuse_way == 2'h2 ? valid_0_73 : _GEN_2387; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3542 = unuse_way == 2'h2 ? valid_0_74 : _GEN_2388; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3543 = unuse_way == 2'h2 ? valid_0_75 : _GEN_2389; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3544 = unuse_way == 2'h2 ? valid_0_76 : _GEN_2390; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3545 = unuse_way == 2'h2 ? valid_0_77 : _GEN_2391; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3546 = unuse_way == 2'h2 ? valid_0_78 : _GEN_2392; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3547 = unuse_way == 2'h2 ? valid_0_79 : _GEN_2393; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3548 = unuse_way == 2'h2 ? valid_0_80 : _GEN_2394; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3549 = unuse_way == 2'h2 ? valid_0_81 : _GEN_2395; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3550 = unuse_way == 2'h2 ? valid_0_82 : _GEN_2396; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3551 = unuse_way == 2'h2 ? valid_0_83 : _GEN_2397; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3552 = unuse_way == 2'h2 ? valid_0_84 : _GEN_2398; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3553 = unuse_way == 2'h2 ? valid_0_85 : _GEN_2399; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3554 = unuse_way == 2'h2 ? valid_0_86 : _GEN_2400; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3555 = unuse_way == 2'h2 ? valid_0_87 : _GEN_2401; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3556 = unuse_way == 2'h2 ? valid_0_88 : _GEN_2402; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3557 = unuse_way == 2'h2 ? valid_0_89 : _GEN_2403; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3558 = unuse_way == 2'h2 ? valid_0_90 : _GEN_2404; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3559 = unuse_way == 2'h2 ? valid_0_91 : _GEN_2405; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3560 = unuse_way == 2'h2 ? valid_0_92 : _GEN_2406; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3561 = unuse_way == 2'h2 ? valid_0_93 : _GEN_2407; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3562 = unuse_way == 2'h2 ? valid_0_94 : _GEN_2408; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3563 = unuse_way == 2'h2 ? valid_0_95 : _GEN_2409; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3564 = unuse_way == 2'h2 ? valid_0_96 : _GEN_2410; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3565 = unuse_way == 2'h2 ? valid_0_97 : _GEN_2411; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3566 = unuse_way == 2'h2 ? valid_0_98 : _GEN_2412; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3567 = unuse_way == 2'h2 ? valid_0_99 : _GEN_2413; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3568 = unuse_way == 2'h2 ? valid_0_100 : _GEN_2414; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3569 = unuse_way == 2'h2 ? valid_0_101 : _GEN_2415; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3570 = unuse_way == 2'h2 ? valid_0_102 : _GEN_2416; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3571 = unuse_way == 2'h2 ? valid_0_103 : _GEN_2417; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3572 = unuse_way == 2'h2 ? valid_0_104 : _GEN_2418; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3573 = unuse_way == 2'h2 ? valid_0_105 : _GEN_2419; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3574 = unuse_way == 2'h2 ? valid_0_106 : _GEN_2420; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3575 = unuse_way == 2'h2 ? valid_0_107 : _GEN_2421; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3576 = unuse_way == 2'h2 ? valid_0_108 : _GEN_2422; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3577 = unuse_way == 2'h2 ? valid_0_109 : _GEN_2423; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3578 = unuse_way == 2'h2 ? valid_0_110 : _GEN_2424; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3579 = unuse_way == 2'h2 ? valid_0_111 : _GEN_2425; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3580 = unuse_way == 2'h2 ? valid_0_112 : _GEN_2426; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3581 = unuse_way == 2'h2 ? valid_0_113 : _GEN_2427; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3582 = unuse_way == 2'h2 ? valid_0_114 : _GEN_2428; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3583 = unuse_way == 2'h2 ? valid_0_115 : _GEN_2429; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3584 = unuse_way == 2'h2 ? valid_0_116 : _GEN_2430; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3585 = unuse_way == 2'h2 ? valid_0_117 : _GEN_2431; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3586 = unuse_way == 2'h2 ? valid_0_118 : _GEN_2432; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3587 = unuse_way == 2'h2 ? valid_0_119 : _GEN_2433; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3588 = unuse_way == 2'h2 ? valid_0_120 : _GEN_2434; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3589 = unuse_way == 2'h2 ? valid_0_121 : _GEN_2435; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3590 = unuse_way == 2'h2 ? valid_0_122 : _GEN_2436; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3591 = unuse_way == 2'h2 ? valid_0_123 : _GEN_2437; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3592 = unuse_way == 2'h2 ? valid_0_124 : _GEN_2438; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3593 = unuse_way == 2'h2 ? valid_0_125 : _GEN_2439; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3594 = unuse_way == 2'h2 ? valid_0_126 : _GEN_2440; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3595 = unuse_way == 2'h2 ? valid_0_127 : _GEN_2441; // @[i_cache.scala 21:26 91:40]
  wire [63:0] _GEN_3596 = unuse_way == 2'h1 ? _GEN_522 : _GEN_3212; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3597 = unuse_way == 2'h1 ? _GEN_523 : _GEN_3213; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3598 = unuse_way == 2'h1 ? _GEN_524 : _GEN_3214; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3599 = unuse_way == 2'h1 ? _GEN_525 : _GEN_3215; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3600 = unuse_way == 2'h1 ? _GEN_526 : _GEN_3216; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3601 = unuse_way == 2'h1 ? _GEN_527 : _GEN_3217; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3602 = unuse_way == 2'h1 ? _GEN_528 : _GEN_3218; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3603 = unuse_way == 2'h1 ? _GEN_529 : _GEN_3219; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3604 = unuse_way == 2'h1 ? _GEN_530 : _GEN_3220; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3605 = unuse_way == 2'h1 ? _GEN_531 : _GEN_3221; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3606 = unuse_way == 2'h1 ? _GEN_532 : _GEN_3222; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3607 = unuse_way == 2'h1 ? _GEN_533 : _GEN_3223; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3608 = unuse_way == 2'h1 ? _GEN_534 : _GEN_3224; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3609 = unuse_way == 2'h1 ? _GEN_535 : _GEN_3225; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3610 = unuse_way == 2'h1 ? _GEN_536 : _GEN_3226; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3611 = unuse_way == 2'h1 ? _GEN_537 : _GEN_3227; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3612 = unuse_way == 2'h1 ? _GEN_538 : _GEN_3228; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3613 = unuse_way == 2'h1 ? _GEN_539 : _GEN_3229; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3614 = unuse_way == 2'h1 ? _GEN_540 : _GEN_3230; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3615 = unuse_way == 2'h1 ? _GEN_541 : _GEN_3231; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3616 = unuse_way == 2'h1 ? _GEN_542 : _GEN_3232; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3617 = unuse_way == 2'h1 ? _GEN_543 : _GEN_3233; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3618 = unuse_way == 2'h1 ? _GEN_544 : _GEN_3234; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3619 = unuse_way == 2'h1 ? _GEN_545 : _GEN_3235; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3620 = unuse_way == 2'h1 ? _GEN_546 : _GEN_3236; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3621 = unuse_way == 2'h1 ? _GEN_547 : _GEN_3237; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3622 = unuse_way == 2'h1 ? _GEN_548 : _GEN_3238; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3623 = unuse_way == 2'h1 ? _GEN_549 : _GEN_3239; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3624 = unuse_way == 2'h1 ? _GEN_550 : _GEN_3240; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3625 = unuse_way == 2'h1 ? _GEN_551 : _GEN_3241; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3626 = unuse_way == 2'h1 ? _GEN_552 : _GEN_3242; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3627 = unuse_way == 2'h1 ? _GEN_553 : _GEN_3243; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3628 = unuse_way == 2'h1 ? _GEN_554 : _GEN_3244; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3629 = unuse_way == 2'h1 ? _GEN_555 : _GEN_3245; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3630 = unuse_way == 2'h1 ? _GEN_556 : _GEN_3246; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3631 = unuse_way == 2'h1 ? _GEN_557 : _GEN_3247; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3632 = unuse_way == 2'h1 ? _GEN_558 : _GEN_3248; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3633 = unuse_way == 2'h1 ? _GEN_559 : _GEN_3249; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3634 = unuse_way == 2'h1 ? _GEN_560 : _GEN_3250; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3635 = unuse_way == 2'h1 ? _GEN_561 : _GEN_3251; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3636 = unuse_way == 2'h1 ? _GEN_562 : _GEN_3252; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3637 = unuse_way == 2'h1 ? _GEN_563 : _GEN_3253; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3638 = unuse_way == 2'h1 ? _GEN_564 : _GEN_3254; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3639 = unuse_way == 2'h1 ? _GEN_565 : _GEN_3255; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3640 = unuse_way == 2'h1 ? _GEN_566 : _GEN_3256; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3641 = unuse_way == 2'h1 ? _GEN_567 : _GEN_3257; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3642 = unuse_way == 2'h1 ? _GEN_568 : _GEN_3258; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3643 = unuse_way == 2'h1 ? _GEN_569 : _GEN_3259; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3644 = unuse_way == 2'h1 ? _GEN_570 : _GEN_3260; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3645 = unuse_way == 2'h1 ? _GEN_571 : _GEN_3261; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3646 = unuse_way == 2'h1 ? _GEN_572 : _GEN_3262; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3647 = unuse_way == 2'h1 ? _GEN_573 : _GEN_3263; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3648 = unuse_way == 2'h1 ? _GEN_574 : _GEN_3264; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3649 = unuse_way == 2'h1 ? _GEN_575 : _GEN_3265; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3650 = unuse_way == 2'h1 ? _GEN_576 : _GEN_3266; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3651 = unuse_way == 2'h1 ? _GEN_577 : _GEN_3267; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3652 = unuse_way == 2'h1 ? _GEN_578 : _GEN_3268; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3653 = unuse_way == 2'h1 ? _GEN_579 : _GEN_3269; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3654 = unuse_way == 2'h1 ? _GEN_580 : _GEN_3270; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3655 = unuse_way == 2'h1 ? _GEN_581 : _GEN_3271; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3656 = unuse_way == 2'h1 ? _GEN_582 : _GEN_3272; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3657 = unuse_way == 2'h1 ? _GEN_583 : _GEN_3273; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3658 = unuse_way == 2'h1 ? _GEN_584 : _GEN_3274; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3659 = unuse_way == 2'h1 ? _GEN_585 : _GEN_3275; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3660 = unuse_way == 2'h1 ? _GEN_586 : _GEN_3276; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3661 = unuse_way == 2'h1 ? _GEN_587 : _GEN_3277; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3662 = unuse_way == 2'h1 ? _GEN_588 : _GEN_3278; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3663 = unuse_way == 2'h1 ? _GEN_589 : _GEN_3279; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3664 = unuse_way == 2'h1 ? _GEN_590 : _GEN_3280; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3665 = unuse_way == 2'h1 ? _GEN_591 : _GEN_3281; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3666 = unuse_way == 2'h1 ? _GEN_592 : _GEN_3282; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3667 = unuse_way == 2'h1 ? _GEN_593 : _GEN_3283; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3668 = unuse_way == 2'h1 ? _GEN_594 : _GEN_3284; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3669 = unuse_way == 2'h1 ? _GEN_595 : _GEN_3285; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3670 = unuse_way == 2'h1 ? _GEN_596 : _GEN_3286; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3671 = unuse_way == 2'h1 ? _GEN_597 : _GEN_3287; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3672 = unuse_way == 2'h1 ? _GEN_598 : _GEN_3288; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3673 = unuse_way == 2'h1 ? _GEN_599 : _GEN_3289; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3674 = unuse_way == 2'h1 ? _GEN_600 : _GEN_3290; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3675 = unuse_way == 2'h1 ? _GEN_601 : _GEN_3291; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3676 = unuse_way == 2'h1 ? _GEN_602 : _GEN_3292; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3677 = unuse_way == 2'h1 ? _GEN_603 : _GEN_3293; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3678 = unuse_way == 2'h1 ? _GEN_604 : _GEN_3294; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3679 = unuse_way == 2'h1 ? _GEN_605 : _GEN_3295; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3680 = unuse_way == 2'h1 ? _GEN_606 : _GEN_3296; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3681 = unuse_way == 2'h1 ? _GEN_607 : _GEN_3297; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3682 = unuse_way == 2'h1 ? _GEN_608 : _GEN_3298; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3683 = unuse_way == 2'h1 ? _GEN_609 : _GEN_3299; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3684 = unuse_way == 2'h1 ? _GEN_610 : _GEN_3300; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3685 = unuse_way == 2'h1 ? _GEN_611 : _GEN_3301; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3686 = unuse_way == 2'h1 ? _GEN_612 : _GEN_3302; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3687 = unuse_way == 2'h1 ? _GEN_613 : _GEN_3303; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3688 = unuse_way == 2'h1 ? _GEN_614 : _GEN_3304; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3689 = unuse_way == 2'h1 ? _GEN_615 : _GEN_3305; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3690 = unuse_way == 2'h1 ? _GEN_616 : _GEN_3306; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3691 = unuse_way == 2'h1 ? _GEN_617 : _GEN_3307; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3692 = unuse_way == 2'h1 ? _GEN_618 : _GEN_3308; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3693 = unuse_way == 2'h1 ? _GEN_619 : _GEN_3309; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3694 = unuse_way == 2'h1 ? _GEN_620 : _GEN_3310; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3695 = unuse_way == 2'h1 ? _GEN_621 : _GEN_3311; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3696 = unuse_way == 2'h1 ? _GEN_622 : _GEN_3312; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3697 = unuse_way == 2'h1 ? _GEN_623 : _GEN_3313; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3698 = unuse_way == 2'h1 ? _GEN_624 : _GEN_3314; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3699 = unuse_way == 2'h1 ? _GEN_625 : _GEN_3315; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3700 = unuse_way == 2'h1 ? _GEN_626 : _GEN_3316; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3701 = unuse_way == 2'h1 ? _GEN_627 : _GEN_3317; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3702 = unuse_way == 2'h1 ? _GEN_628 : _GEN_3318; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3703 = unuse_way == 2'h1 ? _GEN_629 : _GEN_3319; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3704 = unuse_way == 2'h1 ? _GEN_630 : _GEN_3320; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3705 = unuse_way == 2'h1 ? _GEN_631 : _GEN_3321; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3706 = unuse_way == 2'h1 ? _GEN_632 : _GEN_3322; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3707 = unuse_way == 2'h1 ? _GEN_633 : _GEN_3323; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3708 = unuse_way == 2'h1 ? _GEN_634 : _GEN_3324; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3709 = unuse_way == 2'h1 ? _GEN_635 : _GEN_3325; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3710 = unuse_way == 2'h1 ? _GEN_636 : _GEN_3326; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3711 = unuse_way == 2'h1 ? _GEN_637 : _GEN_3327; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3712 = unuse_way == 2'h1 ? _GEN_638 : _GEN_3328; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3713 = unuse_way == 2'h1 ? _GEN_639 : _GEN_3329; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3714 = unuse_way == 2'h1 ? _GEN_640 : _GEN_3330; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3715 = unuse_way == 2'h1 ? _GEN_641 : _GEN_3331; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3716 = unuse_way == 2'h1 ? _GEN_642 : _GEN_3332; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3717 = unuse_way == 2'h1 ? _GEN_643 : _GEN_3333; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3718 = unuse_way == 2'h1 ? _GEN_644 : _GEN_3334; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3719 = unuse_way == 2'h1 ? _GEN_645 : _GEN_3335; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3720 = unuse_way == 2'h1 ? _GEN_646 : _GEN_3336; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3721 = unuse_way == 2'h1 ? _GEN_647 : _GEN_3337; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3722 = unuse_way == 2'h1 ? _GEN_648 : _GEN_3338; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3723 = unuse_way == 2'h1 ? _GEN_649 : _GEN_3339; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3724 = unuse_way == 2'h1 ? _GEN_650 : _GEN_3340; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3725 = unuse_way == 2'h1 ? _GEN_651 : _GEN_3341; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3726 = unuse_way == 2'h1 ? _GEN_652 : _GEN_3342; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3727 = unuse_way == 2'h1 ? _GEN_653 : _GEN_3343; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3728 = unuse_way == 2'h1 ? _GEN_654 : _GEN_3344; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3729 = unuse_way == 2'h1 ? _GEN_655 : _GEN_3345; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3730 = unuse_way == 2'h1 ? _GEN_656 : _GEN_3346; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3731 = unuse_way == 2'h1 ? _GEN_657 : _GEN_3347; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3732 = unuse_way == 2'h1 ? _GEN_658 : _GEN_3348; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3733 = unuse_way == 2'h1 ? _GEN_659 : _GEN_3349; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3734 = unuse_way == 2'h1 ? _GEN_660 : _GEN_3350; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3735 = unuse_way == 2'h1 ? _GEN_661 : _GEN_3351; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3736 = unuse_way == 2'h1 ? _GEN_662 : _GEN_3352; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3737 = unuse_way == 2'h1 ? _GEN_663 : _GEN_3353; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3738 = unuse_way == 2'h1 ? _GEN_664 : _GEN_3354; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3739 = unuse_way == 2'h1 ? _GEN_665 : _GEN_3355; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3740 = unuse_way == 2'h1 ? _GEN_666 : _GEN_3356; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3741 = unuse_way == 2'h1 ? _GEN_667 : _GEN_3357; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3742 = unuse_way == 2'h1 ? _GEN_668 : _GEN_3358; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3743 = unuse_way == 2'h1 ? _GEN_669 : _GEN_3359; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3744 = unuse_way == 2'h1 ? _GEN_670 : _GEN_3360; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3745 = unuse_way == 2'h1 ? _GEN_671 : _GEN_3361; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3746 = unuse_way == 2'h1 ? _GEN_672 : _GEN_3362; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3747 = unuse_way == 2'h1 ? _GEN_673 : _GEN_3363; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3748 = unuse_way == 2'h1 ? _GEN_674 : _GEN_3364; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3749 = unuse_way == 2'h1 ? _GEN_675 : _GEN_3365; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3750 = unuse_way == 2'h1 ? _GEN_676 : _GEN_3366; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3751 = unuse_way == 2'h1 ? _GEN_677 : _GEN_3367; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3752 = unuse_way == 2'h1 ? _GEN_678 : _GEN_3368; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3753 = unuse_way == 2'h1 ? _GEN_679 : _GEN_3369; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3754 = unuse_way == 2'h1 ? _GEN_680 : _GEN_3370; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3755 = unuse_way == 2'h1 ? _GEN_681 : _GEN_3371; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3756 = unuse_way == 2'h1 ? _GEN_682 : _GEN_3372; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3757 = unuse_way == 2'h1 ? _GEN_683 : _GEN_3373; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3758 = unuse_way == 2'h1 ? _GEN_684 : _GEN_3374; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3759 = unuse_way == 2'h1 ? _GEN_685 : _GEN_3375; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3760 = unuse_way == 2'h1 ? _GEN_686 : _GEN_3376; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3761 = unuse_way == 2'h1 ? _GEN_687 : _GEN_3377; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3762 = unuse_way == 2'h1 ? _GEN_688 : _GEN_3378; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3763 = unuse_way == 2'h1 ? _GEN_689 : _GEN_3379; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3764 = unuse_way == 2'h1 ? _GEN_690 : _GEN_3380; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3765 = unuse_way == 2'h1 ? _GEN_691 : _GEN_3381; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3766 = unuse_way == 2'h1 ? _GEN_692 : _GEN_3382; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3767 = unuse_way == 2'h1 ? _GEN_693 : _GEN_3383; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3768 = unuse_way == 2'h1 ? _GEN_694 : _GEN_3384; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3769 = unuse_way == 2'h1 ? _GEN_695 : _GEN_3385; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3770 = unuse_way == 2'h1 ? _GEN_696 : _GEN_3386; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3771 = unuse_way == 2'h1 ? _GEN_697 : _GEN_3387; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3772 = unuse_way == 2'h1 ? _GEN_698 : _GEN_3388; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3773 = unuse_way == 2'h1 ? _GEN_699 : _GEN_3389; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3774 = unuse_way == 2'h1 ? _GEN_700 : _GEN_3390; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3775 = unuse_way == 2'h1 ? _GEN_701 : _GEN_3391; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3776 = unuse_way == 2'h1 ? _GEN_702 : _GEN_3392; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3777 = unuse_way == 2'h1 ? _GEN_703 : _GEN_3393; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3778 = unuse_way == 2'h1 ? _GEN_704 : _GEN_3394; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3779 = unuse_way == 2'h1 ? _GEN_705 : _GEN_3395; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3780 = unuse_way == 2'h1 ? _GEN_706 : _GEN_3396; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3781 = unuse_way == 2'h1 ? _GEN_707 : _GEN_3397; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3782 = unuse_way == 2'h1 ? _GEN_708 : _GEN_3398; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3783 = unuse_way == 2'h1 ? _GEN_709 : _GEN_3399; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3784 = unuse_way == 2'h1 ? _GEN_710 : _GEN_3400; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3785 = unuse_way == 2'h1 ? _GEN_711 : _GEN_3401; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3786 = unuse_way == 2'h1 ? _GEN_712 : _GEN_3402; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3787 = unuse_way == 2'h1 ? _GEN_713 : _GEN_3403; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3788 = unuse_way == 2'h1 ? _GEN_714 : _GEN_3404; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3789 = unuse_way == 2'h1 ? _GEN_715 : _GEN_3405; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3790 = unuse_way == 2'h1 ? _GEN_716 : _GEN_3406; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3791 = unuse_way == 2'h1 ? _GEN_717 : _GEN_3407; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3792 = unuse_way == 2'h1 ? _GEN_718 : _GEN_3408; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3793 = unuse_way == 2'h1 ? _GEN_719 : _GEN_3409; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3794 = unuse_way == 2'h1 ? _GEN_720 : _GEN_3410; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3795 = unuse_way == 2'h1 ? _GEN_721 : _GEN_3411; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3796 = unuse_way == 2'h1 ? _GEN_722 : _GEN_3412; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3797 = unuse_way == 2'h1 ? _GEN_723 : _GEN_3413; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3798 = unuse_way == 2'h1 ? _GEN_724 : _GEN_3414; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3799 = unuse_way == 2'h1 ? _GEN_725 : _GEN_3415; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3800 = unuse_way == 2'h1 ? _GEN_726 : _GEN_3416; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3801 = unuse_way == 2'h1 ? _GEN_727 : _GEN_3417; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3802 = unuse_way == 2'h1 ? _GEN_728 : _GEN_3418; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3803 = unuse_way == 2'h1 ? _GEN_729 : _GEN_3419; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3804 = unuse_way == 2'h1 ? _GEN_730 : _GEN_3420; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3805 = unuse_way == 2'h1 ? _GEN_731 : _GEN_3421; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3806 = unuse_way == 2'h1 ? _GEN_732 : _GEN_3422; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3807 = unuse_way == 2'h1 ? _GEN_733 : _GEN_3423; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3808 = unuse_way == 2'h1 ? _GEN_734 : _GEN_3424; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3809 = unuse_way == 2'h1 ? _GEN_735 : _GEN_3425; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3810 = unuse_way == 2'h1 ? _GEN_736 : _GEN_3426; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3811 = unuse_way == 2'h1 ? _GEN_737 : _GEN_3427; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3812 = unuse_way == 2'h1 ? _GEN_738 : _GEN_3428; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3813 = unuse_way == 2'h1 ? _GEN_739 : _GEN_3429; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3814 = unuse_way == 2'h1 ? _GEN_740 : _GEN_3430; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3815 = unuse_way == 2'h1 ? _GEN_741 : _GEN_3431; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3816 = unuse_way == 2'h1 ? _GEN_742 : _GEN_3432; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3817 = unuse_way == 2'h1 ? _GEN_743 : _GEN_3433; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3818 = unuse_way == 2'h1 ? _GEN_744 : _GEN_3434; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3819 = unuse_way == 2'h1 ? _GEN_745 : _GEN_3435; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3820 = unuse_way == 2'h1 ? _GEN_746 : _GEN_3436; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3821 = unuse_way == 2'h1 ? _GEN_747 : _GEN_3437; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3822 = unuse_way == 2'h1 ? _GEN_748 : _GEN_3438; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3823 = unuse_way == 2'h1 ? _GEN_749 : _GEN_3439; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3824 = unuse_way == 2'h1 ? _GEN_750 : _GEN_3440; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3825 = unuse_way == 2'h1 ? _GEN_751 : _GEN_3441; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3826 = unuse_way == 2'h1 ? _GEN_752 : _GEN_3442; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3827 = unuse_way == 2'h1 ? _GEN_753 : _GEN_3443; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3828 = unuse_way == 2'h1 ? _GEN_754 : _GEN_3444; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3829 = unuse_way == 2'h1 ? _GEN_755 : _GEN_3445; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3830 = unuse_way == 2'h1 ? _GEN_756 : _GEN_3446; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3831 = unuse_way == 2'h1 ? _GEN_757 : _GEN_3447; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3832 = unuse_way == 2'h1 ? _GEN_758 : _GEN_3448; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3833 = unuse_way == 2'h1 ? _GEN_759 : _GEN_3449; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3834 = unuse_way == 2'h1 ? _GEN_760 : _GEN_3450; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3835 = unuse_way == 2'h1 ? _GEN_761 : _GEN_3451; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3836 = unuse_way == 2'h1 ? _GEN_762 : _GEN_3452; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3837 = unuse_way == 2'h1 ? _GEN_763 : _GEN_3453; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3838 = unuse_way == 2'h1 ? _GEN_764 : _GEN_3454; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3839 = unuse_way == 2'h1 ? _GEN_765 : _GEN_3455; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3840 = unuse_way == 2'h1 ? _GEN_766 : _GEN_3456; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3841 = unuse_way == 2'h1 ? _GEN_767 : _GEN_3457; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3842 = unuse_way == 2'h1 ? _GEN_768 : _GEN_3458; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3843 = unuse_way == 2'h1 ? _GEN_769 : _GEN_3459; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3844 = unuse_way == 2'h1 ? _GEN_770 : _GEN_3460; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3845 = unuse_way == 2'h1 ? _GEN_771 : _GEN_3461; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3846 = unuse_way == 2'h1 ? _GEN_772 : _GEN_3462; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3847 = unuse_way == 2'h1 ? _GEN_773 : _GEN_3463; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3848 = unuse_way == 2'h1 ? _GEN_774 : _GEN_3464; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3849 = unuse_way == 2'h1 ? _GEN_775 : _GEN_3465; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3850 = unuse_way == 2'h1 ? _GEN_776 : _GEN_3466; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3851 = unuse_way == 2'h1 ? _GEN_777 : _GEN_3467; // @[i_cache.scala 86:34]
  wire  _GEN_3852 = unuse_way == 2'h1 ? _GEN_778 : _GEN_3468; // @[i_cache.scala 86:34]
  wire  _GEN_3853 = unuse_way == 2'h1 ? _GEN_779 : _GEN_3469; // @[i_cache.scala 86:34]
  wire  _GEN_3854 = unuse_way == 2'h1 ? _GEN_780 : _GEN_3470; // @[i_cache.scala 86:34]
  wire  _GEN_3855 = unuse_way == 2'h1 ? _GEN_781 : _GEN_3471; // @[i_cache.scala 86:34]
  wire  _GEN_3856 = unuse_way == 2'h1 ? _GEN_782 : _GEN_3472; // @[i_cache.scala 86:34]
  wire  _GEN_3857 = unuse_way == 2'h1 ? _GEN_783 : _GEN_3473; // @[i_cache.scala 86:34]
  wire  _GEN_3858 = unuse_way == 2'h1 ? _GEN_784 : _GEN_3474; // @[i_cache.scala 86:34]
  wire  _GEN_3859 = unuse_way == 2'h1 ? _GEN_785 : _GEN_3475; // @[i_cache.scala 86:34]
  wire  _GEN_3860 = unuse_way == 2'h1 ? _GEN_786 : _GEN_3476; // @[i_cache.scala 86:34]
  wire  _GEN_3861 = unuse_way == 2'h1 ? _GEN_787 : _GEN_3477; // @[i_cache.scala 86:34]
  wire  _GEN_3862 = unuse_way == 2'h1 ? _GEN_788 : _GEN_3478; // @[i_cache.scala 86:34]
  wire  _GEN_3863 = unuse_way == 2'h1 ? _GEN_789 : _GEN_3479; // @[i_cache.scala 86:34]
  wire  _GEN_3864 = unuse_way == 2'h1 ? _GEN_790 : _GEN_3480; // @[i_cache.scala 86:34]
  wire  _GEN_3865 = unuse_way == 2'h1 ? _GEN_791 : _GEN_3481; // @[i_cache.scala 86:34]
  wire  _GEN_3866 = unuse_way == 2'h1 ? _GEN_792 : _GEN_3482; // @[i_cache.scala 86:34]
  wire  _GEN_3867 = unuse_way == 2'h1 ? _GEN_793 : _GEN_3483; // @[i_cache.scala 86:34]
  wire  _GEN_3868 = unuse_way == 2'h1 ? _GEN_794 : _GEN_3484; // @[i_cache.scala 86:34]
  wire  _GEN_3869 = unuse_way == 2'h1 ? _GEN_795 : _GEN_3485; // @[i_cache.scala 86:34]
  wire  _GEN_3870 = unuse_way == 2'h1 ? _GEN_796 : _GEN_3486; // @[i_cache.scala 86:34]
  wire  _GEN_3871 = unuse_way == 2'h1 ? _GEN_797 : _GEN_3487; // @[i_cache.scala 86:34]
  wire  _GEN_3872 = unuse_way == 2'h1 ? _GEN_798 : _GEN_3488; // @[i_cache.scala 86:34]
  wire  _GEN_3873 = unuse_way == 2'h1 ? _GEN_799 : _GEN_3489; // @[i_cache.scala 86:34]
  wire  _GEN_3874 = unuse_way == 2'h1 ? _GEN_800 : _GEN_3490; // @[i_cache.scala 86:34]
  wire  _GEN_3875 = unuse_way == 2'h1 ? _GEN_801 : _GEN_3491; // @[i_cache.scala 86:34]
  wire  _GEN_3876 = unuse_way == 2'h1 ? _GEN_802 : _GEN_3492; // @[i_cache.scala 86:34]
  wire  _GEN_3877 = unuse_way == 2'h1 ? _GEN_803 : _GEN_3493; // @[i_cache.scala 86:34]
  wire  _GEN_3878 = unuse_way == 2'h1 ? _GEN_804 : _GEN_3494; // @[i_cache.scala 86:34]
  wire  _GEN_3879 = unuse_way == 2'h1 ? _GEN_805 : _GEN_3495; // @[i_cache.scala 86:34]
  wire  _GEN_3880 = unuse_way == 2'h1 ? _GEN_806 : _GEN_3496; // @[i_cache.scala 86:34]
  wire  _GEN_3881 = unuse_way == 2'h1 ? _GEN_807 : _GEN_3497; // @[i_cache.scala 86:34]
  wire  _GEN_3882 = unuse_way == 2'h1 ? _GEN_808 : _GEN_3498; // @[i_cache.scala 86:34]
  wire  _GEN_3883 = unuse_way == 2'h1 ? _GEN_809 : _GEN_3499; // @[i_cache.scala 86:34]
  wire  _GEN_3884 = unuse_way == 2'h1 ? _GEN_810 : _GEN_3500; // @[i_cache.scala 86:34]
  wire  _GEN_3885 = unuse_way == 2'h1 ? _GEN_811 : _GEN_3501; // @[i_cache.scala 86:34]
  wire  _GEN_3886 = unuse_way == 2'h1 ? _GEN_812 : _GEN_3502; // @[i_cache.scala 86:34]
  wire  _GEN_3887 = unuse_way == 2'h1 ? _GEN_813 : _GEN_3503; // @[i_cache.scala 86:34]
  wire  _GEN_3888 = unuse_way == 2'h1 ? _GEN_814 : _GEN_3504; // @[i_cache.scala 86:34]
  wire  _GEN_3889 = unuse_way == 2'h1 ? _GEN_815 : _GEN_3505; // @[i_cache.scala 86:34]
  wire  _GEN_3890 = unuse_way == 2'h1 ? _GEN_816 : _GEN_3506; // @[i_cache.scala 86:34]
  wire  _GEN_3891 = unuse_way == 2'h1 ? _GEN_817 : _GEN_3507; // @[i_cache.scala 86:34]
  wire  _GEN_3892 = unuse_way == 2'h1 ? _GEN_818 : _GEN_3508; // @[i_cache.scala 86:34]
  wire  _GEN_3893 = unuse_way == 2'h1 ? _GEN_819 : _GEN_3509; // @[i_cache.scala 86:34]
  wire  _GEN_3894 = unuse_way == 2'h1 ? _GEN_820 : _GEN_3510; // @[i_cache.scala 86:34]
  wire  _GEN_3895 = unuse_way == 2'h1 ? _GEN_821 : _GEN_3511; // @[i_cache.scala 86:34]
  wire  _GEN_3896 = unuse_way == 2'h1 ? _GEN_822 : _GEN_3512; // @[i_cache.scala 86:34]
  wire  _GEN_3897 = unuse_way == 2'h1 ? _GEN_823 : _GEN_3513; // @[i_cache.scala 86:34]
  wire  _GEN_3898 = unuse_way == 2'h1 ? _GEN_824 : _GEN_3514; // @[i_cache.scala 86:34]
  wire  _GEN_3899 = unuse_way == 2'h1 ? _GEN_825 : _GEN_3515; // @[i_cache.scala 86:34]
  wire  _GEN_3900 = unuse_way == 2'h1 ? _GEN_826 : _GEN_3516; // @[i_cache.scala 86:34]
  wire  _GEN_3901 = unuse_way == 2'h1 ? _GEN_827 : _GEN_3517; // @[i_cache.scala 86:34]
  wire  _GEN_3902 = unuse_way == 2'h1 ? _GEN_828 : _GEN_3518; // @[i_cache.scala 86:34]
  wire  _GEN_3903 = unuse_way == 2'h1 ? _GEN_829 : _GEN_3519; // @[i_cache.scala 86:34]
  wire  _GEN_3904 = unuse_way == 2'h1 ? _GEN_830 : _GEN_3520; // @[i_cache.scala 86:34]
  wire  _GEN_3905 = unuse_way == 2'h1 ? _GEN_831 : _GEN_3521; // @[i_cache.scala 86:34]
  wire  _GEN_3906 = unuse_way == 2'h1 ? _GEN_832 : _GEN_3522; // @[i_cache.scala 86:34]
  wire  _GEN_3907 = unuse_way == 2'h1 ? _GEN_833 : _GEN_3523; // @[i_cache.scala 86:34]
  wire  _GEN_3908 = unuse_way == 2'h1 ? _GEN_834 : _GEN_3524; // @[i_cache.scala 86:34]
  wire  _GEN_3909 = unuse_way == 2'h1 ? _GEN_835 : _GEN_3525; // @[i_cache.scala 86:34]
  wire  _GEN_3910 = unuse_way == 2'h1 ? _GEN_836 : _GEN_3526; // @[i_cache.scala 86:34]
  wire  _GEN_3911 = unuse_way == 2'h1 ? _GEN_837 : _GEN_3527; // @[i_cache.scala 86:34]
  wire  _GEN_3912 = unuse_way == 2'h1 ? _GEN_838 : _GEN_3528; // @[i_cache.scala 86:34]
  wire  _GEN_3913 = unuse_way == 2'h1 ? _GEN_839 : _GEN_3529; // @[i_cache.scala 86:34]
  wire  _GEN_3914 = unuse_way == 2'h1 ? _GEN_840 : _GEN_3530; // @[i_cache.scala 86:34]
  wire  _GEN_3915 = unuse_way == 2'h1 ? _GEN_841 : _GEN_3531; // @[i_cache.scala 86:34]
  wire  _GEN_3916 = unuse_way == 2'h1 ? _GEN_842 : _GEN_3532; // @[i_cache.scala 86:34]
  wire  _GEN_3917 = unuse_way == 2'h1 ? _GEN_843 : _GEN_3533; // @[i_cache.scala 86:34]
  wire  _GEN_3918 = unuse_way == 2'h1 ? _GEN_844 : _GEN_3534; // @[i_cache.scala 86:34]
  wire  _GEN_3919 = unuse_way == 2'h1 ? _GEN_845 : _GEN_3535; // @[i_cache.scala 86:34]
  wire  _GEN_3920 = unuse_way == 2'h1 ? _GEN_846 : _GEN_3536; // @[i_cache.scala 86:34]
  wire  _GEN_3921 = unuse_way == 2'h1 ? _GEN_847 : _GEN_3537; // @[i_cache.scala 86:34]
  wire  _GEN_3922 = unuse_way == 2'h1 ? _GEN_848 : _GEN_3538; // @[i_cache.scala 86:34]
  wire  _GEN_3923 = unuse_way == 2'h1 ? _GEN_849 : _GEN_3539; // @[i_cache.scala 86:34]
  wire  _GEN_3924 = unuse_way == 2'h1 ? _GEN_850 : _GEN_3540; // @[i_cache.scala 86:34]
  wire  _GEN_3925 = unuse_way == 2'h1 ? _GEN_851 : _GEN_3541; // @[i_cache.scala 86:34]
  wire  _GEN_3926 = unuse_way == 2'h1 ? _GEN_852 : _GEN_3542; // @[i_cache.scala 86:34]
  wire  _GEN_3927 = unuse_way == 2'h1 ? _GEN_853 : _GEN_3543; // @[i_cache.scala 86:34]
  wire  _GEN_3928 = unuse_way == 2'h1 ? _GEN_854 : _GEN_3544; // @[i_cache.scala 86:34]
  wire  _GEN_3929 = unuse_way == 2'h1 ? _GEN_855 : _GEN_3545; // @[i_cache.scala 86:34]
  wire  _GEN_3930 = unuse_way == 2'h1 ? _GEN_856 : _GEN_3546; // @[i_cache.scala 86:34]
  wire  _GEN_3931 = unuse_way == 2'h1 ? _GEN_857 : _GEN_3547; // @[i_cache.scala 86:34]
  wire  _GEN_3932 = unuse_way == 2'h1 ? _GEN_858 : _GEN_3548; // @[i_cache.scala 86:34]
  wire  _GEN_3933 = unuse_way == 2'h1 ? _GEN_859 : _GEN_3549; // @[i_cache.scala 86:34]
  wire  _GEN_3934 = unuse_way == 2'h1 ? _GEN_860 : _GEN_3550; // @[i_cache.scala 86:34]
  wire  _GEN_3935 = unuse_way == 2'h1 ? _GEN_861 : _GEN_3551; // @[i_cache.scala 86:34]
  wire  _GEN_3936 = unuse_way == 2'h1 ? _GEN_862 : _GEN_3552; // @[i_cache.scala 86:34]
  wire  _GEN_3937 = unuse_way == 2'h1 ? _GEN_863 : _GEN_3553; // @[i_cache.scala 86:34]
  wire  _GEN_3938 = unuse_way == 2'h1 ? _GEN_864 : _GEN_3554; // @[i_cache.scala 86:34]
  wire  _GEN_3939 = unuse_way == 2'h1 ? _GEN_865 : _GEN_3555; // @[i_cache.scala 86:34]
  wire  _GEN_3940 = unuse_way == 2'h1 ? _GEN_866 : _GEN_3556; // @[i_cache.scala 86:34]
  wire  _GEN_3941 = unuse_way == 2'h1 ? _GEN_867 : _GEN_3557; // @[i_cache.scala 86:34]
  wire  _GEN_3942 = unuse_way == 2'h1 ? _GEN_868 : _GEN_3558; // @[i_cache.scala 86:34]
  wire  _GEN_3943 = unuse_way == 2'h1 ? _GEN_869 : _GEN_3559; // @[i_cache.scala 86:34]
  wire  _GEN_3944 = unuse_way == 2'h1 ? _GEN_870 : _GEN_3560; // @[i_cache.scala 86:34]
  wire  _GEN_3945 = unuse_way == 2'h1 ? _GEN_871 : _GEN_3561; // @[i_cache.scala 86:34]
  wire  _GEN_3946 = unuse_way == 2'h1 ? _GEN_872 : _GEN_3562; // @[i_cache.scala 86:34]
  wire  _GEN_3947 = unuse_way == 2'h1 ? _GEN_873 : _GEN_3563; // @[i_cache.scala 86:34]
  wire  _GEN_3948 = unuse_way == 2'h1 ? _GEN_874 : _GEN_3564; // @[i_cache.scala 86:34]
  wire  _GEN_3949 = unuse_way == 2'h1 ? _GEN_875 : _GEN_3565; // @[i_cache.scala 86:34]
  wire  _GEN_3950 = unuse_way == 2'h1 ? _GEN_876 : _GEN_3566; // @[i_cache.scala 86:34]
  wire  _GEN_3951 = unuse_way == 2'h1 ? _GEN_877 : _GEN_3567; // @[i_cache.scala 86:34]
  wire  _GEN_3952 = unuse_way == 2'h1 ? _GEN_878 : _GEN_3568; // @[i_cache.scala 86:34]
  wire  _GEN_3953 = unuse_way == 2'h1 ? _GEN_879 : _GEN_3569; // @[i_cache.scala 86:34]
  wire  _GEN_3954 = unuse_way == 2'h1 ? _GEN_880 : _GEN_3570; // @[i_cache.scala 86:34]
  wire  _GEN_3955 = unuse_way == 2'h1 ? _GEN_881 : _GEN_3571; // @[i_cache.scala 86:34]
  wire  _GEN_3956 = unuse_way == 2'h1 ? _GEN_882 : _GEN_3572; // @[i_cache.scala 86:34]
  wire  _GEN_3957 = unuse_way == 2'h1 ? _GEN_883 : _GEN_3573; // @[i_cache.scala 86:34]
  wire  _GEN_3958 = unuse_way == 2'h1 ? _GEN_884 : _GEN_3574; // @[i_cache.scala 86:34]
  wire  _GEN_3959 = unuse_way == 2'h1 ? _GEN_885 : _GEN_3575; // @[i_cache.scala 86:34]
  wire  _GEN_3960 = unuse_way == 2'h1 ? _GEN_886 : _GEN_3576; // @[i_cache.scala 86:34]
  wire  _GEN_3961 = unuse_way == 2'h1 ? _GEN_887 : _GEN_3577; // @[i_cache.scala 86:34]
  wire  _GEN_3962 = unuse_way == 2'h1 ? _GEN_888 : _GEN_3578; // @[i_cache.scala 86:34]
  wire  _GEN_3963 = unuse_way == 2'h1 ? _GEN_889 : _GEN_3579; // @[i_cache.scala 86:34]
  wire  _GEN_3964 = unuse_way == 2'h1 ? _GEN_890 : _GEN_3580; // @[i_cache.scala 86:34]
  wire  _GEN_3965 = unuse_way == 2'h1 ? _GEN_891 : _GEN_3581; // @[i_cache.scala 86:34]
  wire  _GEN_3966 = unuse_way == 2'h1 ? _GEN_892 : _GEN_3582; // @[i_cache.scala 86:34]
  wire  _GEN_3967 = unuse_way == 2'h1 ? _GEN_893 : _GEN_3583; // @[i_cache.scala 86:34]
  wire  _GEN_3968 = unuse_way == 2'h1 ? _GEN_894 : _GEN_3584; // @[i_cache.scala 86:34]
  wire  _GEN_3969 = unuse_way == 2'h1 ? _GEN_895 : _GEN_3585; // @[i_cache.scala 86:34]
  wire  _GEN_3970 = unuse_way == 2'h1 ? _GEN_896 : _GEN_3586; // @[i_cache.scala 86:34]
  wire  _GEN_3971 = unuse_way == 2'h1 ? _GEN_897 : _GEN_3587; // @[i_cache.scala 86:34]
  wire  _GEN_3972 = unuse_way == 2'h1 ? _GEN_898 : _GEN_3588; // @[i_cache.scala 86:34]
  wire  _GEN_3973 = unuse_way == 2'h1 ? _GEN_899 : _GEN_3589; // @[i_cache.scala 86:34]
  wire  _GEN_3974 = unuse_way == 2'h1 ? _GEN_900 : _GEN_3590; // @[i_cache.scala 86:34]
  wire  _GEN_3975 = unuse_way == 2'h1 ? _GEN_901 : _GEN_3591; // @[i_cache.scala 86:34]
  wire  _GEN_3976 = unuse_way == 2'h1 ? _GEN_902 : _GEN_3592; // @[i_cache.scala 86:34]
  wire  _GEN_3977 = unuse_way == 2'h1 ? _GEN_903 : _GEN_3593; // @[i_cache.scala 86:34]
  wire  _GEN_3978 = unuse_way == 2'h1 ? _GEN_904 : _GEN_3594; // @[i_cache.scala 86:34]
  wire  _GEN_3979 = unuse_way == 2'h1 ? _GEN_905 : _GEN_3595; // @[i_cache.scala 86:34]
  wire  _GEN_3980 = unuse_way == 2'h1 | _GEN_3211; // @[i_cache.scala 86:34 90:23]
  wire [63:0] _GEN_3981 = unuse_way == 2'h1 ? ram_1_0 : _GEN_2827; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3982 = unuse_way == 2'h1 ? ram_1_1 : _GEN_2828; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3983 = unuse_way == 2'h1 ? ram_1_2 : _GEN_2829; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3984 = unuse_way == 2'h1 ? ram_1_3 : _GEN_2830; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3985 = unuse_way == 2'h1 ? ram_1_4 : _GEN_2831; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3986 = unuse_way == 2'h1 ? ram_1_5 : _GEN_2832; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3987 = unuse_way == 2'h1 ? ram_1_6 : _GEN_2833; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3988 = unuse_way == 2'h1 ? ram_1_7 : _GEN_2834; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3989 = unuse_way == 2'h1 ? ram_1_8 : _GEN_2835; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3990 = unuse_way == 2'h1 ? ram_1_9 : _GEN_2836; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3991 = unuse_way == 2'h1 ? ram_1_10 : _GEN_2837; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3992 = unuse_way == 2'h1 ? ram_1_11 : _GEN_2838; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3993 = unuse_way == 2'h1 ? ram_1_12 : _GEN_2839; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3994 = unuse_way == 2'h1 ? ram_1_13 : _GEN_2840; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3995 = unuse_way == 2'h1 ? ram_1_14 : _GEN_2841; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3996 = unuse_way == 2'h1 ? ram_1_15 : _GEN_2842; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3997 = unuse_way == 2'h1 ? ram_1_16 : _GEN_2843; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3998 = unuse_way == 2'h1 ? ram_1_17 : _GEN_2844; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3999 = unuse_way == 2'h1 ? ram_1_18 : _GEN_2845; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4000 = unuse_way == 2'h1 ? ram_1_19 : _GEN_2846; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4001 = unuse_way == 2'h1 ? ram_1_20 : _GEN_2847; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4002 = unuse_way == 2'h1 ? ram_1_21 : _GEN_2848; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4003 = unuse_way == 2'h1 ? ram_1_22 : _GEN_2849; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4004 = unuse_way == 2'h1 ? ram_1_23 : _GEN_2850; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4005 = unuse_way == 2'h1 ? ram_1_24 : _GEN_2851; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4006 = unuse_way == 2'h1 ? ram_1_25 : _GEN_2852; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4007 = unuse_way == 2'h1 ? ram_1_26 : _GEN_2853; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4008 = unuse_way == 2'h1 ? ram_1_27 : _GEN_2854; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4009 = unuse_way == 2'h1 ? ram_1_28 : _GEN_2855; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4010 = unuse_way == 2'h1 ? ram_1_29 : _GEN_2856; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4011 = unuse_way == 2'h1 ? ram_1_30 : _GEN_2857; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4012 = unuse_way == 2'h1 ? ram_1_31 : _GEN_2858; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4013 = unuse_way == 2'h1 ? ram_1_32 : _GEN_2859; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4014 = unuse_way == 2'h1 ? ram_1_33 : _GEN_2860; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4015 = unuse_way == 2'h1 ? ram_1_34 : _GEN_2861; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4016 = unuse_way == 2'h1 ? ram_1_35 : _GEN_2862; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4017 = unuse_way == 2'h1 ? ram_1_36 : _GEN_2863; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4018 = unuse_way == 2'h1 ? ram_1_37 : _GEN_2864; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4019 = unuse_way == 2'h1 ? ram_1_38 : _GEN_2865; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4020 = unuse_way == 2'h1 ? ram_1_39 : _GEN_2866; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4021 = unuse_way == 2'h1 ? ram_1_40 : _GEN_2867; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4022 = unuse_way == 2'h1 ? ram_1_41 : _GEN_2868; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4023 = unuse_way == 2'h1 ? ram_1_42 : _GEN_2869; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4024 = unuse_way == 2'h1 ? ram_1_43 : _GEN_2870; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4025 = unuse_way == 2'h1 ? ram_1_44 : _GEN_2871; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4026 = unuse_way == 2'h1 ? ram_1_45 : _GEN_2872; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4027 = unuse_way == 2'h1 ? ram_1_46 : _GEN_2873; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4028 = unuse_way == 2'h1 ? ram_1_47 : _GEN_2874; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4029 = unuse_way == 2'h1 ? ram_1_48 : _GEN_2875; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4030 = unuse_way == 2'h1 ? ram_1_49 : _GEN_2876; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4031 = unuse_way == 2'h1 ? ram_1_50 : _GEN_2877; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4032 = unuse_way == 2'h1 ? ram_1_51 : _GEN_2878; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4033 = unuse_way == 2'h1 ? ram_1_52 : _GEN_2879; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4034 = unuse_way == 2'h1 ? ram_1_53 : _GEN_2880; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4035 = unuse_way == 2'h1 ? ram_1_54 : _GEN_2881; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4036 = unuse_way == 2'h1 ? ram_1_55 : _GEN_2882; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4037 = unuse_way == 2'h1 ? ram_1_56 : _GEN_2883; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4038 = unuse_way == 2'h1 ? ram_1_57 : _GEN_2884; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4039 = unuse_way == 2'h1 ? ram_1_58 : _GEN_2885; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4040 = unuse_way == 2'h1 ? ram_1_59 : _GEN_2886; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4041 = unuse_way == 2'h1 ? ram_1_60 : _GEN_2887; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4042 = unuse_way == 2'h1 ? ram_1_61 : _GEN_2888; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4043 = unuse_way == 2'h1 ? ram_1_62 : _GEN_2889; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4044 = unuse_way == 2'h1 ? ram_1_63 : _GEN_2890; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4045 = unuse_way == 2'h1 ? ram_1_64 : _GEN_2891; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4046 = unuse_way == 2'h1 ? ram_1_65 : _GEN_2892; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4047 = unuse_way == 2'h1 ? ram_1_66 : _GEN_2893; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4048 = unuse_way == 2'h1 ? ram_1_67 : _GEN_2894; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4049 = unuse_way == 2'h1 ? ram_1_68 : _GEN_2895; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4050 = unuse_way == 2'h1 ? ram_1_69 : _GEN_2896; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4051 = unuse_way == 2'h1 ? ram_1_70 : _GEN_2897; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4052 = unuse_way == 2'h1 ? ram_1_71 : _GEN_2898; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4053 = unuse_way == 2'h1 ? ram_1_72 : _GEN_2899; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4054 = unuse_way == 2'h1 ? ram_1_73 : _GEN_2900; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4055 = unuse_way == 2'h1 ? ram_1_74 : _GEN_2901; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4056 = unuse_way == 2'h1 ? ram_1_75 : _GEN_2902; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4057 = unuse_way == 2'h1 ? ram_1_76 : _GEN_2903; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4058 = unuse_way == 2'h1 ? ram_1_77 : _GEN_2904; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4059 = unuse_way == 2'h1 ? ram_1_78 : _GEN_2905; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4060 = unuse_way == 2'h1 ? ram_1_79 : _GEN_2906; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4061 = unuse_way == 2'h1 ? ram_1_80 : _GEN_2907; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4062 = unuse_way == 2'h1 ? ram_1_81 : _GEN_2908; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4063 = unuse_way == 2'h1 ? ram_1_82 : _GEN_2909; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4064 = unuse_way == 2'h1 ? ram_1_83 : _GEN_2910; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4065 = unuse_way == 2'h1 ? ram_1_84 : _GEN_2911; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4066 = unuse_way == 2'h1 ? ram_1_85 : _GEN_2912; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4067 = unuse_way == 2'h1 ? ram_1_86 : _GEN_2913; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4068 = unuse_way == 2'h1 ? ram_1_87 : _GEN_2914; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4069 = unuse_way == 2'h1 ? ram_1_88 : _GEN_2915; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4070 = unuse_way == 2'h1 ? ram_1_89 : _GEN_2916; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4071 = unuse_way == 2'h1 ? ram_1_90 : _GEN_2917; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4072 = unuse_way == 2'h1 ? ram_1_91 : _GEN_2918; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4073 = unuse_way == 2'h1 ? ram_1_92 : _GEN_2919; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4074 = unuse_way == 2'h1 ? ram_1_93 : _GEN_2920; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4075 = unuse_way == 2'h1 ? ram_1_94 : _GEN_2921; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4076 = unuse_way == 2'h1 ? ram_1_95 : _GEN_2922; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4077 = unuse_way == 2'h1 ? ram_1_96 : _GEN_2923; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4078 = unuse_way == 2'h1 ? ram_1_97 : _GEN_2924; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4079 = unuse_way == 2'h1 ? ram_1_98 : _GEN_2925; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4080 = unuse_way == 2'h1 ? ram_1_99 : _GEN_2926; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4081 = unuse_way == 2'h1 ? ram_1_100 : _GEN_2927; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4082 = unuse_way == 2'h1 ? ram_1_101 : _GEN_2928; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4083 = unuse_way == 2'h1 ? ram_1_102 : _GEN_2929; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4084 = unuse_way == 2'h1 ? ram_1_103 : _GEN_2930; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4085 = unuse_way == 2'h1 ? ram_1_104 : _GEN_2931; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4086 = unuse_way == 2'h1 ? ram_1_105 : _GEN_2932; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4087 = unuse_way == 2'h1 ? ram_1_106 : _GEN_2933; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4088 = unuse_way == 2'h1 ? ram_1_107 : _GEN_2934; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4089 = unuse_way == 2'h1 ? ram_1_108 : _GEN_2935; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4090 = unuse_way == 2'h1 ? ram_1_109 : _GEN_2936; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4091 = unuse_way == 2'h1 ? ram_1_110 : _GEN_2937; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4092 = unuse_way == 2'h1 ? ram_1_111 : _GEN_2938; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4093 = unuse_way == 2'h1 ? ram_1_112 : _GEN_2939; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4094 = unuse_way == 2'h1 ? ram_1_113 : _GEN_2940; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4095 = unuse_way == 2'h1 ? ram_1_114 : _GEN_2941; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4096 = unuse_way == 2'h1 ? ram_1_115 : _GEN_2942; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4097 = unuse_way == 2'h1 ? ram_1_116 : _GEN_2943; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4098 = unuse_way == 2'h1 ? ram_1_117 : _GEN_2944; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4099 = unuse_way == 2'h1 ? ram_1_118 : _GEN_2945; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4100 = unuse_way == 2'h1 ? ram_1_119 : _GEN_2946; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4101 = unuse_way == 2'h1 ? ram_1_120 : _GEN_2947; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4102 = unuse_way == 2'h1 ? ram_1_121 : _GEN_2948; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4103 = unuse_way == 2'h1 ? ram_1_122 : _GEN_2949; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4104 = unuse_way == 2'h1 ? ram_1_123 : _GEN_2950; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4105 = unuse_way == 2'h1 ? ram_1_124 : _GEN_2951; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4106 = unuse_way == 2'h1 ? ram_1_125 : _GEN_2952; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4107 = unuse_way == 2'h1 ? ram_1_126 : _GEN_2953; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4108 = unuse_way == 2'h1 ? ram_1_127 : _GEN_2954; // @[i_cache.scala 18:24 86:34]
  wire [31:0] _GEN_4109 = unuse_way == 2'h1 ? tag_1_0 : _GEN_2955; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4110 = unuse_way == 2'h1 ? tag_1_1 : _GEN_2956; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4111 = unuse_way == 2'h1 ? tag_1_2 : _GEN_2957; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4112 = unuse_way == 2'h1 ? tag_1_3 : _GEN_2958; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4113 = unuse_way == 2'h1 ? tag_1_4 : _GEN_2959; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4114 = unuse_way == 2'h1 ? tag_1_5 : _GEN_2960; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4115 = unuse_way == 2'h1 ? tag_1_6 : _GEN_2961; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4116 = unuse_way == 2'h1 ? tag_1_7 : _GEN_2962; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4117 = unuse_way == 2'h1 ? tag_1_8 : _GEN_2963; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4118 = unuse_way == 2'h1 ? tag_1_9 : _GEN_2964; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4119 = unuse_way == 2'h1 ? tag_1_10 : _GEN_2965; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4120 = unuse_way == 2'h1 ? tag_1_11 : _GEN_2966; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4121 = unuse_way == 2'h1 ? tag_1_12 : _GEN_2967; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4122 = unuse_way == 2'h1 ? tag_1_13 : _GEN_2968; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4123 = unuse_way == 2'h1 ? tag_1_14 : _GEN_2969; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4124 = unuse_way == 2'h1 ? tag_1_15 : _GEN_2970; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4125 = unuse_way == 2'h1 ? tag_1_16 : _GEN_2971; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4126 = unuse_way == 2'h1 ? tag_1_17 : _GEN_2972; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4127 = unuse_way == 2'h1 ? tag_1_18 : _GEN_2973; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4128 = unuse_way == 2'h1 ? tag_1_19 : _GEN_2974; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4129 = unuse_way == 2'h1 ? tag_1_20 : _GEN_2975; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4130 = unuse_way == 2'h1 ? tag_1_21 : _GEN_2976; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4131 = unuse_way == 2'h1 ? tag_1_22 : _GEN_2977; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4132 = unuse_way == 2'h1 ? tag_1_23 : _GEN_2978; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4133 = unuse_way == 2'h1 ? tag_1_24 : _GEN_2979; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4134 = unuse_way == 2'h1 ? tag_1_25 : _GEN_2980; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4135 = unuse_way == 2'h1 ? tag_1_26 : _GEN_2981; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4136 = unuse_way == 2'h1 ? tag_1_27 : _GEN_2982; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4137 = unuse_way == 2'h1 ? tag_1_28 : _GEN_2983; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4138 = unuse_way == 2'h1 ? tag_1_29 : _GEN_2984; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4139 = unuse_way == 2'h1 ? tag_1_30 : _GEN_2985; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4140 = unuse_way == 2'h1 ? tag_1_31 : _GEN_2986; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4141 = unuse_way == 2'h1 ? tag_1_32 : _GEN_2987; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4142 = unuse_way == 2'h1 ? tag_1_33 : _GEN_2988; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4143 = unuse_way == 2'h1 ? tag_1_34 : _GEN_2989; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4144 = unuse_way == 2'h1 ? tag_1_35 : _GEN_2990; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4145 = unuse_way == 2'h1 ? tag_1_36 : _GEN_2991; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4146 = unuse_way == 2'h1 ? tag_1_37 : _GEN_2992; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4147 = unuse_way == 2'h1 ? tag_1_38 : _GEN_2993; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4148 = unuse_way == 2'h1 ? tag_1_39 : _GEN_2994; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4149 = unuse_way == 2'h1 ? tag_1_40 : _GEN_2995; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4150 = unuse_way == 2'h1 ? tag_1_41 : _GEN_2996; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4151 = unuse_way == 2'h1 ? tag_1_42 : _GEN_2997; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4152 = unuse_way == 2'h1 ? tag_1_43 : _GEN_2998; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4153 = unuse_way == 2'h1 ? tag_1_44 : _GEN_2999; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4154 = unuse_way == 2'h1 ? tag_1_45 : _GEN_3000; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4155 = unuse_way == 2'h1 ? tag_1_46 : _GEN_3001; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4156 = unuse_way == 2'h1 ? tag_1_47 : _GEN_3002; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4157 = unuse_way == 2'h1 ? tag_1_48 : _GEN_3003; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4158 = unuse_way == 2'h1 ? tag_1_49 : _GEN_3004; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4159 = unuse_way == 2'h1 ? tag_1_50 : _GEN_3005; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4160 = unuse_way == 2'h1 ? tag_1_51 : _GEN_3006; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4161 = unuse_way == 2'h1 ? tag_1_52 : _GEN_3007; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4162 = unuse_way == 2'h1 ? tag_1_53 : _GEN_3008; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4163 = unuse_way == 2'h1 ? tag_1_54 : _GEN_3009; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4164 = unuse_way == 2'h1 ? tag_1_55 : _GEN_3010; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4165 = unuse_way == 2'h1 ? tag_1_56 : _GEN_3011; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4166 = unuse_way == 2'h1 ? tag_1_57 : _GEN_3012; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4167 = unuse_way == 2'h1 ? tag_1_58 : _GEN_3013; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4168 = unuse_way == 2'h1 ? tag_1_59 : _GEN_3014; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4169 = unuse_way == 2'h1 ? tag_1_60 : _GEN_3015; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4170 = unuse_way == 2'h1 ? tag_1_61 : _GEN_3016; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4171 = unuse_way == 2'h1 ? tag_1_62 : _GEN_3017; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4172 = unuse_way == 2'h1 ? tag_1_63 : _GEN_3018; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4173 = unuse_way == 2'h1 ? tag_1_64 : _GEN_3019; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4174 = unuse_way == 2'h1 ? tag_1_65 : _GEN_3020; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4175 = unuse_way == 2'h1 ? tag_1_66 : _GEN_3021; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4176 = unuse_way == 2'h1 ? tag_1_67 : _GEN_3022; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4177 = unuse_way == 2'h1 ? tag_1_68 : _GEN_3023; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4178 = unuse_way == 2'h1 ? tag_1_69 : _GEN_3024; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4179 = unuse_way == 2'h1 ? tag_1_70 : _GEN_3025; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4180 = unuse_way == 2'h1 ? tag_1_71 : _GEN_3026; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4181 = unuse_way == 2'h1 ? tag_1_72 : _GEN_3027; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4182 = unuse_way == 2'h1 ? tag_1_73 : _GEN_3028; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4183 = unuse_way == 2'h1 ? tag_1_74 : _GEN_3029; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4184 = unuse_way == 2'h1 ? tag_1_75 : _GEN_3030; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4185 = unuse_way == 2'h1 ? tag_1_76 : _GEN_3031; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4186 = unuse_way == 2'h1 ? tag_1_77 : _GEN_3032; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4187 = unuse_way == 2'h1 ? tag_1_78 : _GEN_3033; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4188 = unuse_way == 2'h1 ? tag_1_79 : _GEN_3034; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4189 = unuse_way == 2'h1 ? tag_1_80 : _GEN_3035; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4190 = unuse_way == 2'h1 ? tag_1_81 : _GEN_3036; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4191 = unuse_way == 2'h1 ? tag_1_82 : _GEN_3037; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4192 = unuse_way == 2'h1 ? tag_1_83 : _GEN_3038; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4193 = unuse_way == 2'h1 ? tag_1_84 : _GEN_3039; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4194 = unuse_way == 2'h1 ? tag_1_85 : _GEN_3040; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4195 = unuse_way == 2'h1 ? tag_1_86 : _GEN_3041; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4196 = unuse_way == 2'h1 ? tag_1_87 : _GEN_3042; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4197 = unuse_way == 2'h1 ? tag_1_88 : _GEN_3043; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4198 = unuse_way == 2'h1 ? tag_1_89 : _GEN_3044; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4199 = unuse_way == 2'h1 ? tag_1_90 : _GEN_3045; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4200 = unuse_way == 2'h1 ? tag_1_91 : _GEN_3046; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4201 = unuse_way == 2'h1 ? tag_1_92 : _GEN_3047; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4202 = unuse_way == 2'h1 ? tag_1_93 : _GEN_3048; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4203 = unuse_way == 2'h1 ? tag_1_94 : _GEN_3049; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4204 = unuse_way == 2'h1 ? tag_1_95 : _GEN_3050; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4205 = unuse_way == 2'h1 ? tag_1_96 : _GEN_3051; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4206 = unuse_way == 2'h1 ? tag_1_97 : _GEN_3052; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4207 = unuse_way == 2'h1 ? tag_1_98 : _GEN_3053; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4208 = unuse_way == 2'h1 ? tag_1_99 : _GEN_3054; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4209 = unuse_way == 2'h1 ? tag_1_100 : _GEN_3055; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4210 = unuse_way == 2'h1 ? tag_1_101 : _GEN_3056; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4211 = unuse_way == 2'h1 ? tag_1_102 : _GEN_3057; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4212 = unuse_way == 2'h1 ? tag_1_103 : _GEN_3058; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4213 = unuse_way == 2'h1 ? tag_1_104 : _GEN_3059; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4214 = unuse_way == 2'h1 ? tag_1_105 : _GEN_3060; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4215 = unuse_way == 2'h1 ? tag_1_106 : _GEN_3061; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4216 = unuse_way == 2'h1 ? tag_1_107 : _GEN_3062; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4217 = unuse_way == 2'h1 ? tag_1_108 : _GEN_3063; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4218 = unuse_way == 2'h1 ? tag_1_109 : _GEN_3064; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4219 = unuse_way == 2'h1 ? tag_1_110 : _GEN_3065; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4220 = unuse_way == 2'h1 ? tag_1_111 : _GEN_3066; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4221 = unuse_way == 2'h1 ? tag_1_112 : _GEN_3067; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4222 = unuse_way == 2'h1 ? tag_1_113 : _GEN_3068; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4223 = unuse_way == 2'h1 ? tag_1_114 : _GEN_3069; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4224 = unuse_way == 2'h1 ? tag_1_115 : _GEN_3070; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4225 = unuse_way == 2'h1 ? tag_1_116 : _GEN_3071; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4226 = unuse_way == 2'h1 ? tag_1_117 : _GEN_3072; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4227 = unuse_way == 2'h1 ? tag_1_118 : _GEN_3073; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4228 = unuse_way == 2'h1 ? tag_1_119 : _GEN_3074; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4229 = unuse_way == 2'h1 ? tag_1_120 : _GEN_3075; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4230 = unuse_way == 2'h1 ? tag_1_121 : _GEN_3076; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4231 = unuse_way == 2'h1 ? tag_1_122 : _GEN_3077; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4232 = unuse_way == 2'h1 ? tag_1_123 : _GEN_3078; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4233 = unuse_way == 2'h1 ? tag_1_124 : _GEN_3079; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4234 = unuse_way == 2'h1 ? tag_1_125 : _GEN_3080; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4235 = unuse_way == 2'h1 ? tag_1_126 : _GEN_3081; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4236 = unuse_way == 2'h1 ? tag_1_127 : _GEN_3082; // @[i_cache.scala 20:24 86:34]
  wire  _GEN_4237 = unuse_way == 2'h1 ? valid_1_0 : _GEN_3083; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4238 = unuse_way == 2'h1 ? valid_1_1 : _GEN_3084; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4239 = unuse_way == 2'h1 ? valid_1_2 : _GEN_3085; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4240 = unuse_way == 2'h1 ? valid_1_3 : _GEN_3086; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4241 = unuse_way == 2'h1 ? valid_1_4 : _GEN_3087; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4242 = unuse_way == 2'h1 ? valid_1_5 : _GEN_3088; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4243 = unuse_way == 2'h1 ? valid_1_6 : _GEN_3089; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4244 = unuse_way == 2'h1 ? valid_1_7 : _GEN_3090; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4245 = unuse_way == 2'h1 ? valid_1_8 : _GEN_3091; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4246 = unuse_way == 2'h1 ? valid_1_9 : _GEN_3092; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4247 = unuse_way == 2'h1 ? valid_1_10 : _GEN_3093; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4248 = unuse_way == 2'h1 ? valid_1_11 : _GEN_3094; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4249 = unuse_way == 2'h1 ? valid_1_12 : _GEN_3095; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4250 = unuse_way == 2'h1 ? valid_1_13 : _GEN_3096; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4251 = unuse_way == 2'h1 ? valid_1_14 : _GEN_3097; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4252 = unuse_way == 2'h1 ? valid_1_15 : _GEN_3098; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4253 = unuse_way == 2'h1 ? valid_1_16 : _GEN_3099; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4254 = unuse_way == 2'h1 ? valid_1_17 : _GEN_3100; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4255 = unuse_way == 2'h1 ? valid_1_18 : _GEN_3101; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4256 = unuse_way == 2'h1 ? valid_1_19 : _GEN_3102; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4257 = unuse_way == 2'h1 ? valid_1_20 : _GEN_3103; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4258 = unuse_way == 2'h1 ? valid_1_21 : _GEN_3104; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4259 = unuse_way == 2'h1 ? valid_1_22 : _GEN_3105; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4260 = unuse_way == 2'h1 ? valid_1_23 : _GEN_3106; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4261 = unuse_way == 2'h1 ? valid_1_24 : _GEN_3107; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4262 = unuse_way == 2'h1 ? valid_1_25 : _GEN_3108; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4263 = unuse_way == 2'h1 ? valid_1_26 : _GEN_3109; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4264 = unuse_way == 2'h1 ? valid_1_27 : _GEN_3110; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4265 = unuse_way == 2'h1 ? valid_1_28 : _GEN_3111; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4266 = unuse_way == 2'h1 ? valid_1_29 : _GEN_3112; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4267 = unuse_way == 2'h1 ? valid_1_30 : _GEN_3113; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4268 = unuse_way == 2'h1 ? valid_1_31 : _GEN_3114; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4269 = unuse_way == 2'h1 ? valid_1_32 : _GEN_3115; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4270 = unuse_way == 2'h1 ? valid_1_33 : _GEN_3116; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4271 = unuse_way == 2'h1 ? valid_1_34 : _GEN_3117; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4272 = unuse_way == 2'h1 ? valid_1_35 : _GEN_3118; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4273 = unuse_way == 2'h1 ? valid_1_36 : _GEN_3119; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4274 = unuse_way == 2'h1 ? valid_1_37 : _GEN_3120; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4275 = unuse_way == 2'h1 ? valid_1_38 : _GEN_3121; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4276 = unuse_way == 2'h1 ? valid_1_39 : _GEN_3122; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4277 = unuse_way == 2'h1 ? valid_1_40 : _GEN_3123; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4278 = unuse_way == 2'h1 ? valid_1_41 : _GEN_3124; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4279 = unuse_way == 2'h1 ? valid_1_42 : _GEN_3125; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4280 = unuse_way == 2'h1 ? valid_1_43 : _GEN_3126; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4281 = unuse_way == 2'h1 ? valid_1_44 : _GEN_3127; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4282 = unuse_way == 2'h1 ? valid_1_45 : _GEN_3128; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4283 = unuse_way == 2'h1 ? valid_1_46 : _GEN_3129; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4284 = unuse_way == 2'h1 ? valid_1_47 : _GEN_3130; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4285 = unuse_way == 2'h1 ? valid_1_48 : _GEN_3131; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4286 = unuse_way == 2'h1 ? valid_1_49 : _GEN_3132; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4287 = unuse_way == 2'h1 ? valid_1_50 : _GEN_3133; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4288 = unuse_way == 2'h1 ? valid_1_51 : _GEN_3134; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4289 = unuse_way == 2'h1 ? valid_1_52 : _GEN_3135; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4290 = unuse_way == 2'h1 ? valid_1_53 : _GEN_3136; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4291 = unuse_way == 2'h1 ? valid_1_54 : _GEN_3137; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4292 = unuse_way == 2'h1 ? valid_1_55 : _GEN_3138; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4293 = unuse_way == 2'h1 ? valid_1_56 : _GEN_3139; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4294 = unuse_way == 2'h1 ? valid_1_57 : _GEN_3140; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4295 = unuse_way == 2'h1 ? valid_1_58 : _GEN_3141; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4296 = unuse_way == 2'h1 ? valid_1_59 : _GEN_3142; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4297 = unuse_way == 2'h1 ? valid_1_60 : _GEN_3143; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4298 = unuse_way == 2'h1 ? valid_1_61 : _GEN_3144; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4299 = unuse_way == 2'h1 ? valid_1_62 : _GEN_3145; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4300 = unuse_way == 2'h1 ? valid_1_63 : _GEN_3146; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4301 = unuse_way == 2'h1 ? valid_1_64 : _GEN_3147; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4302 = unuse_way == 2'h1 ? valid_1_65 : _GEN_3148; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4303 = unuse_way == 2'h1 ? valid_1_66 : _GEN_3149; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4304 = unuse_way == 2'h1 ? valid_1_67 : _GEN_3150; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4305 = unuse_way == 2'h1 ? valid_1_68 : _GEN_3151; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4306 = unuse_way == 2'h1 ? valid_1_69 : _GEN_3152; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4307 = unuse_way == 2'h1 ? valid_1_70 : _GEN_3153; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4308 = unuse_way == 2'h1 ? valid_1_71 : _GEN_3154; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4309 = unuse_way == 2'h1 ? valid_1_72 : _GEN_3155; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4310 = unuse_way == 2'h1 ? valid_1_73 : _GEN_3156; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4311 = unuse_way == 2'h1 ? valid_1_74 : _GEN_3157; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4312 = unuse_way == 2'h1 ? valid_1_75 : _GEN_3158; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4313 = unuse_way == 2'h1 ? valid_1_76 : _GEN_3159; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4314 = unuse_way == 2'h1 ? valid_1_77 : _GEN_3160; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4315 = unuse_way == 2'h1 ? valid_1_78 : _GEN_3161; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4316 = unuse_way == 2'h1 ? valid_1_79 : _GEN_3162; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4317 = unuse_way == 2'h1 ? valid_1_80 : _GEN_3163; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4318 = unuse_way == 2'h1 ? valid_1_81 : _GEN_3164; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4319 = unuse_way == 2'h1 ? valid_1_82 : _GEN_3165; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4320 = unuse_way == 2'h1 ? valid_1_83 : _GEN_3166; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4321 = unuse_way == 2'h1 ? valid_1_84 : _GEN_3167; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4322 = unuse_way == 2'h1 ? valid_1_85 : _GEN_3168; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4323 = unuse_way == 2'h1 ? valid_1_86 : _GEN_3169; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4324 = unuse_way == 2'h1 ? valid_1_87 : _GEN_3170; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4325 = unuse_way == 2'h1 ? valid_1_88 : _GEN_3171; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4326 = unuse_way == 2'h1 ? valid_1_89 : _GEN_3172; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4327 = unuse_way == 2'h1 ? valid_1_90 : _GEN_3173; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4328 = unuse_way == 2'h1 ? valid_1_91 : _GEN_3174; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4329 = unuse_way == 2'h1 ? valid_1_92 : _GEN_3175; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4330 = unuse_way == 2'h1 ? valid_1_93 : _GEN_3176; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4331 = unuse_way == 2'h1 ? valid_1_94 : _GEN_3177; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4332 = unuse_way == 2'h1 ? valid_1_95 : _GEN_3178; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4333 = unuse_way == 2'h1 ? valid_1_96 : _GEN_3179; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4334 = unuse_way == 2'h1 ? valid_1_97 : _GEN_3180; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4335 = unuse_way == 2'h1 ? valid_1_98 : _GEN_3181; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4336 = unuse_way == 2'h1 ? valid_1_99 : _GEN_3182; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4337 = unuse_way == 2'h1 ? valid_1_100 : _GEN_3183; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4338 = unuse_way == 2'h1 ? valid_1_101 : _GEN_3184; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4339 = unuse_way == 2'h1 ? valid_1_102 : _GEN_3185; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4340 = unuse_way == 2'h1 ? valid_1_103 : _GEN_3186; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4341 = unuse_way == 2'h1 ? valid_1_104 : _GEN_3187; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4342 = unuse_way == 2'h1 ? valid_1_105 : _GEN_3188; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4343 = unuse_way == 2'h1 ? valid_1_106 : _GEN_3189; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4344 = unuse_way == 2'h1 ? valid_1_107 : _GEN_3190; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4345 = unuse_way == 2'h1 ? valid_1_108 : _GEN_3191; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4346 = unuse_way == 2'h1 ? valid_1_109 : _GEN_3192; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4347 = unuse_way == 2'h1 ? valid_1_110 : _GEN_3193; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4348 = unuse_way == 2'h1 ? valid_1_111 : _GEN_3194; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4349 = unuse_way == 2'h1 ? valid_1_112 : _GEN_3195; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4350 = unuse_way == 2'h1 ? valid_1_113 : _GEN_3196; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4351 = unuse_way == 2'h1 ? valid_1_114 : _GEN_3197; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4352 = unuse_way == 2'h1 ? valid_1_115 : _GEN_3198; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4353 = unuse_way == 2'h1 ? valid_1_116 : _GEN_3199; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4354 = unuse_way == 2'h1 ? valid_1_117 : _GEN_3200; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4355 = unuse_way == 2'h1 ? valid_1_118 : _GEN_3201; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4356 = unuse_way == 2'h1 ? valid_1_119 : _GEN_3202; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4357 = unuse_way == 2'h1 ? valid_1_120 : _GEN_3203; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4358 = unuse_way == 2'h1 ? valid_1_121 : _GEN_3204; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4359 = unuse_way == 2'h1 ? valid_1_122 : _GEN_3205; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4360 = unuse_way == 2'h1 ? valid_1_123 : _GEN_3206; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4361 = unuse_way == 2'h1 ? valid_1_124 : _GEN_3207; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4362 = unuse_way == 2'h1 ? valid_1_125 : _GEN_3208; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4363 = unuse_way == 2'h1 ? valid_1_126 : _GEN_3209; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4364 = unuse_way == 2'h1 ? valid_1_127 : _GEN_3210; // @[i_cache.scala 22:26 86:34]
  wire [2:0] _GEN_4365 = 3'h4 == state ? 3'h1 : state; // @[i_cache.scala 55:18 111:19 53:24]
  wire [2:0] _GEN_4366 = 3'h3 == state ? 3'h4 : _GEN_4365; // @[i_cache.scala 55:18 85:19]
  wire [63:0] _GEN_4367 = 3'h3 == state ? _GEN_3596 : ram_0_0; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4368 = 3'h3 == state ? _GEN_3597 : ram_0_1; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4369 = 3'h3 == state ? _GEN_3598 : ram_0_2; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4370 = 3'h3 == state ? _GEN_3599 : ram_0_3; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4371 = 3'h3 == state ? _GEN_3600 : ram_0_4; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4372 = 3'h3 == state ? _GEN_3601 : ram_0_5; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4373 = 3'h3 == state ? _GEN_3602 : ram_0_6; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4374 = 3'h3 == state ? _GEN_3603 : ram_0_7; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4375 = 3'h3 == state ? _GEN_3604 : ram_0_8; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4376 = 3'h3 == state ? _GEN_3605 : ram_0_9; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4377 = 3'h3 == state ? _GEN_3606 : ram_0_10; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4378 = 3'h3 == state ? _GEN_3607 : ram_0_11; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4379 = 3'h3 == state ? _GEN_3608 : ram_0_12; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4380 = 3'h3 == state ? _GEN_3609 : ram_0_13; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4381 = 3'h3 == state ? _GEN_3610 : ram_0_14; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4382 = 3'h3 == state ? _GEN_3611 : ram_0_15; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4383 = 3'h3 == state ? _GEN_3612 : ram_0_16; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4384 = 3'h3 == state ? _GEN_3613 : ram_0_17; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4385 = 3'h3 == state ? _GEN_3614 : ram_0_18; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4386 = 3'h3 == state ? _GEN_3615 : ram_0_19; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4387 = 3'h3 == state ? _GEN_3616 : ram_0_20; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4388 = 3'h3 == state ? _GEN_3617 : ram_0_21; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4389 = 3'h3 == state ? _GEN_3618 : ram_0_22; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4390 = 3'h3 == state ? _GEN_3619 : ram_0_23; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4391 = 3'h3 == state ? _GEN_3620 : ram_0_24; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4392 = 3'h3 == state ? _GEN_3621 : ram_0_25; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4393 = 3'h3 == state ? _GEN_3622 : ram_0_26; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4394 = 3'h3 == state ? _GEN_3623 : ram_0_27; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4395 = 3'h3 == state ? _GEN_3624 : ram_0_28; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4396 = 3'h3 == state ? _GEN_3625 : ram_0_29; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4397 = 3'h3 == state ? _GEN_3626 : ram_0_30; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4398 = 3'h3 == state ? _GEN_3627 : ram_0_31; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4399 = 3'h3 == state ? _GEN_3628 : ram_0_32; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4400 = 3'h3 == state ? _GEN_3629 : ram_0_33; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4401 = 3'h3 == state ? _GEN_3630 : ram_0_34; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4402 = 3'h3 == state ? _GEN_3631 : ram_0_35; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4403 = 3'h3 == state ? _GEN_3632 : ram_0_36; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4404 = 3'h3 == state ? _GEN_3633 : ram_0_37; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4405 = 3'h3 == state ? _GEN_3634 : ram_0_38; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4406 = 3'h3 == state ? _GEN_3635 : ram_0_39; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4407 = 3'h3 == state ? _GEN_3636 : ram_0_40; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4408 = 3'h3 == state ? _GEN_3637 : ram_0_41; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4409 = 3'h3 == state ? _GEN_3638 : ram_0_42; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4410 = 3'h3 == state ? _GEN_3639 : ram_0_43; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4411 = 3'h3 == state ? _GEN_3640 : ram_0_44; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4412 = 3'h3 == state ? _GEN_3641 : ram_0_45; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4413 = 3'h3 == state ? _GEN_3642 : ram_0_46; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4414 = 3'h3 == state ? _GEN_3643 : ram_0_47; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4415 = 3'h3 == state ? _GEN_3644 : ram_0_48; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4416 = 3'h3 == state ? _GEN_3645 : ram_0_49; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4417 = 3'h3 == state ? _GEN_3646 : ram_0_50; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4418 = 3'h3 == state ? _GEN_3647 : ram_0_51; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4419 = 3'h3 == state ? _GEN_3648 : ram_0_52; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4420 = 3'h3 == state ? _GEN_3649 : ram_0_53; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4421 = 3'h3 == state ? _GEN_3650 : ram_0_54; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4422 = 3'h3 == state ? _GEN_3651 : ram_0_55; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4423 = 3'h3 == state ? _GEN_3652 : ram_0_56; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4424 = 3'h3 == state ? _GEN_3653 : ram_0_57; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4425 = 3'h3 == state ? _GEN_3654 : ram_0_58; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4426 = 3'h3 == state ? _GEN_3655 : ram_0_59; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4427 = 3'h3 == state ? _GEN_3656 : ram_0_60; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4428 = 3'h3 == state ? _GEN_3657 : ram_0_61; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4429 = 3'h3 == state ? _GEN_3658 : ram_0_62; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4430 = 3'h3 == state ? _GEN_3659 : ram_0_63; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4431 = 3'h3 == state ? _GEN_3660 : ram_0_64; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4432 = 3'h3 == state ? _GEN_3661 : ram_0_65; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4433 = 3'h3 == state ? _GEN_3662 : ram_0_66; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4434 = 3'h3 == state ? _GEN_3663 : ram_0_67; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4435 = 3'h3 == state ? _GEN_3664 : ram_0_68; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4436 = 3'h3 == state ? _GEN_3665 : ram_0_69; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4437 = 3'h3 == state ? _GEN_3666 : ram_0_70; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4438 = 3'h3 == state ? _GEN_3667 : ram_0_71; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4439 = 3'h3 == state ? _GEN_3668 : ram_0_72; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4440 = 3'h3 == state ? _GEN_3669 : ram_0_73; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4441 = 3'h3 == state ? _GEN_3670 : ram_0_74; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4442 = 3'h3 == state ? _GEN_3671 : ram_0_75; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4443 = 3'h3 == state ? _GEN_3672 : ram_0_76; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4444 = 3'h3 == state ? _GEN_3673 : ram_0_77; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4445 = 3'h3 == state ? _GEN_3674 : ram_0_78; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4446 = 3'h3 == state ? _GEN_3675 : ram_0_79; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4447 = 3'h3 == state ? _GEN_3676 : ram_0_80; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4448 = 3'h3 == state ? _GEN_3677 : ram_0_81; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4449 = 3'h3 == state ? _GEN_3678 : ram_0_82; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4450 = 3'h3 == state ? _GEN_3679 : ram_0_83; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4451 = 3'h3 == state ? _GEN_3680 : ram_0_84; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4452 = 3'h3 == state ? _GEN_3681 : ram_0_85; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4453 = 3'h3 == state ? _GEN_3682 : ram_0_86; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4454 = 3'h3 == state ? _GEN_3683 : ram_0_87; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4455 = 3'h3 == state ? _GEN_3684 : ram_0_88; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4456 = 3'h3 == state ? _GEN_3685 : ram_0_89; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4457 = 3'h3 == state ? _GEN_3686 : ram_0_90; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4458 = 3'h3 == state ? _GEN_3687 : ram_0_91; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4459 = 3'h3 == state ? _GEN_3688 : ram_0_92; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4460 = 3'h3 == state ? _GEN_3689 : ram_0_93; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4461 = 3'h3 == state ? _GEN_3690 : ram_0_94; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4462 = 3'h3 == state ? _GEN_3691 : ram_0_95; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4463 = 3'h3 == state ? _GEN_3692 : ram_0_96; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4464 = 3'h3 == state ? _GEN_3693 : ram_0_97; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4465 = 3'h3 == state ? _GEN_3694 : ram_0_98; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4466 = 3'h3 == state ? _GEN_3695 : ram_0_99; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4467 = 3'h3 == state ? _GEN_3696 : ram_0_100; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4468 = 3'h3 == state ? _GEN_3697 : ram_0_101; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4469 = 3'h3 == state ? _GEN_3698 : ram_0_102; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4470 = 3'h3 == state ? _GEN_3699 : ram_0_103; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4471 = 3'h3 == state ? _GEN_3700 : ram_0_104; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4472 = 3'h3 == state ? _GEN_3701 : ram_0_105; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4473 = 3'h3 == state ? _GEN_3702 : ram_0_106; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4474 = 3'h3 == state ? _GEN_3703 : ram_0_107; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4475 = 3'h3 == state ? _GEN_3704 : ram_0_108; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4476 = 3'h3 == state ? _GEN_3705 : ram_0_109; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4477 = 3'h3 == state ? _GEN_3706 : ram_0_110; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4478 = 3'h3 == state ? _GEN_3707 : ram_0_111; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4479 = 3'h3 == state ? _GEN_3708 : ram_0_112; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4480 = 3'h3 == state ? _GEN_3709 : ram_0_113; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4481 = 3'h3 == state ? _GEN_3710 : ram_0_114; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4482 = 3'h3 == state ? _GEN_3711 : ram_0_115; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4483 = 3'h3 == state ? _GEN_3712 : ram_0_116; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4484 = 3'h3 == state ? _GEN_3713 : ram_0_117; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4485 = 3'h3 == state ? _GEN_3714 : ram_0_118; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4486 = 3'h3 == state ? _GEN_3715 : ram_0_119; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4487 = 3'h3 == state ? _GEN_3716 : ram_0_120; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4488 = 3'h3 == state ? _GEN_3717 : ram_0_121; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4489 = 3'h3 == state ? _GEN_3718 : ram_0_122; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4490 = 3'h3 == state ? _GEN_3719 : ram_0_123; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4491 = 3'h3 == state ? _GEN_3720 : ram_0_124; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4492 = 3'h3 == state ? _GEN_3721 : ram_0_125; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4493 = 3'h3 == state ? _GEN_3722 : ram_0_126; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4494 = 3'h3 == state ? _GEN_3723 : ram_0_127; // @[i_cache.scala 55:18 17:24]
  wire [31:0] _GEN_4495 = 3'h3 == state ? _GEN_3724 : tag_0_0; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4496 = 3'h3 == state ? _GEN_3725 : tag_0_1; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4497 = 3'h3 == state ? _GEN_3726 : tag_0_2; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4498 = 3'h3 == state ? _GEN_3727 : tag_0_3; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4499 = 3'h3 == state ? _GEN_3728 : tag_0_4; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4500 = 3'h3 == state ? _GEN_3729 : tag_0_5; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4501 = 3'h3 == state ? _GEN_3730 : tag_0_6; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4502 = 3'h3 == state ? _GEN_3731 : tag_0_7; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4503 = 3'h3 == state ? _GEN_3732 : tag_0_8; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4504 = 3'h3 == state ? _GEN_3733 : tag_0_9; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4505 = 3'h3 == state ? _GEN_3734 : tag_0_10; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4506 = 3'h3 == state ? _GEN_3735 : tag_0_11; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4507 = 3'h3 == state ? _GEN_3736 : tag_0_12; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4508 = 3'h3 == state ? _GEN_3737 : tag_0_13; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4509 = 3'h3 == state ? _GEN_3738 : tag_0_14; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4510 = 3'h3 == state ? _GEN_3739 : tag_0_15; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4511 = 3'h3 == state ? _GEN_3740 : tag_0_16; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4512 = 3'h3 == state ? _GEN_3741 : tag_0_17; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4513 = 3'h3 == state ? _GEN_3742 : tag_0_18; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4514 = 3'h3 == state ? _GEN_3743 : tag_0_19; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4515 = 3'h3 == state ? _GEN_3744 : tag_0_20; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4516 = 3'h3 == state ? _GEN_3745 : tag_0_21; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4517 = 3'h3 == state ? _GEN_3746 : tag_0_22; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4518 = 3'h3 == state ? _GEN_3747 : tag_0_23; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4519 = 3'h3 == state ? _GEN_3748 : tag_0_24; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4520 = 3'h3 == state ? _GEN_3749 : tag_0_25; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4521 = 3'h3 == state ? _GEN_3750 : tag_0_26; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4522 = 3'h3 == state ? _GEN_3751 : tag_0_27; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4523 = 3'h3 == state ? _GEN_3752 : tag_0_28; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4524 = 3'h3 == state ? _GEN_3753 : tag_0_29; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4525 = 3'h3 == state ? _GEN_3754 : tag_0_30; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4526 = 3'h3 == state ? _GEN_3755 : tag_0_31; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4527 = 3'h3 == state ? _GEN_3756 : tag_0_32; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4528 = 3'h3 == state ? _GEN_3757 : tag_0_33; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4529 = 3'h3 == state ? _GEN_3758 : tag_0_34; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4530 = 3'h3 == state ? _GEN_3759 : tag_0_35; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4531 = 3'h3 == state ? _GEN_3760 : tag_0_36; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4532 = 3'h3 == state ? _GEN_3761 : tag_0_37; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4533 = 3'h3 == state ? _GEN_3762 : tag_0_38; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4534 = 3'h3 == state ? _GEN_3763 : tag_0_39; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4535 = 3'h3 == state ? _GEN_3764 : tag_0_40; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4536 = 3'h3 == state ? _GEN_3765 : tag_0_41; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4537 = 3'h3 == state ? _GEN_3766 : tag_0_42; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4538 = 3'h3 == state ? _GEN_3767 : tag_0_43; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4539 = 3'h3 == state ? _GEN_3768 : tag_0_44; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4540 = 3'h3 == state ? _GEN_3769 : tag_0_45; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4541 = 3'h3 == state ? _GEN_3770 : tag_0_46; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4542 = 3'h3 == state ? _GEN_3771 : tag_0_47; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4543 = 3'h3 == state ? _GEN_3772 : tag_0_48; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4544 = 3'h3 == state ? _GEN_3773 : tag_0_49; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4545 = 3'h3 == state ? _GEN_3774 : tag_0_50; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4546 = 3'h3 == state ? _GEN_3775 : tag_0_51; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4547 = 3'h3 == state ? _GEN_3776 : tag_0_52; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4548 = 3'h3 == state ? _GEN_3777 : tag_0_53; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4549 = 3'h3 == state ? _GEN_3778 : tag_0_54; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4550 = 3'h3 == state ? _GEN_3779 : tag_0_55; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4551 = 3'h3 == state ? _GEN_3780 : tag_0_56; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4552 = 3'h3 == state ? _GEN_3781 : tag_0_57; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4553 = 3'h3 == state ? _GEN_3782 : tag_0_58; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4554 = 3'h3 == state ? _GEN_3783 : tag_0_59; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4555 = 3'h3 == state ? _GEN_3784 : tag_0_60; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4556 = 3'h3 == state ? _GEN_3785 : tag_0_61; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4557 = 3'h3 == state ? _GEN_3786 : tag_0_62; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4558 = 3'h3 == state ? _GEN_3787 : tag_0_63; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4559 = 3'h3 == state ? _GEN_3788 : tag_0_64; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4560 = 3'h3 == state ? _GEN_3789 : tag_0_65; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4561 = 3'h3 == state ? _GEN_3790 : tag_0_66; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4562 = 3'h3 == state ? _GEN_3791 : tag_0_67; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4563 = 3'h3 == state ? _GEN_3792 : tag_0_68; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4564 = 3'h3 == state ? _GEN_3793 : tag_0_69; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4565 = 3'h3 == state ? _GEN_3794 : tag_0_70; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4566 = 3'h3 == state ? _GEN_3795 : tag_0_71; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4567 = 3'h3 == state ? _GEN_3796 : tag_0_72; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4568 = 3'h3 == state ? _GEN_3797 : tag_0_73; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4569 = 3'h3 == state ? _GEN_3798 : tag_0_74; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4570 = 3'h3 == state ? _GEN_3799 : tag_0_75; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4571 = 3'h3 == state ? _GEN_3800 : tag_0_76; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4572 = 3'h3 == state ? _GEN_3801 : tag_0_77; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4573 = 3'h3 == state ? _GEN_3802 : tag_0_78; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4574 = 3'h3 == state ? _GEN_3803 : tag_0_79; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4575 = 3'h3 == state ? _GEN_3804 : tag_0_80; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4576 = 3'h3 == state ? _GEN_3805 : tag_0_81; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4577 = 3'h3 == state ? _GEN_3806 : tag_0_82; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4578 = 3'h3 == state ? _GEN_3807 : tag_0_83; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4579 = 3'h3 == state ? _GEN_3808 : tag_0_84; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4580 = 3'h3 == state ? _GEN_3809 : tag_0_85; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4581 = 3'h3 == state ? _GEN_3810 : tag_0_86; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4582 = 3'h3 == state ? _GEN_3811 : tag_0_87; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4583 = 3'h3 == state ? _GEN_3812 : tag_0_88; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4584 = 3'h3 == state ? _GEN_3813 : tag_0_89; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4585 = 3'h3 == state ? _GEN_3814 : tag_0_90; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4586 = 3'h3 == state ? _GEN_3815 : tag_0_91; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4587 = 3'h3 == state ? _GEN_3816 : tag_0_92; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4588 = 3'h3 == state ? _GEN_3817 : tag_0_93; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4589 = 3'h3 == state ? _GEN_3818 : tag_0_94; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4590 = 3'h3 == state ? _GEN_3819 : tag_0_95; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4591 = 3'h3 == state ? _GEN_3820 : tag_0_96; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4592 = 3'h3 == state ? _GEN_3821 : tag_0_97; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4593 = 3'h3 == state ? _GEN_3822 : tag_0_98; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4594 = 3'h3 == state ? _GEN_3823 : tag_0_99; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4595 = 3'h3 == state ? _GEN_3824 : tag_0_100; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4596 = 3'h3 == state ? _GEN_3825 : tag_0_101; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4597 = 3'h3 == state ? _GEN_3826 : tag_0_102; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4598 = 3'h3 == state ? _GEN_3827 : tag_0_103; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4599 = 3'h3 == state ? _GEN_3828 : tag_0_104; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4600 = 3'h3 == state ? _GEN_3829 : tag_0_105; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4601 = 3'h3 == state ? _GEN_3830 : tag_0_106; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4602 = 3'h3 == state ? _GEN_3831 : tag_0_107; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4603 = 3'h3 == state ? _GEN_3832 : tag_0_108; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4604 = 3'h3 == state ? _GEN_3833 : tag_0_109; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4605 = 3'h3 == state ? _GEN_3834 : tag_0_110; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4606 = 3'h3 == state ? _GEN_3835 : tag_0_111; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4607 = 3'h3 == state ? _GEN_3836 : tag_0_112; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4608 = 3'h3 == state ? _GEN_3837 : tag_0_113; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4609 = 3'h3 == state ? _GEN_3838 : tag_0_114; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4610 = 3'h3 == state ? _GEN_3839 : tag_0_115; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4611 = 3'h3 == state ? _GEN_3840 : tag_0_116; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4612 = 3'h3 == state ? _GEN_3841 : tag_0_117; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4613 = 3'h3 == state ? _GEN_3842 : tag_0_118; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4614 = 3'h3 == state ? _GEN_3843 : tag_0_119; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4615 = 3'h3 == state ? _GEN_3844 : tag_0_120; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4616 = 3'h3 == state ? _GEN_3845 : tag_0_121; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4617 = 3'h3 == state ? _GEN_3846 : tag_0_122; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4618 = 3'h3 == state ? _GEN_3847 : tag_0_123; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4619 = 3'h3 == state ? _GEN_3848 : tag_0_124; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4620 = 3'h3 == state ? _GEN_3849 : tag_0_125; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4621 = 3'h3 == state ? _GEN_3850 : tag_0_126; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4622 = 3'h3 == state ? _GEN_3851 : tag_0_127; // @[i_cache.scala 55:18 19:24]
  wire  _GEN_4623 = 3'h3 == state ? _GEN_3852 : valid_0_0; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4624 = 3'h3 == state ? _GEN_3853 : valid_0_1; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4625 = 3'h3 == state ? _GEN_3854 : valid_0_2; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4626 = 3'h3 == state ? _GEN_3855 : valid_0_3; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4627 = 3'h3 == state ? _GEN_3856 : valid_0_4; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4628 = 3'h3 == state ? _GEN_3857 : valid_0_5; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4629 = 3'h3 == state ? _GEN_3858 : valid_0_6; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4630 = 3'h3 == state ? _GEN_3859 : valid_0_7; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4631 = 3'h3 == state ? _GEN_3860 : valid_0_8; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4632 = 3'h3 == state ? _GEN_3861 : valid_0_9; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4633 = 3'h3 == state ? _GEN_3862 : valid_0_10; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4634 = 3'h3 == state ? _GEN_3863 : valid_0_11; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4635 = 3'h3 == state ? _GEN_3864 : valid_0_12; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4636 = 3'h3 == state ? _GEN_3865 : valid_0_13; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4637 = 3'h3 == state ? _GEN_3866 : valid_0_14; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4638 = 3'h3 == state ? _GEN_3867 : valid_0_15; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4639 = 3'h3 == state ? _GEN_3868 : valid_0_16; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4640 = 3'h3 == state ? _GEN_3869 : valid_0_17; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4641 = 3'h3 == state ? _GEN_3870 : valid_0_18; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4642 = 3'h3 == state ? _GEN_3871 : valid_0_19; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4643 = 3'h3 == state ? _GEN_3872 : valid_0_20; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4644 = 3'h3 == state ? _GEN_3873 : valid_0_21; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4645 = 3'h3 == state ? _GEN_3874 : valid_0_22; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4646 = 3'h3 == state ? _GEN_3875 : valid_0_23; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4647 = 3'h3 == state ? _GEN_3876 : valid_0_24; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4648 = 3'h3 == state ? _GEN_3877 : valid_0_25; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4649 = 3'h3 == state ? _GEN_3878 : valid_0_26; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4650 = 3'h3 == state ? _GEN_3879 : valid_0_27; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4651 = 3'h3 == state ? _GEN_3880 : valid_0_28; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4652 = 3'h3 == state ? _GEN_3881 : valid_0_29; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4653 = 3'h3 == state ? _GEN_3882 : valid_0_30; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4654 = 3'h3 == state ? _GEN_3883 : valid_0_31; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4655 = 3'h3 == state ? _GEN_3884 : valid_0_32; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4656 = 3'h3 == state ? _GEN_3885 : valid_0_33; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4657 = 3'h3 == state ? _GEN_3886 : valid_0_34; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4658 = 3'h3 == state ? _GEN_3887 : valid_0_35; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4659 = 3'h3 == state ? _GEN_3888 : valid_0_36; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4660 = 3'h3 == state ? _GEN_3889 : valid_0_37; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4661 = 3'h3 == state ? _GEN_3890 : valid_0_38; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4662 = 3'h3 == state ? _GEN_3891 : valid_0_39; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4663 = 3'h3 == state ? _GEN_3892 : valid_0_40; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4664 = 3'h3 == state ? _GEN_3893 : valid_0_41; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4665 = 3'h3 == state ? _GEN_3894 : valid_0_42; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4666 = 3'h3 == state ? _GEN_3895 : valid_0_43; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4667 = 3'h3 == state ? _GEN_3896 : valid_0_44; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4668 = 3'h3 == state ? _GEN_3897 : valid_0_45; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4669 = 3'h3 == state ? _GEN_3898 : valid_0_46; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4670 = 3'h3 == state ? _GEN_3899 : valid_0_47; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4671 = 3'h3 == state ? _GEN_3900 : valid_0_48; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4672 = 3'h3 == state ? _GEN_3901 : valid_0_49; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4673 = 3'h3 == state ? _GEN_3902 : valid_0_50; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4674 = 3'h3 == state ? _GEN_3903 : valid_0_51; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4675 = 3'h3 == state ? _GEN_3904 : valid_0_52; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4676 = 3'h3 == state ? _GEN_3905 : valid_0_53; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4677 = 3'h3 == state ? _GEN_3906 : valid_0_54; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4678 = 3'h3 == state ? _GEN_3907 : valid_0_55; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4679 = 3'h3 == state ? _GEN_3908 : valid_0_56; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4680 = 3'h3 == state ? _GEN_3909 : valid_0_57; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4681 = 3'h3 == state ? _GEN_3910 : valid_0_58; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4682 = 3'h3 == state ? _GEN_3911 : valid_0_59; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4683 = 3'h3 == state ? _GEN_3912 : valid_0_60; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4684 = 3'h3 == state ? _GEN_3913 : valid_0_61; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4685 = 3'h3 == state ? _GEN_3914 : valid_0_62; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4686 = 3'h3 == state ? _GEN_3915 : valid_0_63; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4687 = 3'h3 == state ? _GEN_3916 : valid_0_64; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4688 = 3'h3 == state ? _GEN_3917 : valid_0_65; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4689 = 3'h3 == state ? _GEN_3918 : valid_0_66; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4690 = 3'h3 == state ? _GEN_3919 : valid_0_67; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4691 = 3'h3 == state ? _GEN_3920 : valid_0_68; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4692 = 3'h3 == state ? _GEN_3921 : valid_0_69; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4693 = 3'h3 == state ? _GEN_3922 : valid_0_70; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4694 = 3'h3 == state ? _GEN_3923 : valid_0_71; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4695 = 3'h3 == state ? _GEN_3924 : valid_0_72; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4696 = 3'h3 == state ? _GEN_3925 : valid_0_73; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4697 = 3'h3 == state ? _GEN_3926 : valid_0_74; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4698 = 3'h3 == state ? _GEN_3927 : valid_0_75; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4699 = 3'h3 == state ? _GEN_3928 : valid_0_76; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4700 = 3'h3 == state ? _GEN_3929 : valid_0_77; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4701 = 3'h3 == state ? _GEN_3930 : valid_0_78; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4702 = 3'h3 == state ? _GEN_3931 : valid_0_79; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4703 = 3'h3 == state ? _GEN_3932 : valid_0_80; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4704 = 3'h3 == state ? _GEN_3933 : valid_0_81; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4705 = 3'h3 == state ? _GEN_3934 : valid_0_82; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4706 = 3'h3 == state ? _GEN_3935 : valid_0_83; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4707 = 3'h3 == state ? _GEN_3936 : valid_0_84; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4708 = 3'h3 == state ? _GEN_3937 : valid_0_85; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4709 = 3'h3 == state ? _GEN_3938 : valid_0_86; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4710 = 3'h3 == state ? _GEN_3939 : valid_0_87; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4711 = 3'h3 == state ? _GEN_3940 : valid_0_88; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4712 = 3'h3 == state ? _GEN_3941 : valid_0_89; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4713 = 3'h3 == state ? _GEN_3942 : valid_0_90; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4714 = 3'h3 == state ? _GEN_3943 : valid_0_91; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4715 = 3'h3 == state ? _GEN_3944 : valid_0_92; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4716 = 3'h3 == state ? _GEN_3945 : valid_0_93; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4717 = 3'h3 == state ? _GEN_3946 : valid_0_94; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4718 = 3'h3 == state ? _GEN_3947 : valid_0_95; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4719 = 3'h3 == state ? _GEN_3948 : valid_0_96; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4720 = 3'h3 == state ? _GEN_3949 : valid_0_97; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4721 = 3'h3 == state ? _GEN_3950 : valid_0_98; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4722 = 3'h3 == state ? _GEN_3951 : valid_0_99; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4723 = 3'h3 == state ? _GEN_3952 : valid_0_100; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4724 = 3'h3 == state ? _GEN_3953 : valid_0_101; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4725 = 3'h3 == state ? _GEN_3954 : valid_0_102; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4726 = 3'h3 == state ? _GEN_3955 : valid_0_103; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4727 = 3'h3 == state ? _GEN_3956 : valid_0_104; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4728 = 3'h3 == state ? _GEN_3957 : valid_0_105; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4729 = 3'h3 == state ? _GEN_3958 : valid_0_106; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4730 = 3'h3 == state ? _GEN_3959 : valid_0_107; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4731 = 3'h3 == state ? _GEN_3960 : valid_0_108; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4732 = 3'h3 == state ? _GEN_3961 : valid_0_109; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4733 = 3'h3 == state ? _GEN_3962 : valid_0_110; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4734 = 3'h3 == state ? _GEN_3963 : valid_0_111; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4735 = 3'h3 == state ? _GEN_3964 : valid_0_112; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4736 = 3'h3 == state ? _GEN_3965 : valid_0_113; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4737 = 3'h3 == state ? _GEN_3966 : valid_0_114; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4738 = 3'h3 == state ? _GEN_3967 : valid_0_115; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4739 = 3'h3 == state ? _GEN_3968 : valid_0_116; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4740 = 3'h3 == state ? _GEN_3969 : valid_0_117; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4741 = 3'h3 == state ? _GEN_3970 : valid_0_118; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4742 = 3'h3 == state ? _GEN_3971 : valid_0_119; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4743 = 3'h3 == state ? _GEN_3972 : valid_0_120; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4744 = 3'h3 == state ? _GEN_3973 : valid_0_121; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4745 = 3'h3 == state ? _GEN_3974 : valid_0_122; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4746 = 3'h3 == state ? _GEN_3975 : valid_0_123; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4747 = 3'h3 == state ? _GEN_3976 : valid_0_124; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4748 = 3'h3 == state ? _GEN_3977 : valid_0_125; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4749 = 3'h3 == state ? _GEN_3978 : valid_0_126; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4750 = 3'h3 == state ? _GEN_3979 : valid_0_127; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4751 = 3'h3 == state ? _GEN_3980 : quene; // @[i_cache.scala 55:18 28:24]
  wire [63:0] _GEN_4752 = 3'h3 == state ? _GEN_3981 : ram_1_0; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4753 = 3'h3 == state ? _GEN_3982 : ram_1_1; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4754 = 3'h3 == state ? _GEN_3983 : ram_1_2; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4755 = 3'h3 == state ? _GEN_3984 : ram_1_3; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4756 = 3'h3 == state ? _GEN_3985 : ram_1_4; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4757 = 3'h3 == state ? _GEN_3986 : ram_1_5; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4758 = 3'h3 == state ? _GEN_3987 : ram_1_6; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4759 = 3'h3 == state ? _GEN_3988 : ram_1_7; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4760 = 3'h3 == state ? _GEN_3989 : ram_1_8; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4761 = 3'h3 == state ? _GEN_3990 : ram_1_9; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4762 = 3'h3 == state ? _GEN_3991 : ram_1_10; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4763 = 3'h3 == state ? _GEN_3992 : ram_1_11; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4764 = 3'h3 == state ? _GEN_3993 : ram_1_12; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4765 = 3'h3 == state ? _GEN_3994 : ram_1_13; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4766 = 3'h3 == state ? _GEN_3995 : ram_1_14; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4767 = 3'h3 == state ? _GEN_3996 : ram_1_15; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4768 = 3'h3 == state ? _GEN_3997 : ram_1_16; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4769 = 3'h3 == state ? _GEN_3998 : ram_1_17; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4770 = 3'h3 == state ? _GEN_3999 : ram_1_18; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4771 = 3'h3 == state ? _GEN_4000 : ram_1_19; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4772 = 3'h3 == state ? _GEN_4001 : ram_1_20; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4773 = 3'h3 == state ? _GEN_4002 : ram_1_21; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4774 = 3'h3 == state ? _GEN_4003 : ram_1_22; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4775 = 3'h3 == state ? _GEN_4004 : ram_1_23; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4776 = 3'h3 == state ? _GEN_4005 : ram_1_24; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4777 = 3'h3 == state ? _GEN_4006 : ram_1_25; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4778 = 3'h3 == state ? _GEN_4007 : ram_1_26; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4779 = 3'h3 == state ? _GEN_4008 : ram_1_27; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4780 = 3'h3 == state ? _GEN_4009 : ram_1_28; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4781 = 3'h3 == state ? _GEN_4010 : ram_1_29; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4782 = 3'h3 == state ? _GEN_4011 : ram_1_30; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4783 = 3'h3 == state ? _GEN_4012 : ram_1_31; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4784 = 3'h3 == state ? _GEN_4013 : ram_1_32; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4785 = 3'h3 == state ? _GEN_4014 : ram_1_33; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4786 = 3'h3 == state ? _GEN_4015 : ram_1_34; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4787 = 3'h3 == state ? _GEN_4016 : ram_1_35; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4788 = 3'h3 == state ? _GEN_4017 : ram_1_36; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4789 = 3'h3 == state ? _GEN_4018 : ram_1_37; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4790 = 3'h3 == state ? _GEN_4019 : ram_1_38; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4791 = 3'h3 == state ? _GEN_4020 : ram_1_39; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4792 = 3'h3 == state ? _GEN_4021 : ram_1_40; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4793 = 3'h3 == state ? _GEN_4022 : ram_1_41; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4794 = 3'h3 == state ? _GEN_4023 : ram_1_42; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4795 = 3'h3 == state ? _GEN_4024 : ram_1_43; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4796 = 3'h3 == state ? _GEN_4025 : ram_1_44; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4797 = 3'h3 == state ? _GEN_4026 : ram_1_45; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4798 = 3'h3 == state ? _GEN_4027 : ram_1_46; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4799 = 3'h3 == state ? _GEN_4028 : ram_1_47; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4800 = 3'h3 == state ? _GEN_4029 : ram_1_48; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4801 = 3'h3 == state ? _GEN_4030 : ram_1_49; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4802 = 3'h3 == state ? _GEN_4031 : ram_1_50; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4803 = 3'h3 == state ? _GEN_4032 : ram_1_51; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4804 = 3'h3 == state ? _GEN_4033 : ram_1_52; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4805 = 3'h3 == state ? _GEN_4034 : ram_1_53; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4806 = 3'h3 == state ? _GEN_4035 : ram_1_54; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4807 = 3'h3 == state ? _GEN_4036 : ram_1_55; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4808 = 3'h3 == state ? _GEN_4037 : ram_1_56; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4809 = 3'h3 == state ? _GEN_4038 : ram_1_57; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4810 = 3'h3 == state ? _GEN_4039 : ram_1_58; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4811 = 3'h3 == state ? _GEN_4040 : ram_1_59; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4812 = 3'h3 == state ? _GEN_4041 : ram_1_60; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4813 = 3'h3 == state ? _GEN_4042 : ram_1_61; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4814 = 3'h3 == state ? _GEN_4043 : ram_1_62; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4815 = 3'h3 == state ? _GEN_4044 : ram_1_63; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4816 = 3'h3 == state ? _GEN_4045 : ram_1_64; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4817 = 3'h3 == state ? _GEN_4046 : ram_1_65; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4818 = 3'h3 == state ? _GEN_4047 : ram_1_66; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4819 = 3'h3 == state ? _GEN_4048 : ram_1_67; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4820 = 3'h3 == state ? _GEN_4049 : ram_1_68; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4821 = 3'h3 == state ? _GEN_4050 : ram_1_69; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4822 = 3'h3 == state ? _GEN_4051 : ram_1_70; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4823 = 3'h3 == state ? _GEN_4052 : ram_1_71; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4824 = 3'h3 == state ? _GEN_4053 : ram_1_72; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4825 = 3'h3 == state ? _GEN_4054 : ram_1_73; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4826 = 3'h3 == state ? _GEN_4055 : ram_1_74; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4827 = 3'h3 == state ? _GEN_4056 : ram_1_75; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4828 = 3'h3 == state ? _GEN_4057 : ram_1_76; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4829 = 3'h3 == state ? _GEN_4058 : ram_1_77; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4830 = 3'h3 == state ? _GEN_4059 : ram_1_78; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4831 = 3'h3 == state ? _GEN_4060 : ram_1_79; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4832 = 3'h3 == state ? _GEN_4061 : ram_1_80; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4833 = 3'h3 == state ? _GEN_4062 : ram_1_81; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4834 = 3'h3 == state ? _GEN_4063 : ram_1_82; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4835 = 3'h3 == state ? _GEN_4064 : ram_1_83; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4836 = 3'h3 == state ? _GEN_4065 : ram_1_84; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4837 = 3'h3 == state ? _GEN_4066 : ram_1_85; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4838 = 3'h3 == state ? _GEN_4067 : ram_1_86; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4839 = 3'h3 == state ? _GEN_4068 : ram_1_87; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4840 = 3'h3 == state ? _GEN_4069 : ram_1_88; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4841 = 3'h3 == state ? _GEN_4070 : ram_1_89; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4842 = 3'h3 == state ? _GEN_4071 : ram_1_90; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4843 = 3'h3 == state ? _GEN_4072 : ram_1_91; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4844 = 3'h3 == state ? _GEN_4073 : ram_1_92; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4845 = 3'h3 == state ? _GEN_4074 : ram_1_93; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4846 = 3'h3 == state ? _GEN_4075 : ram_1_94; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4847 = 3'h3 == state ? _GEN_4076 : ram_1_95; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4848 = 3'h3 == state ? _GEN_4077 : ram_1_96; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4849 = 3'h3 == state ? _GEN_4078 : ram_1_97; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4850 = 3'h3 == state ? _GEN_4079 : ram_1_98; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4851 = 3'h3 == state ? _GEN_4080 : ram_1_99; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4852 = 3'h3 == state ? _GEN_4081 : ram_1_100; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4853 = 3'h3 == state ? _GEN_4082 : ram_1_101; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4854 = 3'h3 == state ? _GEN_4083 : ram_1_102; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4855 = 3'h3 == state ? _GEN_4084 : ram_1_103; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4856 = 3'h3 == state ? _GEN_4085 : ram_1_104; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4857 = 3'h3 == state ? _GEN_4086 : ram_1_105; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4858 = 3'h3 == state ? _GEN_4087 : ram_1_106; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4859 = 3'h3 == state ? _GEN_4088 : ram_1_107; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4860 = 3'h3 == state ? _GEN_4089 : ram_1_108; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4861 = 3'h3 == state ? _GEN_4090 : ram_1_109; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4862 = 3'h3 == state ? _GEN_4091 : ram_1_110; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4863 = 3'h3 == state ? _GEN_4092 : ram_1_111; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4864 = 3'h3 == state ? _GEN_4093 : ram_1_112; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4865 = 3'h3 == state ? _GEN_4094 : ram_1_113; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4866 = 3'h3 == state ? _GEN_4095 : ram_1_114; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4867 = 3'h3 == state ? _GEN_4096 : ram_1_115; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4868 = 3'h3 == state ? _GEN_4097 : ram_1_116; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4869 = 3'h3 == state ? _GEN_4098 : ram_1_117; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4870 = 3'h3 == state ? _GEN_4099 : ram_1_118; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4871 = 3'h3 == state ? _GEN_4100 : ram_1_119; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4872 = 3'h3 == state ? _GEN_4101 : ram_1_120; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4873 = 3'h3 == state ? _GEN_4102 : ram_1_121; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4874 = 3'h3 == state ? _GEN_4103 : ram_1_122; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4875 = 3'h3 == state ? _GEN_4104 : ram_1_123; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4876 = 3'h3 == state ? _GEN_4105 : ram_1_124; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4877 = 3'h3 == state ? _GEN_4106 : ram_1_125; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4878 = 3'h3 == state ? _GEN_4107 : ram_1_126; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4879 = 3'h3 == state ? _GEN_4108 : ram_1_127; // @[i_cache.scala 55:18 18:24]
  wire [31:0] _GEN_4880 = 3'h3 == state ? _GEN_4109 : tag_1_0; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4881 = 3'h3 == state ? _GEN_4110 : tag_1_1; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4882 = 3'h3 == state ? _GEN_4111 : tag_1_2; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4883 = 3'h3 == state ? _GEN_4112 : tag_1_3; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4884 = 3'h3 == state ? _GEN_4113 : tag_1_4; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4885 = 3'h3 == state ? _GEN_4114 : tag_1_5; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4886 = 3'h3 == state ? _GEN_4115 : tag_1_6; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4887 = 3'h3 == state ? _GEN_4116 : tag_1_7; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4888 = 3'h3 == state ? _GEN_4117 : tag_1_8; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4889 = 3'h3 == state ? _GEN_4118 : tag_1_9; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4890 = 3'h3 == state ? _GEN_4119 : tag_1_10; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4891 = 3'h3 == state ? _GEN_4120 : tag_1_11; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4892 = 3'h3 == state ? _GEN_4121 : tag_1_12; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4893 = 3'h3 == state ? _GEN_4122 : tag_1_13; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4894 = 3'h3 == state ? _GEN_4123 : tag_1_14; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4895 = 3'h3 == state ? _GEN_4124 : tag_1_15; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4896 = 3'h3 == state ? _GEN_4125 : tag_1_16; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4897 = 3'h3 == state ? _GEN_4126 : tag_1_17; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4898 = 3'h3 == state ? _GEN_4127 : tag_1_18; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4899 = 3'h3 == state ? _GEN_4128 : tag_1_19; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4900 = 3'h3 == state ? _GEN_4129 : tag_1_20; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4901 = 3'h3 == state ? _GEN_4130 : tag_1_21; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4902 = 3'h3 == state ? _GEN_4131 : tag_1_22; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4903 = 3'h3 == state ? _GEN_4132 : tag_1_23; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4904 = 3'h3 == state ? _GEN_4133 : tag_1_24; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4905 = 3'h3 == state ? _GEN_4134 : tag_1_25; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4906 = 3'h3 == state ? _GEN_4135 : tag_1_26; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4907 = 3'h3 == state ? _GEN_4136 : tag_1_27; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4908 = 3'h3 == state ? _GEN_4137 : tag_1_28; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4909 = 3'h3 == state ? _GEN_4138 : tag_1_29; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4910 = 3'h3 == state ? _GEN_4139 : tag_1_30; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4911 = 3'h3 == state ? _GEN_4140 : tag_1_31; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4912 = 3'h3 == state ? _GEN_4141 : tag_1_32; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4913 = 3'h3 == state ? _GEN_4142 : tag_1_33; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4914 = 3'h3 == state ? _GEN_4143 : tag_1_34; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4915 = 3'h3 == state ? _GEN_4144 : tag_1_35; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4916 = 3'h3 == state ? _GEN_4145 : tag_1_36; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4917 = 3'h3 == state ? _GEN_4146 : tag_1_37; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4918 = 3'h3 == state ? _GEN_4147 : tag_1_38; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4919 = 3'h3 == state ? _GEN_4148 : tag_1_39; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4920 = 3'h3 == state ? _GEN_4149 : tag_1_40; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4921 = 3'h3 == state ? _GEN_4150 : tag_1_41; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4922 = 3'h3 == state ? _GEN_4151 : tag_1_42; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4923 = 3'h3 == state ? _GEN_4152 : tag_1_43; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4924 = 3'h3 == state ? _GEN_4153 : tag_1_44; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4925 = 3'h3 == state ? _GEN_4154 : tag_1_45; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4926 = 3'h3 == state ? _GEN_4155 : tag_1_46; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4927 = 3'h3 == state ? _GEN_4156 : tag_1_47; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4928 = 3'h3 == state ? _GEN_4157 : tag_1_48; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4929 = 3'h3 == state ? _GEN_4158 : tag_1_49; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4930 = 3'h3 == state ? _GEN_4159 : tag_1_50; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4931 = 3'h3 == state ? _GEN_4160 : tag_1_51; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4932 = 3'h3 == state ? _GEN_4161 : tag_1_52; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4933 = 3'h3 == state ? _GEN_4162 : tag_1_53; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4934 = 3'h3 == state ? _GEN_4163 : tag_1_54; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4935 = 3'h3 == state ? _GEN_4164 : tag_1_55; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4936 = 3'h3 == state ? _GEN_4165 : tag_1_56; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4937 = 3'h3 == state ? _GEN_4166 : tag_1_57; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4938 = 3'h3 == state ? _GEN_4167 : tag_1_58; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4939 = 3'h3 == state ? _GEN_4168 : tag_1_59; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4940 = 3'h3 == state ? _GEN_4169 : tag_1_60; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4941 = 3'h3 == state ? _GEN_4170 : tag_1_61; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4942 = 3'h3 == state ? _GEN_4171 : tag_1_62; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4943 = 3'h3 == state ? _GEN_4172 : tag_1_63; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4944 = 3'h3 == state ? _GEN_4173 : tag_1_64; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4945 = 3'h3 == state ? _GEN_4174 : tag_1_65; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4946 = 3'h3 == state ? _GEN_4175 : tag_1_66; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4947 = 3'h3 == state ? _GEN_4176 : tag_1_67; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4948 = 3'h3 == state ? _GEN_4177 : tag_1_68; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4949 = 3'h3 == state ? _GEN_4178 : tag_1_69; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4950 = 3'h3 == state ? _GEN_4179 : tag_1_70; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4951 = 3'h3 == state ? _GEN_4180 : tag_1_71; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4952 = 3'h3 == state ? _GEN_4181 : tag_1_72; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4953 = 3'h3 == state ? _GEN_4182 : tag_1_73; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4954 = 3'h3 == state ? _GEN_4183 : tag_1_74; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4955 = 3'h3 == state ? _GEN_4184 : tag_1_75; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4956 = 3'h3 == state ? _GEN_4185 : tag_1_76; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4957 = 3'h3 == state ? _GEN_4186 : tag_1_77; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4958 = 3'h3 == state ? _GEN_4187 : tag_1_78; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4959 = 3'h3 == state ? _GEN_4188 : tag_1_79; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4960 = 3'h3 == state ? _GEN_4189 : tag_1_80; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4961 = 3'h3 == state ? _GEN_4190 : tag_1_81; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4962 = 3'h3 == state ? _GEN_4191 : tag_1_82; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4963 = 3'h3 == state ? _GEN_4192 : tag_1_83; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4964 = 3'h3 == state ? _GEN_4193 : tag_1_84; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4965 = 3'h3 == state ? _GEN_4194 : tag_1_85; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4966 = 3'h3 == state ? _GEN_4195 : tag_1_86; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4967 = 3'h3 == state ? _GEN_4196 : tag_1_87; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4968 = 3'h3 == state ? _GEN_4197 : tag_1_88; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4969 = 3'h3 == state ? _GEN_4198 : tag_1_89; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4970 = 3'h3 == state ? _GEN_4199 : tag_1_90; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4971 = 3'h3 == state ? _GEN_4200 : tag_1_91; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4972 = 3'h3 == state ? _GEN_4201 : tag_1_92; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4973 = 3'h3 == state ? _GEN_4202 : tag_1_93; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4974 = 3'h3 == state ? _GEN_4203 : tag_1_94; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4975 = 3'h3 == state ? _GEN_4204 : tag_1_95; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4976 = 3'h3 == state ? _GEN_4205 : tag_1_96; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4977 = 3'h3 == state ? _GEN_4206 : tag_1_97; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4978 = 3'h3 == state ? _GEN_4207 : tag_1_98; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4979 = 3'h3 == state ? _GEN_4208 : tag_1_99; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4980 = 3'h3 == state ? _GEN_4209 : tag_1_100; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4981 = 3'h3 == state ? _GEN_4210 : tag_1_101; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4982 = 3'h3 == state ? _GEN_4211 : tag_1_102; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4983 = 3'h3 == state ? _GEN_4212 : tag_1_103; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4984 = 3'h3 == state ? _GEN_4213 : tag_1_104; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4985 = 3'h3 == state ? _GEN_4214 : tag_1_105; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4986 = 3'h3 == state ? _GEN_4215 : tag_1_106; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4987 = 3'h3 == state ? _GEN_4216 : tag_1_107; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4988 = 3'h3 == state ? _GEN_4217 : tag_1_108; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4989 = 3'h3 == state ? _GEN_4218 : tag_1_109; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4990 = 3'h3 == state ? _GEN_4219 : tag_1_110; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4991 = 3'h3 == state ? _GEN_4220 : tag_1_111; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4992 = 3'h3 == state ? _GEN_4221 : tag_1_112; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4993 = 3'h3 == state ? _GEN_4222 : tag_1_113; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4994 = 3'h3 == state ? _GEN_4223 : tag_1_114; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4995 = 3'h3 == state ? _GEN_4224 : tag_1_115; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4996 = 3'h3 == state ? _GEN_4225 : tag_1_116; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4997 = 3'h3 == state ? _GEN_4226 : tag_1_117; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4998 = 3'h3 == state ? _GEN_4227 : tag_1_118; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4999 = 3'h3 == state ? _GEN_4228 : tag_1_119; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5000 = 3'h3 == state ? _GEN_4229 : tag_1_120; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5001 = 3'h3 == state ? _GEN_4230 : tag_1_121; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5002 = 3'h3 == state ? _GEN_4231 : tag_1_122; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5003 = 3'h3 == state ? _GEN_4232 : tag_1_123; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5004 = 3'h3 == state ? _GEN_4233 : tag_1_124; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5005 = 3'h3 == state ? _GEN_4234 : tag_1_125; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5006 = 3'h3 == state ? _GEN_4235 : tag_1_126; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5007 = 3'h3 == state ? _GEN_4236 : tag_1_127; // @[i_cache.scala 55:18 20:24]
  wire  _GEN_5008 = 3'h3 == state ? _GEN_4237 : valid_1_0; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5009 = 3'h3 == state ? _GEN_4238 : valid_1_1; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5010 = 3'h3 == state ? _GEN_4239 : valid_1_2; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5011 = 3'h3 == state ? _GEN_4240 : valid_1_3; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5012 = 3'h3 == state ? _GEN_4241 : valid_1_4; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5013 = 3'h3 == state ? _GEN_4242 : valid_1_5; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5014 = 3'h3 == state ? _GEN_4243 : valid_1_6; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5015 = 3'h3 == state ? _GEN_4244 : valid_1_7; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5016 = 3'h3 == state ? _GEN_4245 : valid_1_8; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5017 = 3'h3 == state ? _GEN_4246 : valid_1_9; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5018 = 3'h3 == state ? _GEN_4247 : valid_1_10; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5019 = 3'h3 == state ? _GEN_4248 : valid_1_11; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5020 = 3'h3 == state ? _GEN_4249 : valid_1_12; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5021 = 3'h3 == state ? _GEN_4250 : valid_1_13; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5022 = 3'h3 == state ? _GEN_4251 : valid_1_14; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5023 = 3'h3 == state ? _GEN_4252 : valid_1_15; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5024 = 3'h3 == state ? _GEN_4253 : valid_1_16; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5025 = 3'h3 == state ? _GEN_4254 : valid_1_17; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5026 = 3'h3 == state ? _GEN_4255 : valid_1_18; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5027 = 3'h3 == state ? _GEN_4256 : valid_1_19; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5028 = 3'h3 == state ? _GEN_4257 : valid_1_20; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5029 = 3'h3 == state ? _GEN_4258 : valid_1_21; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5030 = 3'h3 == state ? _GEN_4259 : valid_1_22; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5031 = 3'h3 == state ? _GEN_4260 : valid_1_23; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5032 = 3'h3 == state ? _GEN_4261 : valid_1_24; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5033 = 3'h3 == state ? _GEN_4262 : valid_1_25; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5034 = 3'h3 == state ? _GEN_4263 : valid_1_26; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5035 = 3'h3 == state ? _GEN_4264 : valid_1_27; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5036 = 3'h3 == state ? _GEN_4265 : valid_1_28; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5037 = 3'h3 == state ? _GEN_4266 : valid_1_29; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5038 = 3'h3 == state ? _GEN_4267 : valid_1_30; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5039 = 3'h3 == state ? _GEN_4268 : valid_1_31; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5040 = 3'h3 == state ? _GEN_4269 : valid_1_32; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5041 = 3'h3 == state ? _GEN_4270 : valid_1_33; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5042 = 3'h3 == state ? _GEN_4271 : valid_1_34; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5043 = 3'h3 == state ? _GEN_4272 : valid_1_35; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5044 = 3'h3 == state ? _GEN_4273 : valid_1_36; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5045 = 3'h3 == state ? _GEN_4274 : valid_1_37; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5046 = 3'h3 == state ? _GEN_4275 : valid_1_38; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5047 = 3'h3 == state ? _GEN_4276 : valid_1_39; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5048 = 3'h3 == state ? _GEN_4277 : valid_1_40; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5049 = 3'h3 == state ? _GEN_4278 : valid_1_41; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5050 = 3'h3 == state ? _GEN_4279 : valid_1_42; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5051 = 3'h3 == state ? _GEN_4280 : valid_1_43; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5052 = 3'h3 == state ? _GEN_4281 : valid_1_44; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5053 = 3'h3 == state ? _GEN_4282 : valid_1_45; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5054 = 3'h3 == state ? _GEN_4283 : valid_1_46; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5055 = 3'h3 == state ? _GEN_4284 : valid_1_47; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5056 = 3'h3 == state ? _GEN_4285 : valid_1_48; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5057 = 3'h3 == state ? _GEN_4286 : valid_1_49; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5058 = 3'h3 == state ? _GEN_4287 : valid_1_50; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5059 = 3'h3 == state ? _GEN_4288 : valid_1_51; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5060 = 3'h3 == state ? _GEN_4289 : valid_1_52; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5061 = 3'h3 == state ? _GEN_4290 : valid_1_53; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5062 = 3'h3 == state ? _GEN_4291 : valid_1_54; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5063 = 3'h3 == state ? _GEN_4292 : valid_1_55; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5064 = 3'h3 == state ? _GEN_4293 : valid_1_56; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5065 = 3'h3 == state ? _GEN_4294 : valid_1_57; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5066 = 3'h3 == state ? _GEN_4295 : valid_1_58; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5067 = 3'h3 == state ? _GEN_4296 : valid_1_59; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5068 = 3'h3 == state ? _GEN_4297 : valid_1_60; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5069 = 3'h3 == state ? _GEN_4298 : valid_1_61; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5070 = 3'h3 == state ? _GEN_4299 : valid_1_62; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5071 = 3'h3 == state ? _GEN_4300 : valid_1_63; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5072 = 3'h3 == state ? _GEN_4301 : valid_1_64; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5073 = 3'h3 == state ? _GEN_4302 : valid_1_65; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5074 = 3'h3 == state ? _GEN_4303 : valid_1_66; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5075 = 3'h3 == state ? _GEN_4304 : valid_1_67; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5076 = 3'h3 == state ? _GEN_4305 : valid_1_68; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5077 = 3'h3 == state ? _GEN_4306 : valid_1_69; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5078 = 3'h3 == state ? _GEN_4307 : valid_1_70; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5079 = 3'h3 == state ? _GEN_4308 : valid_1_71; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5080 = 3'h3 == state ? _GEN_4309 : valid_1_72; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5081 = 3'h3 == state ? _GEN_4310 : valid_1_73; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5082 = 3'h3 == state ? _GEN_4311 : valid_1_74; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5083 = 3'h3 == state ? _GEN_4312 : valid_1_75; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5084 = 3'h3 == state ? _GEN_4313 : valid_1_76; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5085 = 3'h3 == state ? _GEN_4314 : valid_1_77; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5086 = 3'h3 == state ? _GEN_4315 : valid_1_78; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5087 = 3'h3 == state ? _GEN_4316 : valid_1_79; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5088 = 3'h3 == state ? _GEN_4317 : valid_1_80; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5089 = 3'h3 == state ? _GEN_4318 : valid_1_81; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5090 = 3'h3 == state ? _GEN_4319 : valid_1_82; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5091 = 3'h3 == state ? _GEN_4320 : valid_1_83; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5092 = 3'h3 == state ? _GEN_4321 : valid_1_84; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5093 = 3'h3 == state ? _GEN_4322 : valid_1_85; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5094 = 3'h3 == state ? _GEN_4323 : valid_1_86; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5095 = 3'h3 == state ? _GEN_4324 : valid_1_87; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5096 = 3'h3 == state ? _GEN_4325 : valid_1_88; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5097 = 3'h3 == state ? _GEN_4326 : valid_1_89; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5098 = 3'h3 == state ? _GEN_4327 : valid_1_90; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5099 = 3'h3 == state ? _GEN_4328 : valid_1_91; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5100 = 3'h3 == state ? _GEN_4329 : valid_1_92; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5101 = 3'h3 == state ? _GEN_4330 : valid_1_93; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5102 = 3'h3 == state ? _GEN_4331 : valid_1_94; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5103 = 3'h3 == state ? _GEN_4332 : valid_1_95; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5104 = 3'h3 == state ? _GEN_4333 : valid_1_96; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5105 = 3'h3 == state ? _GEN_4334 : valid_1_97; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5106 = 3'h3 == state ? _GEN_4335 : valid_1_98; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5107 = 3'h3 == state ? _GEN_4336 : valid_1_99; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5108 = 3'h3 == state ? _GEN_4337 : valid_1_100; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5109 = 3'h3 == state ? _GEN_4338 : valid_1_101; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5110 = 3'h3 == state ? _GEN_4339 : valid_1_102; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5111 = 3'h3 == state ? _GEN_4340 : valid_1_103; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5112 = 3'h3 == state ? _GEN_4341 : valid_1_104; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5113 = 3'h3 == state ? _GEN_4342 : valid_1_105; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5114 = 3'h3 == state ? _GEN_4343 : valid_1_106; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5115 = 3'h3 == state ? _GEN_4344 : valid_1_107; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5116 = 3'h3 == state ? _GEN_4345 : valid_1_108; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5117 = 3'h3 == state ? _GEN_4346 : valid_1_109; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5118 = 3'h3 == state ? _GEN_4347 : valid_1_110; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5119 = 3'h3 == state ? _GEN_4348 : valid_1_111; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5120 = 3'h3 == state ? _GEN_4349 : valid_1_112; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5121 = 3'h3 == state ? _GEN_4350 : valid_1_113; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5122 = 3'h3 == state ? _GEN_4351 : valid_1_114; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5123 = 3'h3 == state ? _GEN_4352 : valid_1_115; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5124 = 3'h3 == state ? _GEN_4353 : valid_1_116; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5125 = 3'h3 == state ? _GEN_4354 : valid_1_117; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5126 = 3'h3 == state ? _GEN_4355 : valid_1_118; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5127 = 3'h3 == state ? _GEN_4356 : valid_1_119; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5128 = 3'h3 == state ? _GEN_4357 : valid_1_120; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5129 = 3'h3 == state ? _GEN_4358 : valid_1_121; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5130 = 3'h3 == state ? _GEN_4359 : valid_1_122; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5131 = 3'h3 == state ? _GEN_4360 : valid_1_123; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5132 = 3'h3 == state ? _GEN_4361 : valid_1_124; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5133 = 3'h3 == state ? _GEN_4362 : valid_1_125; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5134 = 3'h3 == state ? _GEN_4363 : valid_1_126; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5135 = 3'h3 == state ? _GEN_4364 : valid_1_127; // @[i_cache.scala 55:18 22:26]
  wire [63:0] _GEN_7450 = 7'h1 == index ? ram_0_1 : ram_0_0; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7451 = 7'h2 == index ? ram_0_2 : _GEN_7450; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7452 = 7'h3 == index ? ram_0_3 : _GEN_7451; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7453 = 7'h4 == index ? ram_0_4 : _GEN_7452; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7454 = 7'h5 == index ? ram_0_5 : _GEN_7453; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7455 = 7'h6 == index ? ram_0_6 : _GEN_7454; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7456 = 7'h7 == index ? ram_0_7 : _GEN_7455; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7457 = 7'h8 == index ? ram_0_8 : _GEN_7456; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7458 = 7'h9 == index ? ram_0_9 : _GEN_7457; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7459 = 7'ha == index ? ram_0_10 : _GEN_7458; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7460 = 7'hb == index ? ram_0_11 : _GEN_7459; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7461 = 7'hc == index ? ram_0_12 : _GEN_7460; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7462 = 7'hd == index ? ram_0_13 : _GEN_7461; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7463 = 7'he == index ? ram_0_14 : _GEN_7462; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7464 = 7'hf == index ? ram_0_15 : _GEN_7463; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7465 = 7'h10 == index ? ram_0_16 : _GEN_7464; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7466 = 7'h11 == index ? ram_0_17 : _GEN_7465; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7467 = 7'h12 == index ? ram_0_18 : _GEN_7466; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7468 = 7'h13 == index ? ram_0_19 : _GEN_7467; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7469 = 7'h14 == index ? ram_0_20 : _GEN_7468; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7470 = 7'h15 == index ? ram_0_21 : _GEN_7469; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7471 = 7'h16 == index ? ram_0_22 : _GEN_7470; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7472 = 7'h17 == index ? ram_0_23 : _GEN_7471; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7473 = 7'h18 == index ? ram_0_24 : _GEN_7472; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7474 = 7'h19 == index ? ram_0_25 : _GEN_7473; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7475 = 7'h1a == index ? ram_0_26 : _GEN_7474; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7476 = 7'h1b == index ? ram_0_27 : _GEN_7475; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7477 = 7'h1c == index ? ram_0_28 : _GEN_7476; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7478 = 7'h1d == index ? ram_0_29 : _GEN_7477; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7479 = 7'h1e == index ? ram_0_30 : _GEN_7478; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7480 = 7'h1f == index ? ram_0_31 : _GEN_7479; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7481 = 7'h20 == index ? ram_0_32 : _GEN_7480; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7482 = 7'h21 == index ? ram_0_33 : _GEN_7481; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7483 = 7'h22 == index ? ram_0_34 : _GEN_7482; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7484 = 7'h23 == index ? ram_0_35 : _GEN_7483; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7485 = 7'h24 == index ? ram_0_36 : _GEN_7484; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7486 = 7'h25 == index ? ram_0_37 : _GEN_7485; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7487 = 7'h26 == index ? ram_0_38 : _GEN_7486; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7488 = 7'h27 == index ? ram_0_39 : _GEN_7487; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7489 = 7'h28 == index ? ram_0_40 : _GEN_7488; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7490 = 7'h29 == index ? ram_0_41 : _GEN_7489; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7491 = 7'h2a == index ? ram_0_42 : _GEN_7490; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7492 = 7'h2b == index ? ram_0_43 : _GEN_7491; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7493 = 7'h2c == index ? ram_0_44 : _GEN_7492; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7494 = 7'h2d == index ? ram_0_45 : _GEN_7493; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7495 = 7'h2e == index ? ram_0_46 : _GEN_7494; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7496 = 7'h2f == index ? ram_0_47 : _GEN_7495; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7497 = 7'h30 == index ? ram_0_48 : _GEN_7496; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7498 = 7'h31 == index ? ram_0_49 : _GEN_7497; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7499 = 7'h32 == index ? ram_0_50 : _GEN_7498; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7500 = 7'h33 == index ? ram_0_51 : _GEN_7499; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7501 = 7'h34 == index ? ram_0_52 : _GEN_7500; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7502 = 7'h35 == index ? ram_0_53 : _GEN_7501; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7503 = 7'h36 == index ? ram_0_54 : _GEN_7502; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7504 = 7'h37 == index ? ram_0_55 : _GEN_7503; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7505 = 7'h38 == index ? ram_0_56 : _GEN_7504; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7506 = 7'h39 == index ? ram_0_57 : _GEN_7505; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7507 = 7'h3a == index ? ram_0_58 : _GEN_7506; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7508 = 7'h3b == index ? ram_0_59 : _GEN_7507; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7509 = 7'h3c == index ? ram_0_60 : _GEN_7508; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7510 = 7'h3d == index ? ram_0_61 : _GEN_7509; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7511 = 7'h3e == index ? ram_0_62 : _GEN_7510; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7512 = 7'h3f == index ? ram_0_63 : _GEN_7511; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7513 = 7'h40 == index ? ram_0_64 : _GEN_7512; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7514 = 7'h41 == index ? ram_0_65 : _GEN_7513; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7515 = 7'h42 == index ? ram_0_66 : _GEN_7514; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7516 = 7'h43 == index ? ram_0_67 : _GEN_7515; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7517 = 7'h44 == index ? ram_0_68 : _GEN_7516; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7518 = 7'h45 == index ? ram_0_69 : _GEN_7517; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7519 = 7'h46 == index ? ram_0_70 : _GEN_7518; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7520 = 7'h47 == index ? ram_0_71 : _GEN_7519; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7521 = 7'h48 == index ? ram_0_72 : _GEN_7520; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7522 = 7'h49 == index ? ram_0_73 : _GEN_7521; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7523 = 7'h4a == index ? ram_0_74 : _GEN_7522; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7524 = 7'h4b == index ? ram_0_75 : _GEN_7523; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7525 = 7'h4c == index ? ram_0_76 : _GEN_7524; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7526 = 7'h4d == index ? ram_0_77 : _GEN_7525; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7527 = 7'h4e == index ? ram_0_78 : _GEN_7526; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7528 = 7'h4f == index ? ram_0_79 : _GEN_7527; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7529 = 7'h50 == index ? ram_0_80 : _GEN_7528; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7530 = 7'h51 == index ? ram_0_81 : _GEN_7529; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7531 = 7'h52 == index ? ram_0_82 : _GEN_7530; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7532 = 7'h53 == index ? ram_0_83 : _GEN_7531; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7533 = 7'h54 == index ? ram_0_84 : _GEN_7532; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7534 = 7'h55 == index ? ram_0_85 : _GEN_7533; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7535 = 7'h56 == index ? ram_0_86 : _GEN_7534; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7536 = 7'h57 == index ? ram_0_87 : _GEN_7535; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7537 = 7'h58 == index ? ram_0_88 : _GEN_7536; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7538 = 7'h59 == index ? ram_0_89 : _GEN_7537; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7539 = 7'h5a == index ? ram_0_90 : _GEN_7538; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7540 = 7'h5b == index ? ram_0_91 : _GEN_7539; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7541 = 7'h5c == index ? ram_0_92 : _GEN_7540; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7542 = 7'h5d == index ? ram_0_93 : _GEN_7541; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7543 = 7'h5e == index ? ram_0_94 : _GEN_7542; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7544 = 7'h5f == index ? ram_0_95 : _GEN_7543; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7545 = 7'h60 == index ? ram_0_96 : _GEN_7544; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7546 = 7'h61 == index ? ram_0_97 : _GEN_7545; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7547 = 7'h62 == index ? ram_0_98 : _GEN_7546; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7548 = 7'h63 == index ? ram_0_99 : _GEN_7547; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7549 = 7'h64 == index ? ram_0_100 : _GEN_7548; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7550 = 7'h65 == index ? ram_0_101 : _GEN_7549; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7551 = 7'h66 == index ? ram_0_102 : _GEN_7550; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7552 = 7'h67 == index ? ram_0_103 : _GEN_7551; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7553 = 7'h68 == index ? ram_0_104 : _GEN_7552; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7554 = 7'h69 == index ? ram_0_105 : _GEN_7553; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7555 = 7'h6a == index ? ram_0_106 : _GEN_7554; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7556 = 7'h6b == index ? ram_0_107 : _GEN_7555; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7557 = 7'h6c == index ? ram_0_108 : _GEN_7556; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7558 = 7'h6d == index ? ram_0_109 : _GEN_7557; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7559 = 7'h6e == index ? ram_0_110 : _GEN_7558; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7560 = 7'h6f == index ? ram_0_111 : _GEN_7559; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7561 = 7'h70 == index ? ram_0_112 : _GEN_7560; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7562 = 7'h71 == index ? ram_0_113 : _GEN_7561; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7563 = 7'h72 == index ? ram_0_114 : _GEN_7562; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7564 = 7'h73 == index ? ram_0_115 : _GEN_7563; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7565 = 7'h74 == index ? ram_0_116 : _GEN_7564; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7566 = 7'h75 == index ? ram_0_117 : _GEN_7565; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7567 = 7'h76 == index ? ram_0_118 : _GEN_7566; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7568 = 7'h77 == index ? ram_0_119 : _GEN_7567; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7569 = 7'h78 == index ? ram_0_120 : _GEN_7568; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7570 = 7'h79 == index ? ram_0_121 : _GEN_7569; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7571 = 7'h7a == index ? ram_0_122 : _GEN_7570; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7572 = 7'h7b == index ? ram_0_123 : _GEN_7571; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7573 = 7'h7c == index ? ram_0_124 : _GEN_7572; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7574 = 7'h7d == index ? ram_0_125 : _GEN_7573; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7575 = 7'h7e == index ? ram_0_126 : _GEN_7574; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7576 = 7'h7f == index ? ram_0_127 : _GEN_7575; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7578 = 7'h1 == index ? ram_1_1 : ram_1_0; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7579 = 7'h2 == index ? ram_1_2 : _GEN_7578; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7580 = 7'h3 == index ? ram_1_3 : _GEN_7579; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7581 = 7'h4 == index ? ram_1_4 : _GEN_7580; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7582 = 7'h5 == index ? ram_1_5 : _GEN_7581; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7583 = 7'h6 == index ? ram_1_6 : _GEN_7582; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7584 = 7'h7 == index ? ram_1_7 : _GEN_7583; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7585 = 7'h8 == index ? ram_1_8 : _GEN_7584; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7586 = 7'h9 == index ? ram_1_9 : _GEN_7585; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7587 = 7'ha == index ? ram_1_10 : _GEN_7586; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7588 = 7'hb == index ? ram_1_11 : _GEN_7587; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7589 = 7'hc == index ? ram_1_12 : _GEN_7588; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7590 = 7'hd == index ? ram_1_13 : _GEN_7589; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7591 = 7'he == index ? ram_1_14 : _GEN_7590; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7592 = 7'hf == index ? ram_1_15 : _GEN_7591; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7593 = 7'h10 == index ? ram_1_16 : _GEN_7592; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7594 = 7'h11 == index ? ram_1_17 : _GEN_7593; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7595 = 7'h12 == index ? ram_1_18 : _GEN_7594; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7596 = 7'h13 == index ? ram_1_19 : _GEN_7595; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7597 = 7'h14 == index ? ram_1_20 : _GEN_7596; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7598 = 7'h15 == index ? ram_1_21 : _GEN_7597; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7599 = 7'h16 == index ? ram_1_22 : _GEN_7598; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7600 = 7'h17 == index ? ram_1_23 : _GEN_7599; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7601 = 7'h18 == index ? ram_1_24 : _GEN_7600; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7602 = 7'h19 == index ? ram_1_25 : _GEN_7601; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7603 = 7'h1a == index ? ram_1_26 : _GEN_7602; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7604 = 7'h1b == index ? ram_1_27 : _GEN_7603; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7605 = 7'h1c == index ? ram_1_28 : _GEN_7604; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7606 = 7'h1d == index ? ram_1_29 : _GEN_7605; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7607 = 7'h1e == index ? ram_1_30 : _GEN_7606; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7608 = 7'h1f == index ? ram_1_31 : _GEN_7607; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7609 = 7'h20 == index ? ram_1_32 : _GEN_7608; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7610 = 7'h21 == index ? ram_1_33 : _GEN_7609; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7611 = 7'h22 == index ? ram_1_34 : _GEN_7610; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7612 = 7'h23 == index ? ram_1_35 : _GEN_7611; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7613 = 7'h24 == index ? ram_1_36 : _GEN_7612; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7614 = 7'h25 == index ? ram_1_37 : _GEN_7613; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7615 = 7'h26 == index ? ram_1_38 : _GEN_7614; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7616 = 7'h27 == index ? ram_1_39 : _GEN_7615; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7617 = 7'h28 == index ? ram_1_40 : _GEN_7616; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7618 = 7'h29 == index ? ram_1_41 : _GEN_7617; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7619 = 7'h2a == index ? ram_1_42 : _GEN_7618; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7620 = 7'h2b == index ? ram_1_43 : _GEN_7619; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7621 = 7'h2c == index ? ram_1_44 : _GEN_7620; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7622 = 7'h2d == index ? ram_1_45 : _GEN_7621; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7623 = 7'h2e == index ? ram_1_46 : _GEN_7622; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7624 = 7'h2f == index ? ram_1_47 : _GEN_7623; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7625 = 7'h30 == index ? ram_1_48 : _GEN_7624; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7626 = 7'h31 == index ? ram_1_49 : _GEN_7625; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7627 = 7'h32 == index ? ram_1_50 : _GEN_7626; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7628 = 7'h33 == index ? ram_1_51 : _GEN_7627; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7629 = 7'h34 == index ? ram_1_52 : _GEN_7628; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7630 = 7'h35 == index ? ram_1_53 : _GEN_7629; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7631 = 7'h36 == index ? ram_1_54 : _GEN_7630; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7632 = 7'h37 == index ? ram_1_55 : _GEN_7631; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7633 = 7'h38 == index ? ram_1_56 : _GEN_7632; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7634 = 7'h39 == index ? ram_1_57 : _GEN_7633; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7635 = 7'h3a == index ? ram_1_58 : _GEN_7634; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7636 = 7'h3b == index ? ram_1_59 : _GEN_7635; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7637 = 7'h3c == index ? ram_1_60 : _GEN_7636; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7638 = 7'h3d == index ? ram_1_61 : _GEN_7637; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7639 = 7'h3e == index ? ram_1_62 : _GEN_7638; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7640 = 7'h3f == index ? ram_1_63 : _GEN_7639; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7641 = 7'h40 == index ? ram_1_64 : _GEN_7640; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7642 = 7'h41 == index ? ram_1_65 : _GEN_7641; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7643 = 7'h42 == index ? ram_1_66 : _GEN_7642; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7644 = 7'h43 == index ? ram_1_67 : _GEN_7643; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7645 = 7'h44 == index ? ram_1_68 : _GEN_7644; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7646 = 7'h45 == index ? ram_1_69 : _GEN_7645; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7647 = 7'h46 == index ? ram_1_70 : _GEN_7646; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7648 = 7'h47 == index ? ram_1_71 : _GEN_7647; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7649 = 7'h48 == index ? ram_1_72 : _GEN_7648; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7650 = 7'h49 == index ? ram_1_73 : _GEN_7649; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7651 = 7'h4a == index ? ram_1_74 : _GEN_7650; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7652 = 7'h4b == index ? ram_1_75 : _GEN_7651; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7653 = 7'h4c == index ? ram_1_76 : _GEN_7652; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7654 = 7'h4d == index ? ram_1_77 : _GEN_7653; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7655 = 7'h4e == index ? ram_1_78 : _GEN_7654; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7656 = 7'h4f == index ? ram_1_79 : _GEN_7655; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7657 = 7'h50 == index ? ram_1_80 : _GEN_7656; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7658 = 7'h51 == index ? ram_1_81 : _GEN_7657; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7659 = 7'h52 == index ? ram_1_82 : _GEN_7658; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7660 = 7'h53 == index ? ram_1_83 : _GEN_7659; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7661 = 7'h54 == index ? ram_1_84 : _GEN_7660; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7662 = 7'h55 == index ? ram_1_85 : _GEN_7661; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7663 = 7'h56 == index ? ram_1_86 : _GEN_7662; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7664 = 7'h57 == index ? ram_1_87 : _GEN_7663; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7665 = 7'h58 == index ? ram_1_88 : _GEN_7664; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7666 = 7'h59 == index ? ram_1_89 : _GEN_7665; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7667 = 7'h5a == index ? ram_1_90 : _GEN_7666; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7668 = 7'h5b == index ? ram_1_91 : _GEN_7667; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7669 = 7'h5c == index ? ram_1_92 : _GEN_7668; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7670 = 7'h5d == index ? ram_1_93 : _GEN_7669; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7671 = 7'h5e == index ? ram_1_94 : _GEN_7670; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7672 = 7'h5f == index ? ram_1_95 : _GEN_7671; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7673 = 7'h60 == index ? ram_1_96 : _GEN_7672; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7674 = 7'h61 == index ? ram_1_97 : _GEN_7673; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7675 = 7'h62 == index ? ram_1_98 : _GEN_7674; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7676 = 7'h63 == index ? ram_1_99 : _GEN_7675; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7677 = 7'h64 == index ? ram_1_100 : _GEN_7676; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7678 = 7'h65 == index ? ram_1_101 : _GEN_7677; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7679 = 7'h66 == index ? ram_1_102 : _GEN_7678; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7680 = 7'h67 == index ? ram_1_103 : _GEN_7679; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7681 = 7'h68 == index ? ram_1_104 : _GEN_7680; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7682 = 7'h69 == index ? ram_1_105 : _GEN_7681; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7683 = 7'h6a == index ? ram_1_106 : _GEN_7682; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7684 = 7'h6b == index ? ram_1_107 : _GEN_7683; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7685 = 7'h6c == index ? ram_1_108 : _GEN_7684; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7686 = 7'h6d == index ? ram_1_109 : _GEN_7685; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7687 = 7'h6e == index ? ram_1_110 : _GEN_7686; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7688 = 7'h6f == index ? ram_1_111 : _GEN_7687; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7689 = 7'h70 == index ? ram_1_112 : _GEN_7688; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7690 = 7'h71 == index ? ram_1_113 : _GEN_7689; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7691 = 7'h72 == index ? ram_1_114 : _GEN_7690; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7692 = 7'h73 == index ? ram_1_115 : _GEN_7691; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7693 = 7'h74 == index ? ram_1_116 : _GEN_7692; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7694 = 7'h75 == index ? ram_1_117 : _GEN_7693; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7695 = 7'h76 == index ? ram_1_118 : _GEN_7694; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7696 = 7'h77 == index ? ram_1_119 : _GEN_7695; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7697 = 7'h78 == index ? ram_1_120 : _GEN_7696; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7698 = 7'h79 == index ? ram_1_121 : _GEN_7697; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7699 = 7'h7a == index ? ram_1_122 : _GEN_7698; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7700 = 7'h7b == index ? ram_1_123 : _GEN_7699; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7701 = 7'h7c == index ? ram_1_124 : _GEN_7700; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7702 = 7'h7d == index ? ram_1_125 : _GEN_7701; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7703 = 7'h7e == index ? ram_1_126 : _GEN_7702; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7704 = 7'h7f == index ? ram_1_127 : _GEN_7703; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7705 = way1_hit ? _GEN_7704 : 64'h0; // @[i_cache.scala 148:33 149:33 156:33]
  wire [63:0] _GEN_7709 = way0_hit ? _GEN_7576 : _GEN_7705; // @[i_cache.scala 140:23 141:33]
  wire  _GEN_7711 = way0_hit | way1_hit; // @[i_cache.scala 140:23 143:34]
  wire  _T_18 = state == 3'h2; // @[i_cache.scala 163:21]
  wire  _GEN_7722 = state == 3'h1 ? 1'h0 : _T_18; // @[i_cache.scala 130:31 131:27]
  wire  _GEN_7724 = state == 3'h1 ? 1'h0 : io_from_ifu_rready; // @[i_cache.scala 130:31 133:26]
  wire [63:0] _GEN_7726 = state == 3'h1 ? _GEN_7709 : 64'h0; // @[i_cache.scala 130:31]
  wire  _GEN_7728 = state == 3'h1 & _GEN_7711; // @[i_cache.scala 130:31]
  assign io_to_ifu_rdata = state == 3'h0 ? 64'h0 : _GEN_7726; // @[i_cache.scala 114:23 115:25]
  assign io_to_ifu_rvalid = state == 3'h0 ? 1'h0 : _GEN_7728; // @[i_cache.scala 114:23 117:26]
  assign io_to_axi_araddr = io_from_ifu_araddr; // @[i_cache.scala 114:23 122:26]
  assign io_to_axi_arvalid = state == 3'h0 ? 1'h0 : _GEN_7722; // @[i_cache.scala 114:23 121:27]
  assign io_to_axi_rready = state == 3'h0 ? io_from_ifu_rready : _GEN_7724; // @[i_cache.scala 114:23 123:26]
  always @(posedge clock) begin
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_0 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_0 <= _GEN_4367;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_1 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_1 <= _GEN_4368;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_2 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_2 <= _GEN_4369;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_3 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_3 <= _GEN_4370;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_4 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_4 <= _GEN_4371;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_5 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_5 <= _GEN_4372;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_6 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_6 <= _GEN_4373;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_7 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_7 <= _GEN_4374;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_8 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_8 <= _GEN_4375;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_9 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_9 <= _GEN_4376;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_10 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_10 <= _GEN_4377;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_11 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_11 <= _GEN_4378;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_12 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_12 <= _GEN_4379;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_13 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_13 <= _GEN_4380;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_14 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_14 <= _GEN_4381;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_15 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_15 <= _GEN_4382;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_16 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_16 <= _GEN_4383;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_17 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_17 <= _GEN_4384;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_18 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_18 <= _GEN_4385;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_19 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_19 <= _GEN_4386;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_20 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_20 <= _GEN_4387;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_21 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_21 <= _GEN_4388;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_22 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_22 <= _GEN_4389;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_23 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_23 <= _GEN_4390;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_24 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_24 <= _GEN_4391;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_25 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_25 <= _GEN_4392;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_26 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_26 <= _GEN_4393;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_27 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_27 <= _GEN_4394;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_28 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_28 <= _GEN_4395;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_29 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_29 <= _GEN_4396;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_30 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_30 <= _GEN_4397;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_31 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_31 <= _GEN_4398;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_32 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_32 <= _GEN_4399;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_33 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_33 <= _GEN_4400;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_34 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_34 <= _GEN_4401;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_35 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_35 <= _GEN_4402;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_36 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_36 <= _GEN_4403;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_37 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_37 <= _GEN_4404;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_38 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_38 <= _GEN_4405;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_39 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_39 <= _GEN_4406;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_40 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_40 <= _GEN_4407;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_41 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_41 <= _GEN_4408;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_42 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_42 <= _GEN_4409;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_43 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_43 <= _GEN_4410;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_44 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_44 <= _GEN_4411;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_45 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_45 <= _GEN_4412;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_46 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_46 <= _GEN_4413;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_47 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_47 <= _GEN_4414;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_48 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_48 <= _GEN_4415;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_49 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_49 <= _GEN_4416;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_50 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_50 <= _GEN_4417;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_51 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_51 <= _GEN_4418;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_52 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_52 <= _GEN_4419;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_53 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_53 <= _GEN_4420;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_54 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_54 <= _GEN_4421;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_55 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_55 <= _GEN_4422;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_56 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_56 <= _GEN_4423;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_57 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_57 <= _GEN_4424;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_58 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_58 <= _GEN_4425;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_59 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_59 <= _GEN_4426;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_60 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_60 <= _GEN_4427;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_61 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_61 <= _GEN_4428;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_62 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_62 <= _GEN_4429;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_63 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_63 <= _GEN_4430;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_64 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_64 <= _GEN_4431;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_65 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_65 <= _GEN_4432;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_66 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_66 <= _GEN_4433;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_67 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_67 <= _GEN_4434;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_68 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_68 <= _GEN_4435;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_69 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_69 <= _GEN_4436;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_70 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_70 <= _GEN_4437;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_71 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_71 <= _GEN_4438;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_72 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_72 <= _GEN_4439;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_73 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_73 <= _GEN_4440;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_74 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_74 <= _GEN_4441;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_75 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_75 <= _GEN_4442;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_76 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_76 <= _GEN_4443;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_77 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_77 <= _GEN_4444;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_78 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_78 <= _GEN_4445;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_79 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_79 <= _GEN_4446;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_80 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_80 <= _GEN_4447;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_81 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_81 <= _GEN_4448;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_82 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_82 <= _GEN_4449;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_83 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_83 <= _GEN_4450;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_84 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_84 <= _GEN_4451;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_85 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_85 <= _GEN_4452;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_86 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_86 <= _GEN_4453;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_87 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_87 <= _GEN_4454;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_88 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_88 <= _GEN_4455;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_89 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_89 <= _GEN_4456;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_90 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_90 <= _GEN_4457;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_91 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_91 <= _GEN_4458;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_92 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_92 <= _GEN_4459;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_93 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_93 <= _GEN_4460;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_94 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_94 <= _GEN_4461;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_95 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_95 <= _GEN_4462;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_96 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_96 <= _GEN_4463;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_97 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_97 <= _GEN_4464;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_98 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_98 <= _GEN_4465;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_99 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_99 <= _GEN_4466;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_100 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_100 <= _GEN_4467;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_101 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_101 <= _GEN_4468;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_102 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_102 <= _GEN_4469;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_103 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_103 <= _GEN_4470;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_104 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_104 <= _GEN_4471;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_105 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_105 <= _GEN_4472;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_106 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_106 <= _GEN_4473;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_107 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_107 <= _GEN_4474;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_108 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_108 <= _GEN_4475;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_109 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_109 <= _GEN_4476;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_110 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_110 <= _GEN_4477;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_111 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_111 <= _GEN_4478;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_112 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_112 <= _GEN_4479;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_113 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_113 <= _GEN_4480;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_114 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_114 <= _GEN_4481;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_115 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_115 <= _GEN_4482;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_116 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_116 <= _GEN_4483;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_117 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_117 <= _GEN_4484;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_118 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_118 <= _GEN_4485;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_119 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_119 <= _GEN_4486;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_120 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_120 <= _GEN_4487;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_121 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_121 <= _GEN_4488;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_122 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_122 <= _GEN_4489;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_123 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_123 <= _GEN_4490;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_124 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_124 <= _GEN_4491;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_125 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_125 <= _GEN_4492;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_126 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_126 <= _GEN_4493;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_127 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_127 <= _GEN_4494;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_0 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_0 <= _GEN_4752;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_1 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_1 <= _GEN_4753;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_2 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_2 <= _GEN_4754;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_3 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_3 <= _GEN_4755;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_4 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_4 <= _GEN_4756;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_5 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_5 <= _GEN_4757;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_6 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_6 <= _GEN_4758;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_7 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_7 <= _GEN_4759;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_8 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_8 <= _GEN_4760;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_9 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_9 <= _GEN_4761;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_10 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_10 <= _GEN_4762;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_11 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_11 <= _GEN_4763;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_12 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_12 <= _GEN_4764;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_13 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_13 <= _GEN_4765;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_14 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_14 <= _GEN_4766;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_15 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_15 <= _GEN_4767;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_16 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_16 <= _GEN_4768;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_17 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_17 <= _GEN_4769;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_18 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_18 <= _GEN_4770;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_19 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_19 <= _GEN_4771;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_20 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_20 <= _GEN_4772;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_21 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_21 <= _GEN_4773;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_22 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_22 <= _GEN_4774;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_23 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_23 <= _GEN_4775;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_24 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_24 <= _GEN_4776;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_25 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_25 <= _GEN_4777;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_26 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_26 <= _GEN_4778;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_27 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_27 <= _GEN_4779;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_28 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_28 <= _GEN_4780;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_29 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_29 <= _GEN_4781;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_30 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_30 <= _GEN_4782;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_31 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_31 <= _GEN_4783;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_32 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_32 <= _GEN_4784;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_33 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_33 <= _GEN_4785;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_34 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_34 <= _GEN_4786;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_35 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_35 <= _GEN_4787;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_36 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_36 <= _GEN_4788;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_37 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_37 <= _GEN_4789;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_38 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_38 <= _GEN_4790;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_39 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_39 <= _GEN_4791;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_40 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_40 <= _GEN_4792;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_41 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_41 <= _GEN_4793;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_42 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_42 <= _GEN_4794;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_43 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_43 <= _GEN_4795;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_44 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_44 <= _GEN_4796;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_45 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_45 <= _GEN_4797;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_46 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_46 <= _GEN_4798;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_47 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_47 <= _GEN_4799;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_48 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_48 <= _GEN_4800;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_49 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_49 <= _GEN_4801;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_50 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_50 <= _GEN_4802;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_51 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_51 <= _GEN_4803;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_52 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_52 <= _GEN_4804;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_53 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_53 <= _GEN_4805;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_54 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_54 <= _GEN_4806;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_55 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_55 <= _GEN_4807;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_56 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_56 <= _GEN_4808;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_57 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_57 <= _GEN_4809;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_58 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_58 <= _GEN_4810;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_59 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_59 <= _GEN_4811;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_60 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_60 <= _GEN_4812;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_61 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_61 <= _GEN_4813;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_62 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_62 <= _GEN_4814;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_63 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_63 <= _GEN_4815;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_64 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_64 <= _GEN_4816;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_65 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_65 <= _GEN_4817;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_66 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_66 <= _GEN_4818;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_67 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_67 <= _GEN_4819;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_68 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_68 <= _GEN_4820;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_69 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_69 <= _GEN_4821;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_70 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_70 <= _GEN_4822;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_71 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_71 <= _GEN_4823;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_72 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_72 <= _GEN_4824;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_73 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_73 <= _GEN_4825;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_74 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_74 <= _GEN_4826;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_75 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_75 <= _GEN_4827;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_76 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_76 <= _GEN_4828;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_77 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_77 <= _GEN_4829;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_78 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_78 <= _GEN_4830;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_79 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_79 <= _GEN_4831;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_80 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_80 <= _GEN_4832;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_81 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_81 <= _GEN_4833;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_82 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_82 <= _GEN_4834;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_83 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_83 <= _GEN_4835;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_84 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_84 <= _GEN_4836;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_85 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_85 <= _GEN_4837;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_86 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_86 <= _GEN_4838;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_87 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_87 <= _GEN_4839;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_88 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_88 <= _GEN_4840;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_89 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_89 <= _GEN_4841;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_90 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_90 <= _GEN_4842;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_91 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_91 <= _GEN_4843;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_92 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_92 <= _GEN_4844;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_93 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_93 <= _GEN_4845;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_94 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_94 <= _GEN_4846;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_95 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_95 <= _GEN_4847;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_96 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_96 <= _GEN_4848;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_97 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_97 <= _GEN_4849;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_98 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_98 <= _GEN_4850;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_99 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_99 <= _GEN_4851;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_100 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_100 <= _GEN_4852;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_101 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_101 <= _GEN_4853;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_102 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_102 <= _GEN_4854;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_103 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_103 <= _GEN_4855;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_104 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_104 <= _GEN_4856;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_105 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_105 <= _GEN_4857;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_106 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_106 <= _GEN_4858;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_107 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_107 <= _GEN_4859;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_108 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_108 <= _GEN_4860;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_109 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_109 <= _GEN_4861;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_110 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_110 <= _GEN_4862;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_111 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_111 <= _GEN_4863;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_112 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_112 <= _GEN_4864;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_113 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_113 <= _GEN_4865;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_114 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_114 <= _GEN_4866;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_115 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_115 <= _GEN_4867;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_116 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_116 <= _GEN_4868;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_117 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_117 <= _GEN_4869;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_118 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_118 <= _GEN_4870;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_119 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_119 <= _GEN_4871;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_120 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_120 <= _GEN_4872;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_121 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_121 <= _GEN_4873;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_122 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_122 <= _GEN_4874;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_123 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_123 <= _GEN_4875;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_124 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_124 <= _GEN_4876;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_125 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_125 <= _GEN_4877;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_126 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_126 <= _GEN_4878;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_127 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_127 <= _GEN_4879;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_0 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_0 <= _GEN_4495;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_1 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_1 <= _GEN_4496;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_2 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_2 <= _GEN_4497;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_3 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_3 <= _GEN_4498;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_4 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_4 <= _GEN_4499;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_5 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_5 <= _GEN_4500;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_6 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_6 <= _GEN_4501;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_7 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_7 <= _GEN_4502;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_8 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_8 <= _GEN_4503;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_9 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_9 <= _GEN_4504;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_10 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_10 <= _GEN_4505;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_11 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_11 <= _GEN_4506;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_12 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_12 <= _GEN_4507;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_13 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_13 <= _GEN_4508;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_14 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_14 <= _GEN_4509;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_15 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_15 <= _GEN_4510;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_16 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_16 <= _GEN_4511;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_17 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_17 <= _GEN_4512;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_18 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_18 <= _GEN_4513;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_19 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_19 <= _GEN_4514;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_20 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_20 <= _GEN_4515;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_21 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_21 <= _GEN_4516;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_22 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_22 <= _GEN_4517;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_23 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_23 <= _GEN_4518;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_24 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_24 <= _GEN_4519;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_25 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_25 <= _GEN_4520;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_26 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_26 <= _GEN_4521;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_27 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_27 <= _GEN_4522;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_28 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_28 <= _GEN_4523;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_29 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_29 <= _GEN_4524;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_30 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_30 <= _GEN_4525;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_31 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_31 <= _GEN_4526;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_32 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_32 <= _GEN_4527;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_33 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_33 <= _GEN_4528;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_34 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_34 <= _GEN_4529;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_35 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_35 <= _GEN_4530;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_36 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_36 <= _GEN_4531;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_37 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_37 <= _GEN_4532;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_38 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_38 <= _GEN_4533;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_39 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_39 <= _GEN_4534;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_40 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_40 <= _GEN_4535;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_41 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_41 <= _GEN_4536;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_42 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_42 <= _GEN_4537;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_43 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_43 <= _GEN_4538;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_44 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_44 <= _GEN_4539;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_45 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_45 <= _GEN_4540;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_46 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_46 <= _GEN_4541;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_47 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_47 <= _GEN_4542;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_48 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_48 <= _GEN_4543;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_49 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_49 <= _GEN_4544;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_50 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_50 <= _GEN_4545;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_51 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_51 <= _GEN_4546;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_52 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_52 <= _GEN_4547;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_53 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_53 <= _GEN_4548;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_54 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_54 <= _GEN_4549;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_55 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_55 <= _GEN_4550;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_56 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_56 <= _GEN_4551;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_57 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_57 <= _GEN_4552;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_58 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_58 <= _GEN_4553;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_59 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_59 <= _GEN_4554;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_60 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_60 <= _GEN_4555;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_61 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_61 <= _GEN_4556;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_62 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_62 <= _GEN_4557;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_63 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_63 <= _GEN_4558;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_64 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_64 <= _GEN_4559;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_65 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_65 <= _GEN_4560;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_66 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_66 <= _GEN_4561;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_67 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_67 <= _GEN_4562;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_68 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_68 <= _GEN_4563;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_69 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_69 <= _GEN_4564;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_70 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_70 <= _GEN_4565;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_71 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_71 <= _GEN_4566;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_72 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_72 <= _GEN_4567;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_73 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_73 <= _GEN_4568;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_74 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_74 <= _GEN_4569;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_75 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_75 <= _GEN_4570;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_76 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_76 <= _GEN_4571;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_77 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_77 <= _GEN_4572;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_78 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_78 <= _GEN_4573;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_79 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_79 <= _GEN_4574;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_80 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_80 <= _GEN_4575;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_81 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_81 <= _GEN_4576;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_82 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_82 <= _GEN_4577;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_83 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_83 <= _GEN_4578;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_84 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_84 <= _GEN_4579;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_85 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_85 <= _GEN_4580;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_86 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_86 <= _GEN_4581;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_87 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_87 <= _GEN_4582;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_88 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_88 <= _GEN_4583;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_89 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_89 <= _GEN_4584;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_90 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_90 <= _GEN_4585;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_91 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_91 <= _GEN_4586;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_92 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_92 <= _GEN_4587;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_93 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_93 <= _GEN_4588;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_94 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_94 <= _GEN_4589;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_95 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_95 <= _GEN_4590;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_96 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_96 <= _GEN_4591;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_97 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_97 <= _GEN_4592;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_98 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_98 <= _GEN_4593;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_99 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_99 <= _GEN_4594;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_100 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_100 <= _GEN_4595;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_101 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_101 <= _GEN_4596;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_102 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_102 <= _GEN_4597;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_103 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_103 <= _GEN_4598;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_104 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_104 <= _GEN_4599;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_105 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_105 <= _GEN_4600;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_106 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_106 <= _GEN_4601;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_107 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_107 <= _GEN_4602;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_108 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_108 <= _GEN_4603;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_109 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_109 <= _GEN_4604;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_110 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_110 <= _GEN_4605;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_111 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_111 <= _GEN_4606;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_112 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_112 <= _GEN_4607;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_113 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_113 <= _GEN_4608;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_114 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_114 <= _GEN_4609;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_115 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_115 <= _GEN_4610;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_116 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_116 <= _GEN_4611;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_117 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_117 <= _GEN_4612;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_118 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_118 <= _GEN_4613;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_119 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_119 <= _GEN_4614;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_120 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_120 <= _GEN_4615;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_121 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_121 <= _GEN_4616;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_122 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_122 <= _GEN_4617;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_123 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_123 <= _GEN_4618;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_124 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_124 <= _GEN_4619;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_125 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_125 <= _GEN_4620;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_126 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_126 <= _GEN_4621;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_127 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_127 <= _GEN_4622;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_0 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_0 <= _GEN_4880;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_1 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_1 <= _GEN_4881;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_2 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_2 <= _GEN_4882;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_3 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_3 <= _GEN_4883;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_4 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_4 <= _GEN_4884;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_5 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_5 <= _GEN_4885;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_6 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_6 <= _GEN_4886;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_7 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_7 <= _GEN_4887;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_8 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_8 <= _GEN_4888;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_9 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_9 <= _GEN_4889;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_10 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_10 <= _GEN_4890;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_11 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_11 <= _GEN_4891;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_12 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_12 <= _GEN_4892;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_13 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_13 <= _GEN_4893;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_14 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_14 <= _GEN_4894;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_15 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_15 <= _GEN_4895;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_16 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_16 <= _GEN_4896;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_17 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_17 <= _GEN_4897;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_18 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_18 <= _GEN_4898;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_19 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_19 <= _GEN_4899;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_20 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_20 <= _GEN_4900;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_21 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_21 <= _GEN_4901;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_22 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_22 <= _GEN_4902;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_23 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_23 <= _GEN_4903;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_24 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_24 <= _GEN_4904;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_25 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_25 <= _GEN_4905;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_26 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_26 <= _GEN_4906;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_27 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_27 <= _GEN_4907;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_28 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_28 <= _GEN_4908;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_29 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_29 <= _GEN_4909;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_30 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_30 <= _GEN_4910;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_31 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_31 <= _GEN_4911;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_32 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_32 <= _GEN_4912;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_33 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_33 <= _GEN_4913;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_34 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_34 <= _GEN_4914;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_35 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_35 <= _GEN_4915;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_36 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_36 <= _GEN_4916;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_37 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_37 <= _GEN_4917;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_38 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_38 <= _GEN_4918;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_39 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_39 <= _GEN_4919;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_40 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_40 <= _GEN_4920;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_41 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_41 <= _GEN_4921;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_42 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_42 <= _GEN_4922;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_43 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_43 <= _GEN_4923;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_44 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_44 <= _GEN_4924;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_45 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_45 <= _GEN_4925;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_46 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_46 <= _GEN_4926;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_47 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_47 <= _GEN_4927;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_48 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_48 <= _GEN_4928;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_49 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_49 <= _GEN_4929;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_50 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_50 <= _GEN_4930;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_51 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_51 <= _GEN_4931;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_52 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_52 <= _GEN_4932;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_53 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_53 <= _GEN_4933;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_54 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_54 <= _GEN_4934;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_55 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_55 <= _GEN_4935;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_56 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_56 <= _GEN_4936;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_57 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_57 <= _GEN_4937;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_58 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_58 <= _GEN_4938;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_59 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_59 <= _GEN_4939;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_60 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_60 <= _GEN_4940;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_61 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_61 <= _GEN_4941;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_62 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_62 <= _GEN_4942;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_63 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_63 <= _GEN_4943;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_64 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_64 <= _GEN_4944;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_65 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_65 <= _GEN_4945;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_66 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_66 <= _GEN_4946;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_67 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_67 <= _GEN_4947;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_68 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_68 <= _GEN_4948;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_69 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_69 <= _GEN_4949;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_70 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_70 <= _GEN_4950;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_71 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_71 <= _GEN_4951;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_72 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_72 <= _GEN_4952;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_73 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_73 <= _GEN_4953;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_74 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_74 <= _GEN_4954;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_75 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_75 <= _GEN_4955;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_76 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_76 <= _GEN_4956;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_77 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_77 <= _GEN_4957;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_78 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_78 <= _GEN_4958;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_79 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_79 <= _GEN_4959;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_80 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_80 <= _GEN_4960;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_81 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_81 <= _GEN_4961;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_82 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_82 <= _GEN_4962;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_83 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_83 <= _GEN_4963;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_84 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_84 <= _GEN_4964;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_85 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_85 <= _GEN_4965;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_86 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_86 <= _GEN_4966;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_87 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_87 <= _GEN_4967;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_88 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_88 <= _GEN_4968;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_89 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_89 <= _GEN_4969;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_90 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_90 <= _GEN_4970;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_91 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_91 <= _GEN_4971;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_92 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_92 <= _GEN_4972;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_93 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_93 <= _GEN_4973;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_94 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_94 <= _GEN_4974;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_95 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_95 <= _GEN_4975;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_96 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_96 <= _GEN_4976;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_97 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_97 <= _GEN_4977;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_98 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_98 <= _GEN_4978;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_99 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_99 <= _GEN_4979;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_100 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_100 <= _GEN_4980;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_101 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_101 <= _GEN_4981;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_102 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_102 <= _GEN_4982;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_103 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_103 <= _GEN_4983;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_104 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_104 <= _GEN_4984;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_105 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_105 <= _GEN_4985;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_106 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_106 <= _GEN_4986;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_107 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_107 <= _GEN_4987;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_108 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_108 <= _GEN_4988;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_109 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_109 <= _GEN_4989;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_110 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_110 <= _GEN_4990;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_111 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_111 <= _GEN_4991;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_112 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_112 <= _GEN_4992;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_113 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_113 <= _GEN_4993;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_114 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_114 <= _GEN_4994;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_115 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_115 <= _GEN_4995;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_116 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_116 <= _GEN_4996;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_117 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_117 <= _GEN_4997;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_118 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_118 <= _GEN_4998;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_119 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_119 <= _GEN_4999;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_120 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_120 <= _GEN_5000;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_121 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_121 <= _GEN_5001;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_122 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_122 <= _GEN_5002;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_123 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_123 <= _GEN_5003;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_124 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_124 <= _GEN_5004;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_125 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_125 <= _GEN_5005;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_126 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_126 <= _GEN_5006;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_127 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_127 <= _GEN_5007;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_0 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_0 <= _GEN_4623;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_1 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_1 <= _GEN_4624;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_2 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_2 <= _GEN_4625;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_3 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_3 <= _GEN_4626;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_4 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_4 <= _GEN_4627;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_5 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_5 <= _GEN_4628;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_6 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_6 <= _GEN_4629;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_7 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_7 <= _GEN_4630;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_8 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_8 <= _GEN_4631;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_9 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_9 <= _GEN_4632;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_10 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_10 <= _GEN_4633;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_11 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_11 <= _GEN_4634;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_12 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_12 <= _GEN_4635;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_13 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_13 <= _GEN_4636;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_14 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_14 <= _GEN_4637;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_15 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_15 <= _GEN_4638;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_16 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_16 <= _GEN_4639;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_17 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_17 <= _GEN_4640;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_18 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_18 <= _GEN_4641;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_19 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_19 <= _GEN_4642;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_20 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_20 <= _GEN_4643;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_21 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_21 <= _GEN_4644;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_22 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_22 <= _GEN_4645;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_23 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_23 <= _GEN_4646;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_24 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_24 <= _GEN_4647;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_25 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_25 <= _GEN_4648;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_26 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_26 <= _GEN_4649;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_27 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_27 <= _GEN_4650;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_28 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_28 <= _GEN_4651;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_29 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_29 <= _GEN_4652;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_30 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_30 <= _GEN_4653;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_31 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_31 <= _GEN_4654;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_32 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_32 <= _GEN_4655;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_33 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_33 <= _GEN_4656;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_34 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_34 <= _GEN_4657;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_35 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_35 <= _GEN_4658;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_36 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_36 <= _GEN_4659;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_37 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_37 <= _GEN_4660;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_38 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_38 <= _GEN_4661;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_39 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_39 <= _GEN_4662;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_40 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_40 <= _GEN_4663;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_41 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_41 <= _GEN_4664;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_42 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_42 <= _GEN_4665;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_43 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_43 <= _GEN_4666;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_44 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_44 <= _GEN_4667;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_45 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_45 <= _GEN_4668;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_46 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_46 <= _GEN_4669;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_47 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_47 <= _GEN_4670;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_48 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_48 <= _GEN_4671;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_49 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_49 <= _GEN_4672;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_50 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_50 <= _GEN_4673;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_51 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_51 <= _GEN_4674;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_52 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_52 <= _GEN_4675;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_53 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_53 <= _GEN_4676;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_54 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_54 <= _GEN_4677;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_55 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_55 <= _GEN_4678;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_56 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_56 <= _GEN_4679;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_57 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_57 <= _GEN_4680;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_58 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_58 <= _GEN_4681;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_59 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_59 <= _GEN_4682;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_60 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_60 <= _GEN_4683;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_61 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_61 <= _GEN_4684;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_62 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_62 <= _GEN_4685;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_63 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_63 <= _GEN_4686;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_64 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_64 <= _GEN_4687;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_65 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_65 <= _GEN_4688;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_66 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_66 <= _GEN_4689;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_67 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_67 <= _GEN_4690;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_68 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_68 <= _GEN_4691;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_69 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_69 <= _GEN_4692;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_70 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_70 <= _GEN_4693;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_71 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_71 <= _GEN_4694;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_72 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_72 <= _GEN_4695;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_73 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_73 <= _GEN_4696;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_74 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_74 <= _GEN_4697;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_75 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_75 <= _GEN_4698;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_76 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_76 <= _GEN_4699;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_77 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_77 <= _GEN_4700;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_78 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_78 <= _GEN_4701;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_79 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_79 <= _GEN_4702;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_80 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_80 <= _GEN_4703;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_81 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_81 <= _GEN_4704;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_82 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_82 <= _GEN_4705;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_83 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_83 <= _GEN_4706;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_84 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_84 <= _GEN_4707;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_85 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_85 <= _GEN_4708;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_86 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_86 <= _GEN_4709;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_87 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_87 <= _GEN_4710;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_88 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_88 <= _GEN_4711;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_89 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_89 <= _GEN_4712;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_90 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_90 <= _GEN_4713;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_91 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_91 <= _GEN_4714;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_92 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_92 <= _GEN_4715;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_93 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_93 <= _GEN_4716;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_94 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_94 <= _GEN_4717;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_95 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_95 <= _GEN_4718;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_96 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_96 <= _GEN_4719;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_97 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_97 <= _GEN_4720;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_98 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_98 <= _GEN_4721;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_99 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_99 <= _GEN_4722;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_100 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_100 <= _GEN_4723;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_101 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_101 <= _GEN_4724;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_102 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_102 <= _GEN_4725;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_103 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_103 <= _GEN_4726;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_104 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_104 <= _GEN_4727;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_105 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_105 <= _GEN_4728;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_106 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_106 <= _GEN_4729;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_107 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_107 <= _GEN_4730;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_108 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_108 <= _GEN_4731;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_109 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_109 <= _GEN_4732;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_110 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_110 <= _GEN_4733;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_111 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_111 <= _GEN_4734;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_112 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_112 <= _GEN_4735;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_113 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_113 <= _GEN_4736;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_114 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_114 <= _GEN_4737;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_115 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_115 <= _GEN_4738;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_116 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_116 <= _GEN_4739;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_117 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_117 <= _GEN_4740;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_118 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_118 <= _GEN_4741;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_119 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_119 <= _GEN_4742;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_120 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_120 <= _GEN_4743;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_121 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_121 <= _GEN_4744;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_122 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_122 <= _GEN_4745;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_123 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_123 <= _GEN_4746;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_124 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_124 <= _GEN_4747;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_125 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_125 <= _GEN_4748;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_126 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_126 <= _GEN_4749;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_127 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_127 <= _GEN_4750;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_0 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_0 <= _GEN_5008;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_1 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_1 <= _GEN_5009;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_2 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_2 <= _GEN_5010;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_3 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_3 <= _GEN_5011;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_4 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_4 <= _GEN_5012;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_5 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_5 <= _GEN_5013;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_6 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_6 <= _GEN_5014;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_7 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_7 <= _GEN_5015;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_8 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_8 <= _GEN_5016;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_9 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_9 <= _GEN_5017;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_10 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_10 <= _GEN_5018;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_11 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_11 <= _GEN_5019;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_12 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_12 <= _GEN_5020;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_13 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_13 <= _GEN_5021;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_14 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_14 <= _GEN_5022;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_15 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_15 <= _GEN_5023;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_16 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_16 <= _GEN_5024;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_17 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_17 <= _GEN_5025;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_18 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_18 <= _GEN_5026;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_19 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_19 <= _GEN_5027;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_20 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_20 <= _GEN_5028;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_21 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_21 <= _GEN_5029;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_22 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_22 <= _GEN_5030;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_23 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_23 <= _GEN_5031;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_24 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_24 <= _GEN_5032;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_25 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_25 <= _GEN_5033;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_26 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_26 <= _GEN_5034;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_27 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_27 <= _GEN_5035;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_28 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_28 <= _GEN_5036;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_29 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_29 <= _GEN_5037;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_30 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_30 <= _GEN_5038;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_31 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_31 <= _GEN_5039;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_32 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_32 <= _GEN_5040;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_33 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_33 <= _GEN_5041;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_34 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_34 <= _GEN_5042;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_35 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_35 <= _GEN_5043;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_36 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_36 <= _GEN_5044;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_37 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_37 <= _GEN_5045;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_38 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_38 <= _GEN_5046;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_39 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_39 <= _GEN_5047;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_40 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_40 <= _GEN_5048;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_41 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_41 <= _GEN_5049;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_42 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_42 <= _GEN_5050;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_43 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_43 <= _GEN_5051;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_44 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_44 <= _GEN_5052;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_45 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_45 <= _GEN_5053;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_46 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_46 <= _GEN_5054;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_47 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_47 <= _GEN_5055;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_48 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_48 <= _GEN_5056;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_49 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_49 <= _GEN_5057;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_50 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_50 <= _GEN_5058;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_51 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_51 <= _GEN_5059;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_52 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_52 <= _GEN_5060;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_53 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_53 <= _GEN_5061;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_54 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_54 <= _GEN_5062;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_55 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_55 <= _GEN_5063;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_56 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_56 <= _GEN_5064;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_57 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_57 <= _GEN_5065;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_58 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_58 <= _GEN_5066;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_59 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_59 <= _GEN_5067;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_60 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_60 <= _GEN_5068;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_61 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_61 <= _GEN_5069;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_62 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_62 <= _GEN_5070;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_63 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_63 <= _GEN_5071;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_64 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_64 <= _GEN_5072;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_65 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_65 <= _GEN_5073;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_66 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_66 <= _GEN_5074;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_67 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_67 <= _GEN_5075;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_68 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_68 <= _GEN_5076;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_69 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_69 <= _GEN_5077;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_70 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_70 <= _GEN_5078;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_71 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_71 <= _GEN_5079;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_72 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_72 <= _GEN_5080;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_73 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_73 <= _GEN_5081;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_74 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_74 <= _GEN_5082;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_75 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_75 <= _GEN_5083;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_76 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_76 <= _GEN_5084;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_77 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_77 <= _GEN_5085;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_78 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_78 <= _GEN_5086;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_79 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_79 <= _GEN_5087;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_80 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_80 <= _GEN_5088;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_81 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_81 <= _GEN_5089;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_82 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_82 <= _GEN_5090;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_83 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_83 <= _GEN_5091;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_84 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_84 <= _GEN_5092;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_85 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_85 <= _GEN_5093;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_86 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_86 <= _GEN_5094;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_87 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_87 <= _GEN_5095;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_88 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_88 <= _GEN_5096;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_89 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_89 <= _GEN_5097;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_90 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_90 <= _GEN_5098;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_91 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_91 <= _GEN_5099;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_92 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_92 <= _GEN_5100;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_93 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_93 <= _GEN_5101;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_94 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_94 <= _GEN_5102;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_95 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_95 <= _GEN_5103;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_96 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_96 <= _GEN_5104;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_97 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_97 <= _GEN_5105;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_98 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_98 <= _GEN_5106;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_99 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_99 <= _GEN_5107;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_100 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_100 <= _GEN_5108;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_101 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_101 <= _GEN_5109;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_102 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_102 <= _GEN_5110;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_103 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_103 <= _GEN_5111;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_104 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_104 <= _GEN_5112;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_105 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_105 <= _GEN_5113;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_106 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_106 <= _GEN_5114;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_107 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_107 <= _GEN_5115;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_108 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_108 <= _GEN_5116;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_109 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_109 <= _GEN_5117;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_110 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_110 <= _GEN_5118;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_111 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_111 <= _GEN_5119;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_112 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_112 <= _GEN_5120;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_113 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_113 <= _GEN_5121;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_114 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_114 <= _GEN_5122;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_115 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_115 <= _GEN_5123;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_116 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_116 <= _GEN_5124;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_117 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_117 <= _GEN_5125;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_118 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_118 <= _GEN_5126;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_119 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_119 <= _GEN_5127;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_120 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_120 <= _GEN_5128;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_121 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_121 <= _GEN_5129;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_122 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_122 <= _GEN_5130;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_123 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_123 <= _GEN_5131;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_124 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_124 <= _GEN_5132;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_125 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_125 <= _GEN_5133;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_126 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_126 <= _GEN_5134;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_127 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_127 <= _GEN_5135;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:27]
      way0_hit <= 1'h0; // @[i_cache.scala 23:27]
    end else begin
      way0_hit <= _T_2;
    end
    if (reset) begin // @[i_cache.scala 24:27]
      way1_hit <= 1'h0; // @[i_cache.scala 24:27]
    end else begin
      way1_hit <= _T_5;
    end
    if (reset) begin // @[i_cache.scala 26:28]
      unuse_way <= 2'h0; // @[i_cache.scala 26:28]
    end else if (~_GEN_255) begin // @[i_cache.scala 45:31]
      unuse_way <= 2'h1; // @[i_cache.scala 46:19]
    end else if (~_GEN_512) begin // @[i_cache.scala 47:37]
      unuse_way <= 2'h2; // @[i_cache.scala 48:19]
    end else begin
      unuse_way <= 2'h0; // @[i_cache.scala 50:19]
    end
    if (reset) begin // @[i_cache.scala 27:31]
      receive_data <= 64'h0; // @[i_cache.scala 27:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (3'h2 == state) begin // @[i_cache.scala 55:18]
          receive_data <= _GEN_521;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:24]
      quene <= 1'h0; // @[i_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          quene <= _GEN_4751;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 53:24]
      state <= 3'h0; // @[i_cache.scala 53:24]
    end else if (3'h0 == state) begin // @[i_cache.scala 55:18]
      if (io_from_ifu_arvalid) begin // @[i_cache.scala 57:38]
        state <= 3'h1; // @[i_cache.scala 58:23]
      end
    end else if (3'h1 == state) begin // @[i_cache.scala 55:18]
      if (way0_hit) begin // @[i_cache.scala 63:27]
        state <= _GEN_517;
      end else begin
        state <= _GEN_518;
      end
    end else if (3'h2 == state) begin // @[i_cache.scala 55:18]
      state <= _GEN_520;
    end else begin
      state <= _GEN_4366;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ram_0_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ram_0_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ram_0_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ram_0_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ram_0_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ram_0_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ram_0_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ram_0_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  ram_0_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  ram_0_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  ram_0_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  ram_0_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  ram_0_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  ram_0_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  ram_0_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  ram_0_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  ram_0_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  ram_0_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  ram_0_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  ram_0_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  ram_0_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  ram_0_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  ram_0_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  ram_0_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  ram_0_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  ram_0_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  ram_0_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  ram_0_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  ram_0_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  ram_0_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  ram_0_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  ram_0_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  ram_0_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  ram_0_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  ram_0_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  ram_0_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  ram_0_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  ram_0_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  ram_0_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  ram_0_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  ram_0_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  ram_0_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  ram_0_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  ram_0_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  ram_0_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  ram_0_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  ram_0_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  ram_0_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  ram_0_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  ram_0_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  ram_0_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  ram_0_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  ram_0_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  ram_0_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  ram_0_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  ram_0_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  ram_0_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  ram_0_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  ram_0_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  ram_0_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  ram_0_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  ram_0_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  ram_0_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  ram_0_63 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  ram_0_64 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  ram_0_65 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  ram_0_66 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  ram_0_67 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  ram_0_68 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  ram_0_69 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  ram_0_70 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  ram_0_71 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  ram_0_72 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  ram_0_73 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  ram_0_74 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  ram_0_75 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  ram_0_76 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  ram_0_77 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  ram_0_78 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  ram_0_79 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  ram_0_80 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  ram_0_81 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  ram_0_82 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  ram_0_83 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  ram_0_84 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  ram_0_85 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  ram_0_86 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  ram_0_87 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  ram_0_88 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  ram_0_89 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  ram_0_90 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  ram_0_91 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  ram_0_92 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  ram_0_93 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  ram_0_94 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  ram_0_95 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  ram_0_96 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  ram_0_97 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  ram_0_98 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  ram_0_99 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  ram_0_100 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  ram_0_101 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  ram_0_102 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  ram_0_103 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  ram_0_104 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  ram_0_105 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  ram_0_106 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  ram_0_107 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  ram_0_108 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  ram_0_109 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  ram_0_110 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  ram_0_111 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  ram_0_112 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  ram_0_113 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  ram_0_114 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  ram_0_115 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  ram_0_116 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  ram_0_117 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  ram_0_118 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  ram_0_119 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  ram_0_120 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  ram_0_121 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  ram_0_122 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  ram_0_123 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  ram_0_124 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  ram_0_125 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  ram_0_126 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  ram_0_127 = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  ram_1_0 = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  ram_1_1 = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  ram_1_2 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  ram_1_3 = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  ram_1_4 = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  ram_1_5 = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  ram_1_6 = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  ram_1_7 = _RAND_135[63:0];
  _RAND_136 = {2{`RANDOM}};
  ram_1_8 = _RAND_136[63:0];
  _RAND_137 = {2{`RANDOM}};
  ram_1_9 = _RAND_137[63:0];
  _RAND_138 = {2{`RANDOM}};
  ram_1_10 = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  ram_1_11 = _RAND_139[63:0];
  _RAND_140 = {2{`RANDOM}};
  ram_1_12 = _RAND_140[63:0];
  _RAND_141 = {2{`RANDOM}};
  ram_1_13 = _RAND_141[63:0];
  _RAND_142 = {2{`RANDOM}};
  ram_1_14 = _RAND_142[63:0];
  _RAND_143 = {2{`RANDOM}};
  ram_1_15 = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  ram_1_16 = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  ram_1_17 = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  ram_1_18 = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  ram_1_19 = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  ram_1_20 = _RAND_148[63:0];
  _RAND_149 = {2{`RANDOM}};
  ram_1_21 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  ram_1_22 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  ram_1_23 = _RAND_151[63:0];
  _RAND_152 = {2{`RANDOM}};
  ram_1_24 = _RAND_152[63:0];
  _RAND_153 = {2{`RANDOM}};
  ram_1_25 = _RAND_153[63:0];
  _RAND_154 = {2{`RANDOM}};
  ram_1_26 = _RAND_154[63:0];
  _RAND_155 = {2{`RANDOM}};
  ram_1_27 = _RAND_155[63:0];
  _RAND_156 = {2{`RANDOM}};
  ram_1_28 = _RAND_156[63:0];
  _RAND_157 = {2{`RANDOM}};
  ram_1_29 = _RAND_157[63:0];
  _RAND_158 = {2{`RANDOM}};
  ram_1_30 = _RAND_158[63:0];
  _RAND_159 = {2{`RANDOM}};
  ram_1_31 = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  ram_1_32 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  ram_1_33 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  ram_1_34 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  ram_1_35 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  ram_1_36 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  ram_1_37 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  ram_1_38 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  ram_1_39 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  ram_1_40 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  ram_1_41 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  ram_1_42 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  ram_1_43 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  ram_1_44 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  ram_1_45 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  ram_1_46 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  ram_1_47 = _RAND_175[63:0];
  _RAND_176 = {2{`RANDOM}};
  ram_1_48 = _RAND_176[63:0];
  _RAND_177 = {2{`RANDOM}};
  ram_1_49 = _RAND_177[63:0];
  _RAND_178 = {2{`RANDOM}};
  ram_1_50 = _RAND_178[63:0];
  _RAND_179 = {2{`RANDOM}};
  ram_1_51 = _RAND_179[63:0];
  _RAND_180 = {2{`RANDOM}};
  ram_1_52 = _RAND_180[63:0];
  _RAND_181 = {2{`RANDOM}};
  ram_1_53 = _RAND_181[63:0];
  _RAND_182 = {2{`RANDOM}};
  ram_1_54 = _RAND_182[63:0];
  _RAND_183 = {2{`RANDOM}};
  ram_1_55 = _RAND_183[63:0];
  _RAND_184 = {2{`RANDOM}};
  ram_1_56 = _RAND_184[63:0];
  _RAND_185 = {2{`RANDOM}};
  ram_1_57 = _RAND_185[63:0];
  _RAND_186 = {2{`RANDOM}};
  ram_1_58 = _RAND_186[63:0];
  _RAND_187 = {2{`RANDOM}};
  ram_1_59 = _RAND_187[63:0];
  _RAND_188 = {2{`RANDOM}};
  ram_1_60 = _RAND_188[63:0];
  _RAND_189 = {2{`RANDOM}};
  ram_1_61 = _RAND_189[63:0];
  _RAND_190 = {2{`RANDOM}};
  ram_1_62 = _RAND_190[63:0];
  _RAND_191 = {2{`RANDOM}};
  ram_1_63 = _RAND_191[63:0];
  _RAND_192 = {2{`RANDOM}};
  ram_1_64 = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  ram_1_65 = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  ram_1_66 = _RAND_194[63:0];
  _RAND_195 = {2{`RANDOM}};
  ram_1_67 = _RAND_195[63:0];
  _RAND_196 = {2{`RANDOM}};
  ram_1_68 = _RAND_196[63:0];
  _RAND_197 = {2{`RANDOM}};
  ram_1_69 = _RAND_197[63:0];
  _RAND_198 = {2{`RANDOM}};
  ram_1_70 = _RAND_198[63:0];
  _RAND_199 = {2{`RANDOM}};
  ram_1_71 = _RAND_199[63:0];
  _RAND_200 = {2{`RANDOM}};
  ram_1_72 = _RAND_200[63:0];
  _RAND_201 = {2{`RANDOM}};
  ram_1_73 = _RAND_201[63:0];
  _RAND_202 = {2{`RANDOM}};
  ram_1_74 = _RAND_202[63:0];
  _RAND_203 = {2{`RANDOM}};
  ram_1_75 = _RAND_203[63:0];
  _RAND_204 = {2{`RANDOM}};
  ram_1_76 = _RAND_204[63:0];
  _RAND_205 = {2{`RANDOM}};
  ram_1_77 = _RAND_205[63:0];
  _RAND_206 = {2{`RANDOM}};
  ram_1_78 = _RAND_206[63:0];
  _RAND_207 = {2{`RANDOM}};
  ram_1_79 = _RAND_207[63:0];
  _RAND_208 = {2{`RANDOM}};
  ram_1_80 = _RAND_208[63:0];
  _RAND_209 = {2{`RANDOM}};
  ram_1_81 = _RAND_209[63:0];
  _RAND_210 = {2{`RANDOM}};
  ram_1_82 = _RAND_210[63:0];
  _RAND_211 = {2{`RANDOM}};
  ram_1_83 = _RAND_211[63:0];
  _RAND_212 = {2{`RANDOM}};
  ram_1_84 = _RAND_212[63:0];
  _RAND_213 = {2{`RANDOM}};
  ram_1_85 = _RAND_213[63:0];
  _RAND_214 = {2{`RANDOM}};
  ram_1_86 = _RAND_214[63:0];
  _RAND_215 = {2{`RANDOM}};
  ram_1_87 = _RAND_215[63:0];
  _RAND_216 = {2{`RANDOM}};
  ram_1_88 = _RAND_216[63:0];
  _RAND_217 = {2{`RANDOM}};
  ram_1_89 = _RAND_217[63:0];
  _RAND_218 = {2{`RANDOM}};
  ram_1_90 = _RAND_218[63:0];
  _RAND_219 = {2{`RANDOM}};
  ram_1_91 = _RAND_219[63:0];
  _RAND_220 = {2{`RANDOM}};
  ram_1_92 = _RAND_220[63:0];
  _RAND_221 = {2{`RANDOM}};
  ram_1_93 = _RAND_221[63:0];
  _RAND_222 = {2{`RANDOM}};
  ram_1_94 = _RAND_222[63:0];
  _RAND_223 = {2{`RANDOM}};
  ram_1_95 = _RAND_223[63:0];
  _RAND_224 = {2{`RANDOM}};
  ram_1_96 = _RAND_224[63:0];
  _RAND_225 = {2{`RANDOM}};
  ram_1_97 = _RAND_225[63:0];
  _RAND_226 = {2{`RANDOM}};
  ram_1_98 = _RAND_226[63:0];
  _RAND_227 = {2{`RANDOM}};
  ram_1_99 = _RAND_227[63:0];
  _RAND_228 = {2{`RANDOM}};
  ram_1_100 = _RAND_228[63:0];
  _RAND_229 = {2{`RANDOM}};
  ram_1_101 = _RAND_229[63:0];
  _RAND_230 = {2{`RANDOM}};
  ram_1_102 = _RAND_230[63:0];
  _RAND_231 = {2{`RANDOM}};
  ram_1_103 = _RAND_231[63:0];
  _RAND_232 = {2{`RANDOM}};
  ram_1_104 = _RAND_232[63:0];
  _RAND_233 = {2{`RANDOM}};
  ram_1_105 = _RAND_233[63:0];
  _RAND_234 = {2{`RANDOM}};
  ram_1_106 = _RAND_234[63:0];
  _RAND_235 = {2{`RANDOM}};
  ram_1_107 = _RAND_235[63:0];
  _RAND_236 = {2{`RANDOM}};
  ram_1_108 = _RAND_236[63:0];
  _RAND_237 = {2{`RANDOM}};
  ram_1_109 = _RAND_237[63:0];
  _RAND_238 = {2{`RANDOM}};
  ram_1_110 = _RAND_238[63:0];
  _RAND_239 = {2{`RANDOM}};
  ram_1_111 = _RAND_239[63:0];
  _RAND_240 = {2{`RANDOM}};
  ram_1_112 = _RAND_240[63:0];
  _RAND_241 = {2{`RANDOM}};
  ram_1_113 = _RAND_241[63:0];
  _RAND_242 = {2{`RANDOM}};
  ram_1_114 = _RAND_242[63:0];
  _RAND_243 = {2{`RANDOM}};
  ram_1_115 = _RAND_243[63:0];
  _RAND_244 = {2{`RANDOM}};
  ram_1_116 = _RAND_244[63:0];
  _RAND_245 = {2{`RANDOM}};
  ram_1_117 = _RAND_245[63:0];
  _RAND_246 = {2{`RANDOM}};
  ram_1_118 = _RAND_246[63:0];
  _RAND_247 = {2{`RANDOM}};
  ram_1_119 = _RAND_247[63:0];
  _RAND_248 = {2{`RANDOM}};
  ram_1_120 = _RAND_248[63:0];
  _RAND_249 = {2{`RANDOM}};
  ram_1_121 = _RAND_249[63:0];
  _RAND_250 = {2{`RANDOM}};
  ram_1_122 = _RAND_250[63:0];
  _RAND_251 = {2{`RANDOM}};
  ram_1_123 = _RAND_251[63:0];
  _RAND_252 = {2{`RANDOM}};
  ram_1_124 = _RAND_252[63:0];
  _RAND_253 = {2{`RANDOM}};
  ram_1_125 = _RAND_253[63:0];
  _RAND_254 = {2{`RANDOM}};
  ram_1_126 = _RAND_254[63:0];
  _RAND_255 = {2{`RANDOM}};
  ram_1_127 = _RAND_255[63:0];
  _RAND_256 = {1{`RANDOM}};
  tag_0_0 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  tag_0_1 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  tag_0_2 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  tag_0_3 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  tag_0_4 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  tag_0_5 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  tag_0_6 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  tag_0_7 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  tag_0_8 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  tag_0_9 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  tag_0_10 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  tag_0_11 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  tag_0_12 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  tag_0_13 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  tag_0_14 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  tag_0_15 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  tag_0_16 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  tag_0_17 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  tag_0_18 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  tag_0_19 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  tag_0_20 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  tag_0_21 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  tag_0_22 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  tag_0_23 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  tag_0_24 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  tag_0_25 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  tag_0_26 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  tag_0_27 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  tag_0_28 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  tag_0_29 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  tag_0_30 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  tag_0_31 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  tag_0_32 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  tag_0_33 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  tag_0_34 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  tag_0_35 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  tag_0_36 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  tag_0_37 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  tag_0_38 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  tag_0_39 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  tag_0_40 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  tag_0_41 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  tag_0_42 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  tag_0_43 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  tag_0_44 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  tag_0_45 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  tag_0_46 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  tag_0_47 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  tag_0_48 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  tag_0_49 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  tag_0_50 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  tag_0_51 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  tag_0_52 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  tag_0_53 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  tag_0_54 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  tag_0_55 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  tag_0_56 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  tag_0_57 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  tag_0_58 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  tag_0_59 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  tag_0_60 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  tag_0_61 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  tag_0_62 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  tag_0_63 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  tag_0_64 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  tag_0_65 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  tag_0_66 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  tag_0_67 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  tag_0_68 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  tag_0_69 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  tag_0_70 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  tag_0_71 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  tag_0_72 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  tag_0_73 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  tag_0_74 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  tag_0_75 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  tag_0_76 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  tag_0_77 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  tag_0_78 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  tag_0_79 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  tag_0_80 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  tag_0_81 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  tag_0_82 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  tag_0_83 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  tag_0_84 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  tag_0_85 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  tag_0_86 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  tag_0_87 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  tag_0_88 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  tag_0_89 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  tag_0_90 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  tag_0_91 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  tag_0_92 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  tag_0_93 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  tag_0_94 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  tag_0_95 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  tag_0_96 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  tag_0_97 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  tag_0_98 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  tag_0_99 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  tag_0_100 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  tag_0_101 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  tag_0_102 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  tag_0_103 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  tag_0_104 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  tag_0_105 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  tag_0_106 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  tag_0_107 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  tag_0_108 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  tag_0_109 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  tag_0_110 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  tag_0_111 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  tag_0_112 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  tag_0_113 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  tag_0_114 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  tag_0_115 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  tag_0_116 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  tag_0_117 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  tag_0_118 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  tag_0_119 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  tag_0_120 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  tag_0_121 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  tag_0_122 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  tag_0_123 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  tag_0_124 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  tag_0_125 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  tag_0_126 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  tag_0_127 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  tag_1_0 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  tag_1_1 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  tag_1_2 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  tag_1_3 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  tag_1_4 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  tag_1_5 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  tag_1_6 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  tag_1_7 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  tag_1_8 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  tag_1_9 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  tag_1_10 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  tag_1_11 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  tag_1_12 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  tag_1_13 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  tag_1_14 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  tag_1_15 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  tag_1_16 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  tag_1_17 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  tag_1_18 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  tag_1_19 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  tag_1_20 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  tag_1_21 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  tag_1_22 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  tag_1_23 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  tag_1_24 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  tag_1_25 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  tag_1_26 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  tag_1_27 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  tag_1_28 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  tag_1_29 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  tag_1_30 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  tag_1_31 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  tag_1_32 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  tag_1_33 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  tag_1_34 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  tag_1_35 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  tag_1_36 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  tag_1_37 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  tag_1_38 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  tag_1_39 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  tag_1_40 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  tag_1_41 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  tag_1_42 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  tag_1_43 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  tag_1_44 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  tag_1_45 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  tag_1_46 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  tag_1_47 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  tag_1_48 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  tag_1_49 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  tag_1_50 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  tag_1_51 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  tag_1_52 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  tag_1_53 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  tag_1_54 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  tag_1_55 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  tag_1_56 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  tag_1_57 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  tag_1_58 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  tag_1_59 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  tag_1_60 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  tag_1_61 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  tag_1_62 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  tag_1_63 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  tag_1_64 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  tag_1_65 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  tag_1_66 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  tag_1_67 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  tag_1_68 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  tag_1_69 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  tag_1_70 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  tag_1_71 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  tag_1_72 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  tag_1_73 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  tag_1_74 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  tag_1_75 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  tag_1_76 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  tag_1_77 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  tag_1_78 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  tag_1_79 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  tag_1_80 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  tag_1_81 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  tag_1_82 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  tag_1_83 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  tag_1_84 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  tag_1_85 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  tag_1_86 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  tag_1_87 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  tag_1_88 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  tag_1_89 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  tag_1_90 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  tag_1_91 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  tag_1_92 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  tag_1_93 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  tag_1_94 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  tag_1_95 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  tag_1_96 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  tag_1_97 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  tag_1_98 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  tag_1_99 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  tag_1_100 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  tag_1_101 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  tag_1_102 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  tag_1_103 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  tag_1_104 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  tag_1_105 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  tag_1_106 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  tag_1_107 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  tag_1_108 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  tag_1_109 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  tag_1_110 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  tag_1_111 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  tag_1_112 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  tag_1_113 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  tag_1_114 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  tag_1_115 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  tag_1_116 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  tag_1_117 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  tag_1_118 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  tag_1_119 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  tag_1_120 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  tag_1_121 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  tag_1_122 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  tag_1_123 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  tag_1_124 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  tag_1_125 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  tag_1_126 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  tag_1_127 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  valid_0_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid_0_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  valid_0_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  valid_0_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  valid_0_4 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  valid_0_5 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  valid_0_6 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  valid_0_7 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  valid_0_8 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  valid_0_9 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  valid_0_10 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  valid_0_11 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  valid_0_12 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  valid_0_13 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  valid_0_14 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  valid_0_15 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  valid_0_16 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  valid_0_17 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  valid_0_18 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  valid_0_19 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  valid_0_20 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  valid_0_21 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  valid_0_22 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  valid_0_23 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  valid_0_24 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  valid_0_25 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  valid_0_26 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  valid_0_27 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  valid_0_28 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  valid_0_29 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  valid_0_30 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  valid_0_31 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  valid_0_32 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  valid_0_33 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  valid_0_34 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  valid_0_35 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  valid_0_36 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  valid_0_37 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  valid_0_38 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  valid_0_39 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  valid_0_40 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  valid_0_41 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  valid_0_42 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  valid_0_43 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  valid_0_44 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  valid_0_45 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  valid_0_46 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  valid_0_47 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  valid_0_48 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  valid_0_49 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  valid_0_50 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  valid_0_51 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  valid_0_52 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  valid_0_53 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  valid_0_54 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  valid_0_55 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  valid_0_56 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  valid_0_57 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  valid_0_58 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  valid_0_59 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  valid_0_60 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  valid_0_61 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  valid_0_62 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  valid_0_63 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  valid_0_64 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  valid_0_65 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  valid_0_66 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  valid_0_67 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  valid_0_68 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  valid_0_69 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  valid_0_70 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  valid_0_71 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  valid_0_72 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  valid_0_73 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  valid_0_74 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  valid_0_75 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  valid_0_76 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  valid_0_77 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  valid_0_78 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  valid_0_79 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  valid_0_80 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  valid_0_81 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  valid_0_82 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  valid_0_83 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  valid_0_84 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  valid_0_85 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  valid_0_86 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  valid_0_87 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  valid_0_88 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  valid_0_89 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  valid_0_90 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  valid_0_91 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  valid_0_92 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  valid_0_93 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  valid_0_94 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  valid_0_95 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  valid_0_96 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  valid_0_97 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  valid_0_98 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  valid_0_99 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  valid_0_100 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  valid_0_101 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  valid_0_102 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  valid_0_103 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  valid_0_104 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  valid_0_105 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  valid_0_106 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  valid_0_107 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  valid_0_108 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  valid_0_109 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  valid_0_110 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  valid_0_111 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  valid_0_112 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  valid_0_113 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  valid_0_114 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  valid_0_115 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  valid_0_116 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  valid_0_117 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  valid_0_118 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  valid_0_119 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  valid_0_120 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  valid_0_121 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  valid_0_122 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  valid_0_123 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  valid_0_124 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  valid_0_125 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  valid_0_126 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  valid_0_127 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  valid_1_0 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  valid_1_1 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  valid_1_2 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  valid_1_3 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  valid_1_4 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  valid_1_5 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  valid_1_6 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  valid_1_7 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  valid_1_8 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  valid_1_9 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  valid_1_10 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  valid_1_11 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  valid_1_12 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  valid_1_13 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  valid_1_14 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  valid_1_15 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  valid_1_16 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  valid_1_17 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  valid_1_18 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  valid_1_19 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  valid_1_20 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  valid_1_21 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  valid_1_22 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  valid_1_23 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  valid_1_24 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  valid_1_25 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  valid_1_26 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  valid_1_27 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  valid_1_28 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  valid_1_29 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  valid_1_30 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  valid_1_31 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  valid_1_32 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  valid_1_33 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  valid_1_34 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  valid_1_35 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  valid_1_36 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  valid_1_37 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  valid_1_38 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  valid_1_39 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  valid_1_40 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  valid_1_41 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  valid_1_42 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  valid_1_43 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  valid_1_44 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  valid_1_45 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  valid_1_46 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  valid_1_47 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  valid_1_48 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  valid_1_49 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  valid_1_50 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  valid_1_51 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  valid_1_52 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  valid_1_53 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  valid_1_54 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  valid_1_55 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  valid_1_56 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  valid_1_57 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  valid_1_58 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  valid_1_59 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  valid_1_60 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  valid_1_61 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  valid_1_62 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  valid_1_63 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  valid_1_64 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  valid_1_65 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  valid_1_66 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  valid_1_67 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  valid_1_68 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  valid_1_69 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  valid_1_70 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  valid_1_71 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  valid_1_72 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  valid_1_73 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  valid_1_74 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  valid_1_75 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  valid_1_76 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  valid_1_77 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  valid_1_78 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  valid_1_79 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  valid_1_80 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  valid_1_81 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  valid_1_82 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  valid_1_83 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  valid_1_84 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  valid_1_85 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  valid_1_86 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  valid_1_87 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  valid_1_88 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  valid_1_89 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  valid_1_90 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  valid_1_91 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  valid_1_92 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  valid_1_93 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  valid_1_94 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  valid_1_95 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  valid_1_96 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  valid_1_97 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  valid_1_98 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  valid_1_99 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  valid_1_100 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  valid_1_101 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  valid_1_102 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  valid_1_103 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  valid_1_104 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  valid_1_105 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  valid_1_106 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  valid_1_107 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  valid_1_108 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  valid_1_109 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  valid_1_110 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  valid_1_111 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  valid_1_112 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  valid_1_113 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  valid_1_114 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  valid_1_115 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  valid_1_116 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  valid_1_117 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  valid_1_118 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  valid_1_119 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  valid_1_120 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  valid_1_121 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  valid_1_122 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  valid_1_123 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  valid_1_124 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  valid_1_125 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  valid_1_126 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  valid_1_127 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  way0_hit = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  way1_hit = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  unuse_way = _RAND_770[1:0];
  _RAND_771 = {2{`RANDOM}};
  receive_data = _RAND_771[63:0];
  _RAND_772 = {1{`RANDOM}};
  quene = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  state = _RAND_773[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module D_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_lsu_araddr,
  input         io_from_lsu_arvalid,
  input         io_from_lsu_rready,
  input  [31:0] io_from_lsu_awaddr,
  input         io_from_lsu_awvalid,
  input  [31:0] io_from_lsu_wdata,
  input  [7:0]  io_from_lsu_wstrb,
  input         io_from_lsu_wvalid,
  input         io_from_lsu_bready,
  output        io_to_lsu_arready,
  output [63:0] io_to_lsu_rdata,
  output        io_to_lsu_rvalid,
  output        io_to_lsu_awready,
  output        io_to_lsu_wready,
  output        io_to_lsu_bvalid,
  output [31:0] io_to_axi_araddr,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  output [31:0] io_to_axi_awaddr,
  output        io_to_axi_awvalid,
  output [31:0] io_to_axi_wdata,
  output [7:0]  io_to_axi_wstrb,
  output        io_to_axi_wvalid,
  output        io_to_axi_bready,
  input         io_from_axi_arready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rvalid,
  input         io_from_axi_awready,
  input         io_from_axi_wready,
  input         io_from_axi_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [63:0] _RAND_256;
  reg [63:0] _RAND_257;
  reg [63:0] _RAND_258;
  reg [63:0] _RAND_259;
  reg [63:0] _RAND_260;
  reg [63:0] _RAND_261;
  reg [63:0] _RAND_262;
  reg [63:0] _RAND_263;
  reg [63:0] _RAND_264;
  reg [63:0] _RAND_265;
  reg [63:0] _RAND_266;
  reg [63:0] _RAND_267;
  reg [63:0] _RAND_268;
  reg [63:0] _RAND_269;
  reg [63:0] _RAND_270;
  reg [63:0] _RAND_271;
  reg [63:0] _RAND_272;
  reg [63:0] _RAND_273;
  reg [63:0] _RAND_274;
  reg [63:0] _RAND_275;
  reg [63:0] _RAND_276;
  reg [63:0] _RAND_277;
  reg [63:0] _RAND_278;
  reg [63:0] _RAND_279;
  reg [63:0] _RAND_280;
  reg [63:0] _RAND_281;
  reg [63:0] _RAND_282;
  reg [63:0] _RAND_283;
  reg [63:0] _RAND_284;
  reg [63:0] _RAND_285;
  reg [63:0] _RAND_286;
  reg [63:0] _RAND_287;
  reg [63:0] _RAND_288;
  reg [63:0] _RAND_289;
  reg [63:0] _RAND_290;
  reg [63:0] _RAND_291;
  reg [63:0] _RAND_292;
  reg [63:0] _RAND_293;
  reg [63:0] _RAND_294;
  reg [63:0] _RAND_295;
  reg [63:0] _RAND_296;
  reg [63:0] _RAND_297;
  reg [63:0] _RAND_298;
  reg [63:0] _RAND_299;
  reg [63:0] _RAND_300;
  reg [63:0] _RAND_301;
  reg [63:0] _RAND_302;
  reg [63:0] _RAND_303;
  reg [63:0] _RAND_304;
  reg [63:0] _RAND_305;
  reg [63:0] _RAND_306;
  reg [63:0] _RAND_307;
  reg [63:0] _RAND_308;
  reg [63:0] _RAND_309;
  reg [63:0] _RAND_310;
  reg [63:0] _RAND_311;
  reg [63:0] _RAND_312;
  reg [63:0] _RAND_313;
  reg [63:0] _RAND_314;
  reg [63:0] _RAND_315;
  reg [63:0] _RAND_316;
  reg [63:0] _RAND_317;
  reg [63:0] _RAND_318;
  reg [63:0] _RAND_319;
  reg [63:0] _RAND_320;
  reg [63:0] _RAND_321;
  reg [63:0] _RAND_322;
  reg [63:0] _RAND_323;
  reg [63:0] _RAND_324;
  reg [63:0] _RAND_325;
  reg [63:0] _RAND_326;
  reg [63:0] _RAND_327;
  reg [63:0] _RAND_328;
  reg [63:0] _RAND_329;
  reg [63:0] _RAND_330;
  reg [63:0] _RAND_331;
  reg [63:0] _RAND_332;
  reg [63:0] _RAND_333;
  reg [63:0] _RAND_334;
  reg [63:0] _RAND_335;
  reg [63:0] _RAND_336;
  reg [63:0] _RAND_337;
  reg [63:0] _RAND_338;
  reg [63:0] _RAND_339;
  reg [63:0] _RAND_340;
  reg [63:0] _RAND_341;
  reg [63:0] _RAND_342;
  reg [63:0] _RAND_343;
  reg [63:0] _RAND_344;
  reg [63:0] _RAND_345;
  reg [63:0] _RAND_346;
  reg [63:0] _RAND_347;
  reg [63:0] _RAND_348;
  reg [63:0] _RAND_349;
  reg [63:0] _RAND_350;
  reg [63:0] _RAND_351;
  reg [63:0] _RAND_352;
  reg [63:0] _RAND_353;
  reg [63:0] _RAND_354;
  reg [63:0] _RAND_355;
  reg [63:0] _RAND_356;
  reg [63:0] _RAND_357;
  reg [63:0] _RAND_358;
  reg [63:0] _RAND_359;
  reg [63:0] _RAND_360;
  reg [63:0] _RAND_361;
  reg [63:0] _RAND_362;
  reg [63:0] _RAND_363;
  reg [63:0] _RAND_364;
  reg [63:0] _RAND_365;
  reg [63:0] _RAND_366;
  reg [63:0] _RAND_367;
  reg [63:0] _RAND_368;
  reg [63:0] _RAND_369;
  reg [63:0] _RAND_370;
  reg [63:0] _RAND_371;
  reg [63:0] _RAND_372;
  reg [63:0] _RAND_373;
  reg [63:0] _RAND_374;
  reg [63:0] _RAND_375;
  reg [63:0] _RAND_376;
  reg [63:0] _RAND_377;
  reg [63:0] _RAND_378;
  reg [63:0] _RAND_379;
  reg [63:0] _RAND_380;
  reg [63:0] _RAND_381;
  reg [63:0] _RAND_382;
  reg [63:0] _RAND_383;
  reg [63:0] _RAND_384;
  reg [63:0] _RAND_385;
  reg [63:0] _RAND_386;
  reg [63:0] _RAND_387;
  reg [63:0] _RAND_388;
  reg [63:0] _RAND_389;
  reg [63:0] _RAND_390;
  reg [63:0] _RAND_391;
  reg [63:0] _RAND_392;
  reg [63:0] _RAND_393;
  reg [63:0] _RAND_394;
  reg [63:0] _RAND_395;
  reg [63:0] _RAND_396;
  reg [63:0] _RAND_397;
  reg [63:0] _RAND_398;
  reg [63:0] _RAND_399;
  reg [63:0] _RAND_400;
  reg [63:0] _RAND_401;
  reg [63:0] _RAND_402;
  reg [63:0] _RAND_403;
  reg [63:0] _RAND_404;
  reg [63:0] _RAND_405;
  reg [63:0] _RAND_406;
  reg [63:0] _RAND_407;
  reg [63:0] _RAND_408;
  reg [63:0] _RAND_409;
  reg [63:0] _RAND_410;
  reg [63:0] _RAND_411;
  reg [63:0] _RAND_412;
  reg [63:0] _RAND_413;
  reg [63:0] _RAND_414;
  reg [63:0] _RAND_415;
  reg [63:0] _RAND_416;
  reg [63:0] _RAND_417;
  reg [63:0] _RAND_418;
  reg [63:0] _RAND_419;
  reg [63:0] _RAND_420;
  reg [63:0] _RAND_421;
  reg [63:0] _RAND_422;
  reg [63:0] _RAND_423;
  reg [63:0] _RAND_424;
  reg [63:0] _RAND_425;
  reg [63:0] _RAND_426;
  reg [63:0] _RAND_427;
  reg [63:0] _RAND_428;
  reg [63:0] _RAND_429;
  reg [63:0] _RAND_430;
  reg [63:0] _RAND_431;
  reg [63:0] _RAND_432;
  reg [63:0] _RAND_433;
  reg [63:0] _RAND_434;
  reg [63:0] _RAND_435;
  reg [63:0] _RAND_436;
  reg [63:0] _RAND_437;
  reg [63:0] _RAND_438;
  reg [63:0] _RAND_439;
  reg [63:0] _RAND_440;
  reg [63:0] _RAND_441;
  reg [63:0] _RAND_442;
  reg [63:0] _RAND_443;
  reg [63:0] _RAND_444;
  reg [63:0] _RAND_445;
  reg [63:0] _RAND_446;
  reg [63:0] _RAND_447;
  reg [63:0] _RAND_448;
  reg [63:0] _RAND_449;
  reg [63:0] _RAND_450;
  reg [63:0] _RAND_451;
  reg [63:0] _RAND_452;
  reg [63:0] _RAND_453;
  reg [63:0] _RAND_454;
  reg [63:0] _RAND_455;
  reg [63:0] _RAND_456;
  reg [63:0] _RAND_457;
  reg [63:0] _RAND_458;
  reg [63:0] _RAND_459;
  reg [63:0] _RAND_460;
  reg [63:0] _RAND_461;
  reg [63:0] _RAND_462;
  reg [63:0] _RAND_463;
  reg [63:0] _RAND_464;
  reg [63:0] _RAND_465;
  reg [63:0] _RAND_466;
  reg [63:0] _RAND_467;
  reg [63:0] _RAND_468;
  reg [63:0] _RAND_469;
  reg [63:0] _RAND_470;
  reg [63:0] _RAND_471;
  reg [63:0] _RAND_472;
  reg [63:0] _RAND_473;
  reg [63:0] _RAND_474;
  reg [63:0] _RAND_475;
  reg [63:0] _RAND_476;
  reg [63:0] _RAND_477;
  reg [63:0] _RAND_478;
  reg [63:0] _RAND_479;
  reg [63:0] _RAND_480;
  reg [63:0] _RAND_481;
  reg [63:0] _RAND_482;
  reg [63:0] _RAND_483;
  reg [63:0] _RAND_484;
  reg [63:0] _RAND_485;
  reg [63:0] _RAND_486;
  reg [63:0] _RAND_487;
  reg [63:0] _RAND_488;
  reg [63:0] _RAND_489;
  reg [63:0] _RAND_490;
  reg [63:0] _RAND_491;
  reg [63:0] _RAND_492;
  reg [63:0] _RAND_493;
  reg [63:0] _RAND_494;
  reg [63:0] _RAND_495;
  reg [63:0] _RAND_496;
  reg [63:0] _RAND_497;
  reg [63:0] _RAND_498;
  reg [63:0] _RAND_499;
  reg [63:0] _RAND_500;
  reg [63:0] _RAND_501;
  reg [63:0] _RAND_502;
  reg [63:0] _RAND_503;
  reg [63:0] _RAND_504;
  reg [63:0] _RAND_505;
  reg [63:0] _RAND_506;
  reg [63:0] _RAND_507;
  reg [63:0] _RAND_508;
  reg [63:0] _RAND_509;
  reg [63:0] _RAND_510;
  reg [63:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [63:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [63:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = ~reset; // @[d_cache.scala 15:11]
  reg [63:0] ram_0_0; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_1; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_2; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_3; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_4; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_5; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_6; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_7; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_8; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_9; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_10; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_11; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_12; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_13; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_14; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_15; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_16; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_17; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_18; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_19; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_20; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_21; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_22; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_23; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_24; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_25; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_26; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_27; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_28; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_29; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_30; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_31; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_32; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_33; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_34; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_35; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_36; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_37; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_38; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_39; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_40; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_41; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_42; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_43; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_44; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_45; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_46; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_47; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_48; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_49; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_50; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_51; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_52; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_53; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_54; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_55; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_56; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_57; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_58; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_59; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_60; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_61; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_62; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_63; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_64; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_65; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_66; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_67; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_68; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_69; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_70; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_71; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_72; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_73; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_74; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_75; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_76; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_77; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_78; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_79; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_80; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_81; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_82; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_83; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_84; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_85; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_86; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_87; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_88; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_89; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_90; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_91; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_92; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_93; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_94; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_95; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_96; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_97; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_98; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_99; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_100; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_101; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_102; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_103; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_104; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_105; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_106; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_107; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_108; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_109; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_110; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_111; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_112; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_113; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_114; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_115; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_116; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_117; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_118; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_119; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_120; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_121; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_122; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_123; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_124; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_125; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_126; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_127; // @[d_cache.scala 18:24]
  reg [63:0] ram_1_0; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_1; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_2; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_3; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_4; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_5; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_6; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_7; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_8; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_9; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_10; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_11; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_12; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_13; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_14; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_15; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_16; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_17; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_18; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_19; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_20; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_21; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_22; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_23; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_24; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_25; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_26; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_27; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_28; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_29; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_30; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_31; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_32; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_33; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_34; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_35; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_36; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_37; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_38; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_39; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_40; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_41; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_42; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_43; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_44; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_45; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_46; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_47; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_48; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_49; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_50; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_51; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_52; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_53; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_54; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_55; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_56; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_57; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_58; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_59; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_60; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_61; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_62; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_63; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_64; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_65; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_66; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_67; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_68; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_69; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_70; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_71; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_72; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_73; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_74; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_75; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_76; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_77; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_78; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_79; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_80; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_81; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_82; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_83; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_84; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_85; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_86; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_87; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_88; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_89; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_90; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_91; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_92; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_93; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_94; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_95; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_96; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_97; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_98; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_99; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_100; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_101; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_102; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_103; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_104; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_105; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_106; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_107; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_108; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_109; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_110; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_111; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_112; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_113; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_114; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_115; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_116; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_117; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_118; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_119; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_120; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_121; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_122; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_123; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_124; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_125; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_126; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_127; // @[d_cache.scala 19:24]
  reg [63:0] recent_wdata0_0; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_1; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_2; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_3; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_4; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_5; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_6; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_7; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_8; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_9; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_10; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_11; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_12; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_13; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_14; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_15; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_16; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_17; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_18; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_19; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_20; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_21; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_22; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_23; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_24; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_25; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_26; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_27; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_28; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_29; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_30; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_31; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_32; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_33; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_34; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_35; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_36; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_37; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_38; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_39; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_40; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_41; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_42; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_43; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_44; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_45; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_46; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_47; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_48; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_49; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_50; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_51; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_52; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_53; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_54; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_55; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_56; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_57; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_58; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_59; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_60; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_61; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_62; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_63; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_64; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_65; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_66; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_67; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_68; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_69; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_70; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_71; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_72; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_73; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_74; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_75; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_76; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_77; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_78; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_79; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_80; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_81; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_82; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_83; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_84; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_85; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_86; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_87; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_88; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_89; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_90; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_91; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_92; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_93; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_94; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_95; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_96; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_97; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_98; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_99; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_100; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_101; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_102; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_103; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_104; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_105; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_106; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_107; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_108; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_109; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_110; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_111; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_112; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_113; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_114; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_115; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_116; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_117; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_118; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_119; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_120; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_121; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_122; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_123; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_124; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_125; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_126; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata0_127; // @[d_cache.scala 20:32]
  reg [63:0] recent_wdata1_0; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_1; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_2; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_3; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_4; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_5; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_6; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_7; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_8; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_9; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_10; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_11; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_12; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_13; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_14; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_15; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_16; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_17; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_18; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_19; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_20; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_21; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_22; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_23; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_24; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_25; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_26; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_27; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_28; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_29; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_30; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_31; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_32; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_33; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_34; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_35; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_36; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_37; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_38; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_39; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_40; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_41; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_42; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_43; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_44; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_45; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_46; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_47; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_48; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_49; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_50; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_51; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_52; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_53; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_54; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_55; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_56; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_57; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_58; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_59; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_60; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_61; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_62; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_63; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_64; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_65; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_66; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_67; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_68; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_69; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_70; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_71; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_72; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_73; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_74; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_75; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_76; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_77; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_78; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_79; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_80; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_81; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_82; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_83; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_84; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_85; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_86; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_87; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_88; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_89; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_90; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_91; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_92; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_93; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_94; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_95; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_96; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_97; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_98; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_99; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_100; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_101; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_102; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_103; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_104; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_105; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_106; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_107; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_108; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_109; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_110; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_111; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_112; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_113; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_114; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_115; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_116; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_117; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_118; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_119; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_120; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_121; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_122; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_123; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_124; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_125; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_126; // @[d_cache.scala 21:32]
  reg [63:0] recent_wdata1_127; // @[d_cache.scala 21:32]
  reg [31:0] tag_0_0; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_1; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_2; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_3; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_4; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_5; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_6; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_7; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_8; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_9; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_10; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_11; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_12; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_13; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_14; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_15; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_16; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_17; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_18; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_19; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_20; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_21; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_22; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_23; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_24; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_25; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_26; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_27; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_28; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_29; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_30; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_31; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_32; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_33; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_34; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_35; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_36; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_37; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_38; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_39; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_40; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_41; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_42; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_43; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_44; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_45; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_46; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_47; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_48; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_49; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_50; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_51; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_52; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_53; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_54; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_55; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_56; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_57; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_58; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_59; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_60; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_61; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_62; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_63; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_64; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_65; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_66; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_67; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_68; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_69; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_70; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_71; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_72; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_73; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_74; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_75; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_76; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_77; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_78; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_79; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_80; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_81; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_82; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_83; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_84; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_85; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_86; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_87; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_88; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_89; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_90; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_91; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_92; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_93; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_94; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_95; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_96; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_97; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_98; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_99; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_100; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_101; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_102; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_103; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_104; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_105; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_106; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_107; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_108; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_109; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_110; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_111; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_112; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_113; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_114; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_115; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_116; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_117; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_118; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_119; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_120; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_121; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_122; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_123; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_124; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_125; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_126; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_127; // @[d_cache.scala 22:24]
  reg [31:0] tag_1_0; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_1; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_2; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_3; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_4; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_5; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_6; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_7; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_8; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_9; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_10; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_11; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_12; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_13; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_14; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_15; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_16; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_17; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_18; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_19; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_20; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_21; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_22; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_23; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_24; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_25; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_26; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_27; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_28; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_29; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_30; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_31; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_32; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_33; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_34; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_35; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_36; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_37; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_38; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_39; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_40; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_41; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_42; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_43; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_44; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_45; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_46; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_47; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_48; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_49; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_50; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_51; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_52; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_53; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_54; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_55; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_56; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_57; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_58; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_59; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_60; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_61; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_62; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_63; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_64; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_65; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_66; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_67; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_68; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_69; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_70; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_71; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_72; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_73; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_74; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_75; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_76; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_77; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_78; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_79; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_80; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_81; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_82; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_83; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_84; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_85; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_86; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_87; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_88; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_89; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_90; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_91; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_92; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_93; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_94; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_95; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_96; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_97; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_98; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_99; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_100; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_101; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_102; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_103; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_104; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_105; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_106; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_107; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_108; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_109; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_110; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_111; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_112; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_113; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_114; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_115; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_116; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_117; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_118; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_119; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_120; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_121; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_122; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_123; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_124; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_125; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_126; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_127; // @[d_cache.scala 23:24]
  reg  valid_0_0; // @[d_cache.scala 24:26]
  reg  valid_0_1; // @[d_cache.scala 24:26]
  reg  valid_0_2; // @[d_cache.scala 24:26]
  reg  valid_0_3; // @[d_cache.scala 24:26]
  reg  valid_0_4; // @[d_cache.scala 24:26]
  reg  valid_0_5; // @[d_cache.scala 24:26]
  reg  valid_0_6; // @[d_cache.scala 24:26]
  reg  valid_0_7; // @[d_cache.scala 24:26]
  reg  valid_0_8; // @[d_cache.scala 24:26]
  reg  valid_0_9; // @[d_cache.scala 24:26]
  reg  valid_0_10; // @[d_cache.scala 24:26]
  reg  valid_0_11; // @[d_cache.scala 24:26]
  reg  valid_0_12; // @[d_cache.scala 24:26]
  reg  valid_0_13; // @[d_cache.scala 24:26]
  reg  valid_0_14; // @[d_cache.scala 24:26]
  reg  valid_0_15; // @[d_cache.scala 24:26]
  reg  valid_0_16; // @[d_cache.scala 24:26]
  reg  valid_0_17; // @[d_cache.scala 24:26]
  reg  valid_0_18; // @[d_cache.scala 24:26]
  reg  valid_0_19; // @[d_cache.scala 24:26]
  reg  valid_0_20; // @[d_cache.scala 24:26]
  reg  valid_0_21; // @[d_cache.scala 24:26]
  reg  valid_0_22; // @[d_cache.scala 24:26]
  reg  valid_0_23; // @[d_cache.scala 24:26]
  reg  valid_0_24; // @[d_cache.scala 24:26]
  reg  valid_0_25; // @[d_cache.scala 24:26]
  reg  valid_0_26; // @[d_cache.scala 24:26]
  reg  valid_0_27; // @[d_cache.scala 24:26]
  reg  valid_0_28; // @[d_cache.scala 24:26]
  reg  valid_0_29; // @[d_cache.scala 24:26]
  reg  valid_0_30; // @[d_cache.scala 24:26]
  reg  valid_0_31; // @[d_cache.scala 24:26]
  reg  valid_0_32; // @[d_cache.scala 24:26]
  reg  valid_0_33; // @[d_cache.scala 24:26]
  reg  valid_0_34; // @[d_cache.scala 24:26]
  reg  valid_0_35; // @[d_cache.scala 24:26]
  reg  valid_0_36; // @[d_cache.scala 24:26]
  reg  valid_0_37; // @[d_cache.scala 24:26]
  reg  valid_0_38; // @[d_cache.scala 24:26]
  reg  valid_0_39; // @[d_cache.scala 24:26]
  reg  valid_0_40; // @[d_cache.scala 24:26]
  reg  valid_0_41; // @[d_cache.scala 24:26]
  reg  valid_0_42; // @[d_cache.scala 24:26]
  reg  valid_0_43; // @[d_cache.scala 24:26]
  reg  valid_0_44; // @[d_cache.scala 24:26]
  reg  valid_0_45; // @[d_cache.scala 24:26]
  reg  valid_0_46; // @[d_cache.scala 24:26]
  reg  valid_0_47; // @[d_cache.scala 24:26]
  reg  valid_0_48; // @[d_cache.scala 24:26]
  reg  valid_0_49; // @[d_cache.scala 24:26]
  reg  valid_0_50; // @[d_cache.scala 24:26]
  reg  valid_0_51; // @[d_cache.scala 24:26]
  reg  valid_0_52; // @[d_cache.scala 24:26]
  reg  valid_0_53; // @[d_cache.scala 24:26]
  reg  valid_0_54; // @[d_cache.scala 24:26]
  reg  valid_0_55; // @[d_cache.scala 24:26]
  reg  valid_0_56; // @[d_cache.scala 24:26]
  reg  valid_0_57; // @[d_cache.scala 24:26]
  reg  valid_0_58; // @[d_cache.scala 24:26]
  reg  valid_0_59; // @[d_cache.scala 24:26]
  reg  valid_0_60; // @[d_cache.scala 24:26]
  reg  valid_0_61; // @[d_cache.scala 24:26]
  reg  valid_0_62; // @[d_cache.scala 24:26]
  reg  valid_0_63; // @[d_cache.scala 24:26]
  reg  valid_0_64; // @[d_cache.scala 24:26]
  reg  valid_0_65; // @[d_cache.scala 24:26]
  reg  valid_0_66; // @[d_cache.scala 24:26]
  reg  valid_0_67; // @[d_cache.scala 24:26]
  reg  valid_0_68; // @[d_cache.scala 24:26]
  reg  valid_0_69; // @[d_cache.scala 24:26]
  reg  valid_0_70; // @[d_cache.scala 24:26]
  reg  valid_0_71; // @[d_cache.scala 24:26]
  reg  valid_0_72; // @[d_cache.scala 24:26]
  reg  valid_0_73; // @[d_cache.scala 24:26]
  reg  valid_0_74; // @[d_cache.scala 24:26]
  reg  valid_0_75; // @[d_cache.scala 24:26]
  reg  valid_0_76; // @[d_cache.scala 24:26]
  reg  valid_0_77; // @[d_cache.scala 24:26]
  reg  valid_0_78; // @[d_cache.scala 24:26]
  reg  valid_0_79; // @[d_cache.scala 24:26]
  reg  valid_0_80; // @[d_cache.scala 24:26]
  reg  valid_0_81; // @[d_cache.scala 24:26]
  reg  valid_0_82; // @[d_cache.scala 24:26]
  reg  valid_0_83; // @[d_cache.scala 24:26]
  reg  valid_0_84; // @[d_cache.scala 24:26]
  reg  valid_0_85; // @[d_cache.scala 24:26]
  reg  valid_0_86; // @[d_cache.scala 24:26]
  reg  valid_0_87; // @[d_cache.scala 24:26]
  reg  valid_0_88; // @[d_cache.scala 24:26]
  reg  valid_0_89; // @[d_cache.scala 24:26]
  reg  valid_0_90; // @[d_cache.scala 24:26]
  reg  valid_0_91; // @[d_cache.scala 24:26]
  reg  valid_0_92; // @[d_cache.scala 24:26]
  reg  valid_0_93; // @[d_cache.scala 24:26]
  reg  valid_0_94; // @[d_cache.scala 24:26]
  reg  valid_0_95; // @[d_cache.scala 24:26]
  reg  valid_0_96; // @[d_cache.scala 24:26]
  reg  valid_0_97; // @[d_cache.scala 24:26]
  reg  valid_0_98; // @[d_cache.scala 24:26]
  reg  valid_0_99; // @[d_cache.scala 24:26]
  reg  valid_0_100; // @[d_cache.scala 24:26]
  reg  valid_0_101; // @[d_cache.scala 24:26]
  reg  valid_0_102; // @[d_cache.scala 24:26]
  reg  valid_0_103; // @[d_cache.scala 24:26]
  reg  valid_0_104; // @[d_cache.scala 24:26]
  reg  valid_0_105; // @[d_cache.scala 24:26]
  reg  valid_0_106; // @[d_cache.scala 24:26]
  reg  valid_0_107; // @[d_cache.scala 24:26]
  reg  valid_0_108; // @[d_cache.scala 24:26]
  reg  valid_0_109; // @[d_cache.scala 24:26]
  reg  valid_0_110; // @[d_cache.scala 24:26]
  reg  valid_0_111; // @[d_cache.scala 24:26]
  reg  valid_0_112; // @[d_cache.scala 24:26]
  reg  valid_0_113; // @[d_cache.scala 24:26]
  reg  valid_0_114; // @[d_cache.scala 24:26]
  reg  valid_0_115; // @[d_cache.scala 24:26]
  reg  valid_0_116; // @[d_cache.scala 24:26]
  reg  valid_0_117; // @[d_cache.scala 24:26]
  reg  valid_0_118; // @[d_cache.scala 24:26]
  reg  valid_0_119; // @[d_cache.scala 24:26]
  reg  valid_0_120; // @[d_cache.scala 24:26]
  reg  valid_0_121; // @[d_cache.scala 24:26]
  reg  valid_0_122; // @[d_cache.scala 24:26]
  reg  valid_0_123; // @[d_cache.scala 24:26]
  reg  valid_0_124; // @[d_cache.scala 24:26]
  reg  valid_0_125; // @[d_cache.scala 24:26]
  reg  valid_0_126; // @[d_cache.scala 24:26]
  reg  valid_0_127; // @[d_cache.scala 24:26]
  reg  valid_1_0; // @[d_cache.scala 25:26]
  reg  valid_1_1; // @[d_cache.scala 25:26]
  reg  valid_1_2; // @[d_cache.scala 25:26]
  reg  valid_1_3; // @[d_cache.scala 25:26]
  reg  valid_1_4; // @[d_cache.scala 25:26]
  reg  valid_1_5; // @[d_cache.scala 25:26]
  reg  valid_1_6; // @[d_cache.scala 25:26]
  reg  valid_1_7; // @[d_cache.scala 25:26]
  reg  valid_1_8; // @[d_cache.scala 25:26]
  reg  valid_1_9; // @[d_cache.scala 25:26]
  reg  valid_1_10; // @[d_cache.scala 25:26]
  reg  valid_1_11; // @[d_cache.scala 25:26]
  reg  valid_1_12; // @[d_cache.scala 25:26]
  reg  valid_1_13; // @[d_cache.scala 25:26]
  reg  valid_1_14; // @[d_cache.scala 25:26]
  reg  valid_1_15; // @[d_cache.scala 25:26]
  reg  valid_1_16; // @[d_cache.scala 25:26]
  reg  valid_1_17; // @[d_cache.scala 25:26]
  reg  valid_1_18; // @[d_cache.scala 25:26]
  reg  valid_1_19; // @[d_cache.scala 25:26]
  reg  valid_1_20; // @[d_cache.scala 25:26]
  reg  valid_1_21; // @[d_cache.scala 25:26]
  reg  valid_1_22; // @[d_cache.scala 25:26]
  reg  valid_1_23; // @[d_cache.scala 25:26]
  reg  valid_1_24; // @[d_cache.scala 25:26]
  reg  valid_1_25; // @[d_cache.scala 25:26]
  reg  valid_1_26; // @[d_cache.scala 25:26]
  reg  valid_1_27; // @[d_cache.scala 25:26]
  reg  valid_1_28; // @[d_cache.scala 25:26]
  reg  valid_1_29; // @[d_cache.scala 25:26]
  reg  valid_1_30; // @[d_cache.scala 25:26]
  reg  valid_1_31; // @[d_cache.scala 25:26]
  reg  valid_1_32; // @[d_cache.scala 25:26]
  reg  valid_1_33; // @[d_cache.scala 25:26]
  reg  valid_1_34; // @[d_cache.scala 25:26]
  reg  valid_1_35; // @[d_cache.scala 25:26]
  reg  valid_1_36; // @[d_cache.scala 25:26]
  reg  valid_1_37; // @[d_cache.scala 25:26]
  reg  valid_1_38; // @[d_cache.scala 25:26]
  reg  valid_1_39; // @[d_cache.scala 25:26]
  reg  valid_1_40; // @[d_cache.scala 25:26]
  reg  valid_1_41; // @[d_cache.scala 25:26]
  reg  valid_1_42; // @[d_cache.scala 25:26]
  reg  valid_1_43; // @[d_cache.scala 25:26]
  reg  valid_1_44; // @[d_cache.scala 25:26]
  reg  valid_1_45; // @[d_cache.scala 25:26]
  reg  valid_1_46; // @[d_cache.scala 25:26]
  reg  valid_1_47; // @[d_cache.scala 25:26]
  reg  valid_1_48; // @[d_cache.scala 25:26]
  reg  valid_1_49; // @[d_cache.scala 25:26]
  reg  valid_1_50; // @[d_cache.scala 25:26]
  reg  valid_1_51; // @[d_cache.scala 25:26]
  reg  valid_1_52; // @[d_cache.scala 25:26]
  reg  valid_1_53; // @[d_cache.scala 25:26]
  reg  valid_1_54; // @[d_cache.scala 25:26]
  reg  valid_1_55; // @[d_cache.scala 25:26]
  reg  valid_1_56; // @[d_cache.scala 25:26]
  reg  valid_1_57; // @[d_cache.scala 25:26]
  reg  valid_1_58; // @[d_cache.scala 25:26]
  reg  valid_1_59; // @[d_cache.scala 25:26]
  reg  valid_1_60; // @[d_cache.scala 25:26]
  reg  valid_1_61; // @[d_cache.scala 25:26]
  reg  valid_1_62; // @[d_cache.scala 25:26]
  reg  valid_1_63; // @[d_cache.scala 25:26]
  reg  valid_1_64; // @[d_cache.scala 25:26]
  reg  valid_1_65; // @[d_cache.scala 25:26]
  reg  valid_1_66; // @[d_cache.scala 25:26]
  reg  valid_1_67; // @[d_cache.scala 25:26]
  reg  valid_1_68; // @[d_cache.scala 25:26]
  reg  valid_1_69; // @[d_cache.scala 25:26]
  reg  valid_1_70; // @[d_cache.scala 25:26]
  reg  valid_1_71; // @[d_cache.scala 25:26]
  reg  valid_1_72; // @[d_cache.scala 25:26]
  reg  valid_1_73; // @[d_cache.scala 25:26]
  reg  valid_1_74; // @[d_cache.scala 25:26]
  reg  valid_1_75; // @[d_cache.scala 25:26]
  reg  valid_1_76; // @[d_cache.scala 25:26]
  reg  valid_1_77; // @[d_cache.scala 25:26]
  reg  valid_1_78; // @[d_cache.scala 25:26]
  reg  valid_1_79; // @[d_cache.scala 25:26]
  reg  valid_1_80; // @[d_cache.scala 25:26]
  reg  valid_1_81; // @[d_cache.scala 25:26]
  reg  valid_1_82; // @[d_cache.scala 25:26]
  reg  valid_1_83; // @[d_cache.scala 25:26]
  reg  valid_1_84; // @[d_cache.scala 25:26]
  reg  valid_1_85; // @[d_cache.scala 25:26]
  reg  valid_1_86; // @[d_cache.scala 25:26]
  reg  valid_1_87; // @[d_cache.scala 25:26]
  reg  valid_1_88; // @[d_cache.scala 25:26]
  reg  valid_1_89; // @[d_cache.scala 25:26]
  reg  valid_1_90; // @[d_cache.scala 25:26]
  reg  valid_1_91; // @[d_cache.scala 25:26]
  reg  valid_1_92; // @[d_cache.scala 25:26]
  reg  valid_1_93; // @[d_cache.scala 25:26]
  reg  valid_1_94; // @[d_cache.scala 25:26]
  reg  valid_1_95; // @[d_cache.scala 25:26]
  reg  valid_1_96; // @[d_cache.scala 25:26]
  reg  valid_1_97; // @[d_cache.scala 25:26]
  reg  valid_1_98; // @[d_cache.scala 25:26]
  reg  valid_1_99; // @[d_cache.scala 25:26]
  reg  valid_1_100; // @[d_cache.scala 25:26]
  reg  valid_1_101; // @[d_cache.scala 25:26]
  reg  valid_1_102; // @[d_cache.scala 25:26]
  reg  valid_1_103; // @[d_cache.scala 25:26]
  reg  valid_1_104; // @[d_cache.scala 25:26]
  reg  valid_1_105; // @[d_cache.scala 25:26]
  reg  valid_1_106; // @[d_cache.scala 25:26]
  reg  valid_1_107; // @[d_cache.scala 25:26]
  reg  valid_1_108; // @[d_cache.scala 25:26]
  reg  valid_1_109; // @[d_cache.scala 25:26]
  reg  valid_1_110; // @[d_cache.scala 25:26]
  reg  valid_1_111; // @[d_cache.scala 25:26]
  reg  valid_1_112; // @[d_cache.scala 25:26]
  reg  valid_1_113; // @[d_cache.scala 25:26]
  reg  valid_1_114; // @[d_cache.scala 25:26]
  reg  valid_1_115; // @[d_cache.scala 25:26]
  reg  valid_1_116; // @[d_cache.scala 25:26]
  reg  valid_1_117; // @[d_cache.scala 25:26]
  reg  valid_1_118; // @[d_cache.scala 25:26]
  reg  valid_1_119; // @[d_cache.scala 25:26]
  reg  valid_1_120; // @[d_cache.scala 25:26]
  reg  valid_1_121; // @[d_cache.scala 25:26]
  reg  valid_1_122; // @[d_cache.scala 25:26]
  reg  valid_1_123; // @[d_cache.scala 25:26]
  reg  valid_1_124; // @[d_cache.scala 25:26]
  reg  valid_1_125; // @[d_cache.scala 25:26]
  reg  valid_1_126; // @[d_cache.scala 25:26]
  reg  valid_1_127; // @[d_cache.scala 25:26]
  reg  dirty_0_0; // @[d_cache.scala 26:26]
  reg  dirty_0_1; // @[d_cache.scala 26:26]
  reg  dirty_0_2; // @[d_cache.scala 26:26]
  reg  dirty_0_3; // @[d_cache.scala 26:26]
  reg  dirty_0_4; // @[d_cache.scala 26:26]
  reg  dirty_0_5; // @[d_cache.scala 26:26]
  reg  dirty_0_6; // @[d_cache.scala 26:26]
  reg  dirty_0_7; // @[d_cache.scala 26:26]
  reg  dirty_0_8; // @[d_cache.scala 26:26]
  reg  dirty_0_9; // @[d_cache.scala 26:26]
  reg  dirty_0_10; // @[d_cache.scala 26:26]
  reg  dirty_0_11; // @[d_cache.scala 26:26]
  reg  dirty_0_12; // @[d_cache.scala 26:26]
  reg  dirty_0_13; // @[d_cache.scala 26:26]
  reg  dirty_0_14; // @[d_cache.scala 26:26]
  reg  dirty_0_15; // @[d_cache.scala 26:26]
  reg  dirty_0_16; // @[d_cache.scala 26:26]
  reg  dirty_0_17; // @[d_cache.scala 26:26]
  reg  dirty_0_18; // @[d_cache.scala 26:26]
  reg  dirty_0_19; // @[d_cache.scala 26:26]
  reg  dirty_0_20; // @[d_cache.scala 26:26]
  reg  dirty_0_21; // @[d_cache.scala 26:26]
  reg  dirty_0_22; // @[d_cache.scala 26:26]
  reg  dirty_0_23; // @[d_cache.scala 26:26]
  reg  dirty_0_24; // @[d_cache.scala 26:26]
  reg  dirty_0_25; // @[d_cache.scala 26:26]
  reg  dirty_0_26; // @[d_cache.scala 26:26]
  reg  dirty_0_27; // @[d_cache.scala 26:26]
  reg  dirty_0_28; // @[d_cache.scala 26:26]
  reg  dirty_0_29; // @[d_cache.scala 26:26]
  reg  dirty_0_30; // @[d_cache.scala 26:26]
  reg  dirty_0_31; // @[d_cache.scala 26:26]
  reg  dirty_0_32; // @[d_cache.scala 26:26]
  reg  dirty_0_33; // @[d_cache.scala 26:26]
  reg  dirty_0_34; // @[d_cache.scala 26:26]
  reg  dirty_0_35; // @[d_cache.scala 26:26]
  reg  dirty_0_36; // @[d_cache.scala 26:26]
  reg  dirty_0_37; // @[d_cache.scala 26:26]
  reg  dirty_0_38; // @[d_cache.scala 26:26]
  reg  dirty_0_39; // @[d_cache.scala 26:26]
  reg  dirty_0_40; // @[d_cache.scala 26:26]
  reg  dirty_0_41; // @[d_cache.scala 26:26]
  reg  dirty_0_42; // @[d_cache.scala 26:26]
  reg  dirty_0_43; // @[d_cache.scala 26:26]
  reg  dirty_0_44; // @[d_cache.scala 26:26]
  reg  dirty_0_45; // @[d_cache.scala 26:26]
  reg  dirty_0_46; // @[d_cache.scala 26:26]
  reg  dirty_0_47; // @[d_cache.scala 26:26]
  reg  dirty_0_48; // @[d_cache.scala 26:26]
  reg  dirty_0_49; // @[d_cache.scala 26:26]
  reg  dirty_0_50; // @[d_cache.scala 26:26]
  reg  dirty_0_51; // @[d_cache.scala 26:26]
  reg  dirty_0_52; // @[d_cache.scala 26:26]
  reg  dirty_0_53; // @[d_cache.scala 26:26]
  reg  dirty_0_54; // @[d_cache.scala 26:26]
  reg  dirty_0_55; // @[d_cache.scala 26:26]
  reg  dirty_0_56; // @[d_cache.scala 26:26]
  reg  dirty_0_57; // @[d_cache.scala 26:26]
  reg  dirty_0_58; // @[d_cache.scala 26:26]
  reg  dirty_0_59; // @[d_cache.scala 26:26]
  reg  dirty_0_60; // @[d_cache.scala 26:26]
  reg  dirty_0_61; // @[d_cache.scala 26:26]
  reg  dirty_0_62; // @[d_cache.scala 26:26]
  reg  dirty_0_63; // @[d_cache.scala 26:26]
  reg  dirty_0_64; // @[d_cache.scala 26:26]
  reg  dirty_0_65; // @[d_cache.scala 26:26]
  reg  dirty_0_66; // @[d_cache.scala 26:26]
  reg  dirty_0_67; // @[d_cache.scala 26:26]
  reg  dirty_0_68; // @[d_cache.scala 26:26]
  reg  dirty_0_69; // @[d_cache.scala 26:26]
  reg  dirty_0_70; // @[d_cache.scala 26:26]
  reg  dirty_0_71; // @[d_cache.scala 26:26]
  reg  dirty_0_72; // @[d_cache.scala 26:26]
  reg  dirty_0_73; // @[d_cache.scala 26:26]
  reg  dirty_0_74; // @[d_cache.scala 26:26]
  reg  dirty_0_75; // @[d_cache.scala 26:26]
  reg  dirty_0_76; // @[d_cache.scala 26:26]
  reg  dirty_0_77; // @[d_cache.scala 26:26]
  reg  dirty_0_78; // @[d_cache.scala 26:26]
  reg  dirty_0_79; // @[d_cache.scala 26:26]
  reg  dirty_0_80; // @[d_cache.scala 26:26]
  reg  dirty_0_81; // @[d_cache.scala 26:26]
  reg  dirty_0_82; // @[d_cache.scala 26:26]
  reg  dirty_0_83; // @[d_cache.scala 26:26]
  reg  dirty_0_84; // @[d_cache.scala 26:26]
  reg  dirty_0_85; // @[d_cache.scala 26:26]
  reg  dirty_0_86; // @[d_cache.scala 26:26]
  reg  dirty_0_87; // @[d_cache.scala 26:26]
  reg  dirty_0_88; // @[d_cache.scala 26:26]
  reg  dirty_0_89; // @[d_cache.scala 26:26]
  reg  dirty_0_90; // @[d_cache.scala 26:26]
  reg  dirty_0_91; // @[d_cache.scala 26:26]
  reg  dirty_0_92; // @[d_cache.scala 26:26]
  reg  dirty_0_93; // @[d_cache.scala 26:26]
  reg  dirty_0_94; // @[d_cache.scala 26:26]
  reg  dirty_0_95; // @[d_cache.scala 26:26]
  reg  dirty_0_96; // @[d_cache.scala 26:26]
  reg  dirty_0_97; // @[d_cache.scala 26:26]
  reg  dirty_0_98; // @[d_cache.scala 26:26]
  reg  dirty_0_99; // @[d_cache.scala 26:26]
  reg  dirty_0_100; // @[d_cache.scala 26:26]
  reg  dirty_0_101; // @[d_cache.scala 26:26]
  reg  dirty_0_102; // @[d_cache.scala 26:26]
  reg  dirty_0_103; // @[d_cache.scala 26:26]
  reg  dirty_0_104; // @[d_cache.scala 26:26]
  reg  dirty_0_105; // @[d_cache.scala 26:26]
  reg  dirty_0_106; // @[d_cache.scala 26:26]
  reg  dirty_0_107; // @[d_cache.scala 26:26]
  reg  dirty_0_108; // @[d_cache.scala 26:26]
  reg  dirty_0_109; // @[d_cache.scala 26:26]
  reg  dirty_0_110; // @[d_cache.scala 26:26]
  reg  dirty_0_111; // @[d_cache.scala 26:26]
  reg  dirty_0_112; // @[d_cache.scala 26:26]
  reg  dirty_0_113; // @[d_cache.scala 26:26]
  reg  dirty_0_114; // @[d_cache.scala 26:26]
  reg  dirty_0_115; // @[d_cache.scala 26:26]
  reg  dirty_0_116; // @[d_cache.scala 26:26]
  reg  dirty_0_117; // @[d_cache.scala 26:26]
  reg  dirty_0_118; // @[d_cache.scala 26:26]
  reg  dirty_0_119; // @[d_cache.scala 26:26]
  reg  dirty_0_120; // @[d_cache.scala 26:26]
  reg  dirty_0_121; // @[d_cache.scala 26:26]
  reg  dirty_0_122; // @[d_cache.scala 26:26]
  reg  dirty_0_123; // @[d_cache.scala 26:26]
  reg  dirty_0_124; // @[d_cache.scala 26:26]
  reg  dirty_0_125; // @[d_cache.scala 26:26]
  reg  dirty_0_126; // @[d_cache.scala 26:26]
  reg  dirty_0_127; // @[d_cache.scala 26:26]
  reg  dirty_1_0; // @[d_cache.scala 27:26]
  reg  dirty_1_1; // @[d_cache.scala 27:26]
  reg  dirty_1_2; // @[d_cache.scala 27:26]
  reg  dirty_1_3; // @[d_cache.scala 27:26]
  reg  dirty_1_4; // @[d_cache.scala 27:26]
  reg  dirty_1_5; // @[d_cache.scala 27:26]
  reg  dirty_1_6; // @[d_cache.scala 27:26]
  reg  dirty_1_7; // @[d_cache.scala 27:26]
  reg  dirty_1_8; // @[d_cache.scala 27:26]
  reg  dirty_1_9; // @[d_cache.scala 27:26]
  reg  dirty_1_10; // @[d_cache.scala 27:26]
  reg  dirty_1_11; // @[d_cache.scala 27:26]
  reg  dirty_1_12; // @[d_cache.scala 27:26]
  reg  dirty_1_13; // @[d_cache.scala 27:26]
  reg  dirty_1_14; // @[d_cache.scala 27:26]
  reg  dirty_1_15; // @[d_cache.scala 27:26]
  reg  dirty_1_16; // @[d_cache.scala 27:26]
  reg  dirty_1_17; // @[d_cache.scala 27:26]
  reg  dirty_1_18; // @[d_cache.scala 27:26]
  reg  dirty_1_19; // @[d_cache.scala 27:26]
  reg  dirty_1_20; // @[d_cache.scala 27:26]
  reg  dirty_1_21; // @[d_cache.scala 27:26]
  reg  dirty_1_22; // @[d_cache.scala 27:26]
  reg  dirty_1_23; // @[d_cache.scala 27:26]
  reg  dirty_1_24; // @[d_cache.scala 27:26]
  reg  dirty_1_25; // @[d_cache.scala 27:26]
  reg  dirty_1_26; // @[d_cache.scala 27:26]
  reg  dirty_1_27; // @[d_cache.scala 27:26]
  reg  dirty_1_28; // @[d_cache.scala 27:26]
  reg  dirty_1_29; // @[d_cache.scala 27:26]
  reg  dirty_1_30; // @[d_cache.scala 27:26]
  reg  dirty_1_31; // @[d_cache.scala 27:26]
  reg  dirty_1_32; // @[d_cache.scala 27:26]
  reg  dirty_1_33; // @[d_cache.scala 27:26]
  reg  dirty_1_34; // @[d_cache.scala 27:26]
  reg  dirty_1_35; // @[d_cache.scala 27:26]
  reg  dirty_1_36; // @[d_cache.scala 27:26]
  reg  dirty_1_37; // @[d_cache.scala 27:26]
  reg  dirty_1_38; // @[d_cache.scala 27:26]
  reg  dirty_1_39; // @[d_cache.scala 27:26]
  reg  dirty_1_40; // @[d_cache.scala 27:26]
  reg  dirty_1_41; // @[d_cache.scala 27:26]
  reg  dirty_1_42; // @[d_cache.scala 27:26]
  reg  dirty_1_43; // @[d_cache.scala 27:26]
  reg  dirty_1_44; // @[d_cache.scala 27:26]
  reg  dirty_1_45; // @[d_cache.scala 27:26]
  reg  dirty_1_46; // @[d_cache.scala 27:26]
  reg  dirty_1_47; // @[d_cache.scala 27:26]
  reg  dirty_1_48; // @[d_cache.scala 27:26]
  reg  dirty_1_49; // @[d_cache.scala 27:26]
  reg  dirty_1_50; // @[d_cache.scala 27:26]
  reg  dirty_1_51; // @[d_cache.scala 27:26]
  reg  dirty_1_52; // @[d_cache.scala 27:26]
  reg  dirty_1_53; // @[d_cache.scala 27:26]
  reg  dirty_1_54; // @[d_cache.scala 27:26]
  reg  dirty_1_55; // @[d_cache.scala 27:26]
  reg  dirty_1_56; // @[d_cache.scala 27:26]
  reg  dirty_1_57; // @[d_cache.scala 27:26]
  reg  dirty_1_58; // @[d_cache.scala 27:26]
  reg  dirty_1_59; // @[d_cache.scala 27:26]
  reg  dirty_1_60; // @[d_cache.scala 27:26]
  reg  dirty_1_61; // @[d_cache.scala 27:26]
  reg  dirty_1_62; // @[d_cache.scala 27:26]
  reg  dirty_1_63; // @[d_cache.scala 27:26]
  reg  dirty_1_64; // @[d_cache.scala 27:26]
  reg  dirty_1_65; // @[d_cache.scala 27:26]
  reg  dirty_1_66; // @[d_cache.scala 27:26]
  reg  dirty_1_67; // @[d_cache.scala 27:26]
  reg  dirty_1_68; // @[d_cache.scala 27:26]
  reg  dirty_1_69; // @[d_cache.scala 27:26]
  reg  dirty_1_70; // @[d_cache.scala 27:26]
  reg  dirty_1_71; // @[d_cache.scala 27:26]
  reg  dirty_1_72; // @[d_cache.scala 27:26]
  reg  dirty_1_73; // @[d_cache.scala 27:26]
  reg  dirty_1_74; // @[d_cache.scala 27:26]
  reg  dirty_1_75; // @[d_cache.scala 27:26]
  reg  dirty_1_76; // @[d_cache.scala 27:26]
  reg  dirty_1_77; // @[d_cache.scala 27:26]
  reg  dirty_1_78; // @[d_cache.scala 27:26]
  reg  dirty_1_79; // @[d_cache.scala 27:26]
  reg  dirty_1_80; // @[d_cache.scala 27:26]
  reg  dirty_1_81; // @[d_cache.scala 27:26]
  reg  dirty_1_82; // @[d_cache.scala 27:26]
  reg  dirty_1_83; // @[d_cache.scala 27:26]
  reg  dirty_1_84; // @[d_cache.scala 27:26]
  reg  dirty_1_85; // @[d_cache.scala 27:26]
  reg  dirty_1_86; // @[d_cache.scala 27:26]
  reg  dirty_1_87; // @[d_cache.scala 27:26]
  reg  dirty_1_88; // @[d_cache.scala 27:26]
  reg  dirty_1_89; // @[d_cache.scala 27:26]
  reg  dirty_1_90; // @[d_cache.scala 27:26]
  reg  dirty_1_91; // @[d_cache.scala 27:26]
  reg  dirty_1_92; // @[d_cache.scala 27:26]
  reg  dirty_1_93; // @[d_cache.scala 27:26]
  reg  dirty_1_94; // @[d_cache.scala 27:26]
  reg  dirty_1_95; // @[d_cache.scala 27:26]
  reg  dirty_1_96; // @[d_cache.scala 27:26]
  reg  dirty_1_97; // @[d_cache.scala 27:26]
  reg  dirty_1_98; // @[d_cache.scala 27:26]
  reg  dirty_1_99; // @[d_cache.scala 27:26]
  reg  dirty_1_100; // @[d_cache.scala 27:26]
  reg  dirty_1_101; // @[d_cache.scala 27:26]
  reg  dirty_1_102; // @[d_cache.scala 27:26]
  reg  dirty_1_103; // @[d_cache.scala 27:26]
  reg  dirty_1_104; // @[d_cache.scala 27:26]
  reg  dirty_1_105; // @[d_cache.scala 27:26]
  reg  dirty_1_106; // @[d_cache.scala 27:26]
  reg  dirty_1_107; // @[d_cache.scala 27:26]
  reg  dirty_1_108; // @[d_cache.scala 27:26]
  reg  dirty_1_109; // @[d_cache.scala 27:26]
  reg  dirty_1_110; // @[d_cache.scala 27:26]
  reg  dirty_1_111; // @[d_cache.scala 27:26]
  reg  dirty_1_112; // @[d_cache.scala 27:26]
  reg  dirty_1_113; // @[d_cache.scala 27:26]
  reg  dirty_1_114; // @[d_cache.scala 27:26]
  reg  dirty_1_115; // @[d_cache.scala 27:26]
  reg  dirty_1_116; // @[d_cache.scala 27:26]
  reg  dirty_1_117; // @[d_cache.scala 27:26]
  reg  dirty_1_118; // @[d_cache.scala 27:26]
  reg  dirty_1_119; // @[d_cache.scala 27:26]
  reg  dirty_1_120; // @[d_cache.scala 27:26]
  reg  dirty_1_121; // @[d_cache.scala 27:26]
  reg  dirty_1_122; // @[d_cache.scala 27:26]
  reg  dirty_1_123; // @[d_cache.scala 27:26]
  reg  dirty_1_124; // @[d_cache.scala 27:26]
  reg  dirty_1_125; // @[d_cache.scala 27:26]
  reg  dirty_1_126; // @[d_cache.scala 27:26]
  reg  dirty_1_127; // @[d_cache.scala 27:26]
  reg  way0_hit; // @[d_cache.scala 28:27]
  reg  way1_hit; // @[d_cache.scala 29:27]
  reg [63:0] write_back_data; // @[d_cache.scala 31:34]
  reg [31:0] write_back_addr; // @[d_cache.scala 32:34]
  reg [1:0] unuse_way; // @[d_cache.scala 35:28]
  reg [63:0] receive_data; // @[d_cache.scala 36:31]
  reg  quene; // @[d_cache.scala 37:24]
  wire [2:0] offset = io_from_lsu_araddr[2:0]; // @[d_cache.scala 39:36]
  wire [21:0] tag = io_from_lsu_araddr[31:10]; // @[d_cache.scala 41:33]
  wire [5:0] _shift_bit_T_8 = offset == 3'h7 ? 6'h38 : 6'h0; // @[d_cache.scala 50:24]
  wire [5:0] _shift_bit_T_9 = offset == 3'h6 ? 6'h30 : _shift_bit_T_8; // @[d_cache.scala 49:24]
  wire [5:0] _shift_bit_T_10 = offset == 3'h5 ? 6'h28 : _shift_bit_T_9; // @[d_cache.scala 48:24]
  wire [5:0] _shift_bit_T_11 = offset == 3'h4 ? 6'h20 : _shift_bit_T_10; // @[d_cache.scala 47:24]
  wire [5:0] _shift_bit_T_12 = offset == 3'h3 ? 6'h18 : _shift_bit_T_11; // @[d_cache.scala 46:24]
  wire [5:0] _shift_bit_T_13 = offset == 3'h2 ? 6'h10 : _shift_bit_T_12; // @[d_cache.scala 45:24]
  wire [5:0] _shift_bit_T_14 = offset == 3'h1 ? 6'h8 : _shift_bit_T_13; // @[d_cache.scala 44:24]
  wire [5:0] shift_bit = offset == 3'h0 ? 6'h0 : _shift_bit_T_14; // @[d_cache.scala 43:24]
  wire [63:0] _wmask_T_4 = io_from_lsu_wstrb == 8'hff ? 64'hffffffffffffffff : 64'h0; // @[d_cache.scala 55:20]
  wire [63:0] _wmask_T_5 = io_from_lsu_wstrb == 8'hf ? 64'hffffffff : _wmask_T_4; // @[d_cache.scala 54:20]
  wire [63:0] _wmask_T_6 = io_from_lsu_wstrb == 8'h3 ? 64'hffff : _wmask_T_5; // @[d_cache.scala 53:20]
  wire [63:0] wmask = io_from_lsu_wstrb == 8'h1 ? 64'hff : _wmask_T_6; // @[d_cache.scala 52:20]
  wire [31:0] index = {{25'd0}, io_from_lsu_araddr[9:3]}; // @[d_cache.scala 38:21 40:11]
  wire [31:0] _GEN_1 = 7'h1 == index[6:0] ? tag_0_1 : tag_0_0; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_2 = 7'h2 == index[6:0] ? tag_0_2 : _GEN_1; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_3 = 7'h3 == index[6:0] ? tag_0_3 : _GEN_2; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_4 = 7'h4 == index[6:0] ? tag_0_4 : _GEN_3; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_5 = 7'h5 == index[6:0] ? tag_0_5 : _GEN_4; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_6 = 7'h6 == index[6:0] ? tag_0_6 : _GEN_5; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_7 = 7'h7 == index[6:0] ? tag_0_7 : _GEN_6; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_8 = 7'h8 == index[6:0] ? tag_0_8 : _GEN_7; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_9 = 7'h9 == index[6:0] ? tag_0_9 : _GEN_8; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_10 = 7'ha == index[6:0] ? tag_0_10 : _GEN_9; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_11 = 7'hb == index[6:0] ? tag_0_11 : _GEN_10; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_12 = 7'hc == index[6:0] ? tag_0_12 : _GEN_11; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_13 = 7'hd == index[6:0] ? tag_0_13 : _GEN_12; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_14 = 7'he == index[6:0] ? tag_0_14 : _GEN_13; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_15 = 7'hf == index[6:0] ? tag_0_15 : _GEN_14; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_16 = 7'h10 == index[6:0] ? tag_0_16 : _GEN_15; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_17 = 7'h11 == index[6:0] ? tag_0_17 : _GEN_16; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_18 = 7'h12 == index[6:0] ? tag_0_18 : _GEN_17; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_19 = 7'h13 == index[6:0] ? tag_0_19 : _GEN_18; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_20 = 7'h14 == index[6:0] ? tag_0_20 : _GEN_19; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_21 = 7'h15 == index[6:0] ? tag_0_21 : _GEN_20; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_22 = 7'h16 == index[6:0] ? tag_0_22 : _GEN_21; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_23 = 7'h17 == index[6:0] ? tag_0_23 : _GEN_22; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_24 = 7'h18 == index[6:0] ? tag_0_24 : _GEN_23; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_25 = 7'h19 == index[6:0] ? tag_0_25 : _GEN_24; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_26 = 7'h1a == index[6:0] ? tag_0_26 : _GEN_25; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_27 = 7'h1b == index[6:0] ? tag_0_27 : _GEN_26; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_28 = 7'h1c == index[6:0] ? tag_0_28 : _GEN_27; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_29 = 7'h1d == index[6:0] ? tag_0_29 : _GEN_28; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_30 = 7'h1e == index[6:0] ? tag_0_30 : _GEN_29; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_31 = 7'h1f == index[6:0] ? tag_0_31 : _GEN_30; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_32 = 7'h20 == index[6:0] ? tag_0_32 : _GEN_31; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_33 = 7'h21 == index[6:0] ? tag_0_33 : _GEN_32; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_34 = 7'h22 == index[6:0] ? tag_0_34 : _GEN_33; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_35 = 7'h23 == index[6:0] ? tag_0_35 : _GEN_34; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_36 = 7'h24 == index[6:0] ? tag_0_36 : _GEN_35; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_37 = 7'h25 == index[6:0] ? tag_0_37 : _GEN_36; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_38 = 7'h26 == index[6:0] ? tag_0_38 : _GEN_37; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_39 = 7'h27 == index[6:0] ? tag_0_39 : _GEN_38; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_40 = 7'h28 == index[6:0] ? tag_0_40 : _GEN_39; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_41 = 7'h29 == index[6:0] ? tag_0_41 : _GEN_40; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_42 = 7'h2a == index[6:0] ? tag_0_42 : _GEN_41; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_43 = 7'h2b == index[6:0] ? tag_0_43 : _GEN_42; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_44 = 7'h2c == index[6:0] ? tag_0_44 : _GEN_43; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_45 = 7'h2d == index[6:0] ? tag_0_45 : _GEN_44; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_46 = 7'h2e == index[6:0] ? tag_0_46 : _GEN_45; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_47 = 7'h2f == index[6:0] ? tag_0_47 : _GEN_46; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_48 = 7'h30 == index[6:0] ? tag_0_48 : _GEN_47; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_49 = 7'h31 == index[6:0] ? tag_0_49 : _GEN_48; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_50 = 7'h32 == index[6:0] ? tag_0_50 : _GEN_49; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_51 = 7'h33 == index[6:0] ? tag_0_51 : _GEN_50; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_52 = 7'h34 == index[6:0] ? tag_0_52 : _GEN_51; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_53 = 7'h35 == index[6:0] ? tag_0_53 : _GEN_52; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_54 = 7'h36 == index[6:0] ? tag_0_54 : _GEN_53; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_55 = 7'h37 == index[6:0] ? tag_0_55 : _GEN_54; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_56 = 7'h38 == index[6:0] ? tag_0_56 : _GEN_55; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_57 = 7'h39 == index[6:0] ? tag_0_57 : _GEN_56; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_58 = 7'h3a == index[6:0] ? tag_0_58 : _GEN_57; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_59 = 7'h3b == index[6:0] ? tag_0_59 : _GEN_58; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_60 = 7'h3c == index[6:0] ? tag_0_60 : _GEN_59; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_61 = 7'h3d == index[6:0] ? tag_0_61 : _GEN_60; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_62 = 7'h3e == index[6:0] ? tag_0_62 : _GEN_61; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_63 = 7'h3f == index[6:0] ? tag_0_63 : _GEN_62; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_64 = 7'h40 == index[6:0] ? tag_0_64 : _GEN_63; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_65 = 7'h41 == index[6:0] ? tag_0_65 : _GEN_64; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_66 = 7'h42 == index[6:0] ? tag_0_66 : _GEN_65; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_67 = 7'h43 == index[6:0] ? tag_0_67 : _GEN_66; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_68 = 7'h44 == index[6:0] ? tag_0_68 : _GEN_67; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_69 = 7'h45 == index[6:0] ? tag_0_69 : _GEN_68; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_70 = 7'h46 == index[6:0] ? tag_0_70 : _GEN_69; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_71 = 7'h47 == index[6:0] ? tag_0_71 : _GEN_70; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_72 = 7'h48 == index[6:0] ? tag_0_72 : _GEN_71; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_73 = 7'h49 == index[6:0] ? tag_0_73 : _GEN_72; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_74 = 7'h4a == index[6:0] ? tag_0_74 : _GEN_73; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_75 = 7'h4b == index[6:0] ? tag_0_75 : _GEN_74; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_76 = 7'h4c == index[6:0] ? tag_0_76 : _GEN_75; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_77 = 7'h4d == index[6:0] ? tag_0_77 : _GEN_76; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_78 = 7'h4e == index[6:0] ? tag_0_78 : _GEN_77; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_79 = 7'h4f == index[6:0] ? tag_0_79 : _GEN_78; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_80 = 7'h50 == index[6:0] ? tag_0_80 : _GEN_79; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_81 = 7'h51 == index[6:0] ? tag_0_81 : _GEN_80; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_82 = 7'h52 == index[6:0] ? tag_0_82 : _GEN_81; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_83 = 7'h53 == index[6:0] ? tag_0_83 : _GEN_82; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_84 = 7'h54 == index[6:0] ? tag_0_84 : _GEN_83; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_85 = 7'h55 == index[6:0] ? tag_0_85 : _GEN_84; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_86 = 7'h56 == index[6:0] ? tag_0_86 : _GEN_85; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_87 = 7'h57 == index[6:0] ? tag_0_87 : _GEN_86; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_88 = 7'h58 == index[6:0] ? tag_0_88 : _GEN_87; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_89 = 7'h59 == index[6:0] ? tag_0_89 : _GEN_88; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_90 = 7'h5a == index[6:0] ? tag_0_90 : _GEN_89; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_91 = 7'h5b == index[6:0] ? tag_0_91 : _GEN_90; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_92 = 7'h5c == index[6:0] ? tag_0_92 : _GEN_91; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_93 = 7'h5d == index[6:0] ? tag_0_93 : _GEN_92; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_94 = 7'h5e == index[6:0] ? tag_0_94 : _GEN_93; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_95 = 7'h5f == index[6:0] ? tag_0_95 : _GEN_94; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_96 = 7'h60 == index[6:0] ? tag_0_96 : _GEN_95; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_97 = 7'h61 == index[6:0] ? tag_0_97 : _GEN_96; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_98 = 7'h62 == index[6:0] ? tag_0_98 : _GEN_97; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_99 = 7'h63 == index[6:0] ? tag_0_99 : _GEN_98; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_100 = 7'h64 == index[6:0] ? tag_0_100 : _GEN_99; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_101 = 7'h65 == index[6:0] ? tag_0_101 : _GEN_100; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_102 = 7'h66 == index[6:0] ? tag_0_102 : _GEN_101; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_103 = 7'h67 == index[6:0] ? tag_0_103 : _GEN_102; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_104 = 7'h68 == index[6:0] ? tag_0_104 : _GEN_103; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_105 = 7'h69 == index[6:0] ? tag_0_105 : _GEN_104; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_106 = 7'h6a == index[6:0] ? tag_0_106 : _GEN_105; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_107 = 7'h6b == index[6:0] ? tag_0_107 : _GEN_106; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_108 = 7'h6c == index[6:0] ? tag_0_108 : _GEN_107; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_109 = 7'h6d == index[6:0] ? tag_0_109 : _GEN_108; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_110 = 7'h6e == index[6:0] ? tag_0_110 : _GEN_109; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_111 = 7'h6f == index[6:0] ? tag_0_111 : _GEN_110; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_112 = 7'h70 == index[6:0] ? tag_0_112 : _GEN_111; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_113 = 7'h71 == index[6:0] ? tag_0_113 : _GEN_112; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_114 = 7'h72 == index[6:0] ? tag_0_114 : _GEN_113; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_115 = 7'h73 == index[6:0] ? tag_0_115 : _GEN_114; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_116 = 7'h74 == index[6:0] ? tag_0_116 : _GEN_115; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_117 = 7'h75 == index[6:0] ? tag_0_117 : _GEN_116; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_118 = 7'h76 == index[6:0] ? tag_0_118 : _GEN_117; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_119 = 7'h77 == index[6:0] ? tag_0_119 : _GEN_118; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_120 = 7'h78 == index[6:0] ? tag_0_120 : _GEN_119; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_121 = 7'h79 == index[6:0] ? tag_0_121 : _GEN_120; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_122 = 7'h7a == index[6:0] ? tag_0_122 : _GEN_121; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_123 = 7'h7b == index[6:0] ? tag_0_123 : _GEN_122; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_124 = 7'h7c == index[6:0] ? tag_0_124 : _GEN_123; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_125 = 7'h7d == index[6:0] ? tag_0_125 : _GEN_124; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_126 = 7'h7e == index[6:0] ? tag_0_126 : _GEN_125; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_127 = 7'h7f == index[6:0] ? tag_0_127 : _GEN_126; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_18465 = {{10'd0}, tag}; // @[d_cache.scala 57:24]
  wire  _GEN_129 = 7'h1 == index[6:0] ? valid_0_1 : valid_0_0; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_130 = 7'h2 == index[6:0] ? valid_0_2 : _GEN_129; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_131 = 7'h3 == index[6:0] ? valid_0_3 : _GEN_130; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_132 = 7'h4 == index[6:0] ? valid_0_4 : _GEN_131; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_133 = 7'h5 == index[6:0] ? valid_0_5 : _GEN_132; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_134 = 7'h6 == index[6:0] ? valid_0_6 : _GEN_133; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_135 = 7'h7 == index[6:0] ? valid_0_7 : _GEN_134; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_136 = 7'h8 == index[6:0] ? valid_0_8 : _GEN_135; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_137 = 7'h9 == index[6:0] ? valid_0_9 : _GEN_136; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_138 = 7'ha == index[6:0] ? valid_0_10 : _GEN_137; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_139 = 7'hb == index[6:0] ? valid_0_11 : _GEN_138; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_140 = 7'hc == index[6:0] ? valid_0_12 : _GEN_139; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_141 = 7'hd == index[6:0] ? valid_0_13 : _GEN_140; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_142 = 7'he == index[6:0] ? valid_0_14 : _GEN_141; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_143 = 7'hf == index[6:0] ? valid_0_15 : _GEN_142; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_144 = 7'h10 == index[6:0] ? valid_0_16 : _GEN_143; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_145 = 7'h11 == index[6:0] ? valid_0_17 : _GEN_144; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_146 = 7'h12 == index[6:0] ? valid_0_18 : _GEN_145; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_147 = 7'h13 == index[6:0] ? valid_0_19 : _GEN_146; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_148 = 7'h14 == index[6:0] ? valid_0_20 : _GEN_147; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_149 = 7'h15 == index[6:0] ? valid_0_21 : _GEN_148; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_150 = 7'h16 == index[6:0] ? valid_0_22 : _GEN_149; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_151 = 7'h17 == index[6:0] ? valid_0_23 : _GEN_150; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_152 = 7'h18 == index[6:0] ? valid_0_24 : _GEN_151; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_153 = 7'h19 == index[6:0] ? valid_0_25 : _GEN_152; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_154 = 7'h1a == index[6:0] ? valid_0_26 : _GEN_153; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_155 = 7'h1b == index[6:0] ? valid_0_27 : _GEN_154; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_156 = 7'h1c == index[6:0] ? valid_0_28 : _GEN_155; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_157 = 7'h1d == index[6:0] ? valid_0_29 : _GEN_156; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_158 = 7'h1e == index[6:0] ? valid_0_30 : _GEN_157; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_159 = 7'h1f == index[6:0] ? valid_0_31 : _GEN_158; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_160 = 7'h20 == index[6:0] ? valid_0_32 : _GEN_159; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_161 = 7'h21 == index[6:0] ? valid_0_33 : _GEN_160; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_162 = 7'h22 == index[6:0] ? valid_0_34 : _GEN_161; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_163 = 7'h23 == index[6:0] ? valid_0_35 : _GEN_162; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_164 = 7'h24 == index[6:0] ? valid_0_36 : _GEN_163; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_165 = 7'h25 == index[6:0] ? valid_0_37 : _GEN_164; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_166 = 7'h26 == index[6:0] ? valid_0_38 : _GEN_165; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_167 = 7'h27 == index[6:0] ? valid_0_39 : _GEN_166; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_168 = 7'h28 == index[6:0] ? valid_0_40 : _GEN_167; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_169 = 7'h29 == index[6:0] ? valid_0_41 : _GEN_168; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_170 = 7'h2a == index[6:0] ? valid_0_42 : _GEN_169; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_171 = 7'h2b == index[6:0] ? valid_0_43 : _GEN_170; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_172 = 7'h2c == index[6:0] ? valid_0_44 : _GEN_171; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_173 = 7'h2d == index[6:0] ? valid_0_45 : _GEN_172; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_174 = 7'h2e == index[6:0] ? valid_0_46 : _GEN_173; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_175 = 7'h2f == index[6:0] ? valid_0_47 : _GEN_174; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_176 = 7'h30 == index[6:0] ? valid_0_48 : _GEN_175; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_177 = 7'h31 == index[6:0] ? valid_0_49 : _GEN_176; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_178 = 7'h32 == index[6:0] ? valid_0_50 : _GEN_177; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_179 = 7'h33 == index[6:0] ? valid_0_51 : _GEN_178; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_180 = 7'h34 == index[6:0] ? valid_0_52 : _GEN_179; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_181 = 7'h35 == index[6:0] ? valid_0_53 : _GEN_180; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_182 = 7'h36 == index[6:0] ? valid_0_54 : _GEN_181; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_183 = 7'h37 == index[6:0] ? valid_0_55 : _GEN_182; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_184 = 7'h38 == index[6:0] ? valid_0_56 : _GEN_183; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_185 = 7'h39 == index[6:0] ? valid_0_57 : _GEN_184; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_186 = 7'h3a == index[6:0] ? valid_0_58 : _GEN_185; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_187 = 7'h3b == index[6:0] ? valid_0_59 : _GEN_186; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_188 = 7'h3c == index[6:0] ? valid_0_60 : _GEN_187; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_189 = 7'h3d == index[6:0] ? valid_0_61 : _GEN_188; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_190 = 7'h3e == index[6:0] ? valid_0_62 : _GEN_189; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_191 = 7'h3f == index[6:0] ? valid_0_63 : _GEN_190; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_192 = 7'h40 == index[6:0] ? valid_0_64 : _GEN_191; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_193 = 7'h41 == index[6:0] ? valid_0_65 : _GEN_192; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_194 = 7'h42 == index[6:0] ? valid_0_66 : _GEN_193; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_195 = 7'h43 == index[6:0] ? valid_0_67 : _GEN_194; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_196 = 7'h44 == index[6:0] ? valid_0_68 : _GEN_195; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_197 = 7'h45 == index[6:0] ? valid_0_69 : _GEN_196; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_198 = 7'h46 == index[6:0] ? valid_0_70 : _GEN_197; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_199 = 7'h47 == index[6:0] ? valid_0_71 : _GEN_198; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_200 = 7'h48 == index[6:0] ? valid_0_72 : _GEN_199; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_201 = 7'h49 == index[6:0] ? valid_0_73 : _GEN_200; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_202 = 7'h4a == index[6:0] ? valid_0_74 : _GEN_201; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_203 = 7'h4b == index[6:0] ? valid_0_75 : _GEN_202; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_204 = 7'h4c == index[6:0] ? valid_0_76 : _GEN_203; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_205 = 7'h4d == index[6:0] ? valid_0_77 : _GEN_204; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_206 = 7'h4e == index[6:0] ? valid_0_78 : _GEN_205; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_207 = 7'h4f == index[6:0] ? valid_0_79 : _GEN_206; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_208 = 7'h50 == index[6:0] ? valid_0_80 : _GEN_207; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_209 = 7'h51 == index[6:0] ? valid_0_81 : _GEN_208; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_210 = 7'h52 == index[6:0] ? valid_0_82 : _GEN_209; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_211 = 7'h53 == index[6:0] ? valid_0_83 : _GEN_210; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_212 = 7'h54 == index[6:0] ? valid_0_84 : _GEN_211; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_213 = 7'h55 == index[6:0] ? valid_0_85 : _GEN_212; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_214 = 7'h56 == index[6:0] ? valid_0_86 : _GEN_213; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_215 = 7'h57 == index[6:0] ? valid_0_87 : _GEN_214; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_216 = 7'h58 == index[6:0] ? valid_0_88 : _GEN_215; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_217 = 7'h59 == index[6:0] ? valid_0_89 : _GEN_216; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_218 = 7'h5a == index[6:0] ? valid_0_90 : _GEN_217; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_219 = 7'h5b == index[6:0] ? valid_0_91 : _GEN_218; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_220 = 7'h5c == index[6:0] ? valid_0_92 : _GEN_219; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_221 = 7'h5d == index[6:0] ? valid_0_93 : _GEN_220; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_222 = 7'h5e == index[6:0] ? valid_0_94 : _GEN_221; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_223 = 7'h5f == index[6:0] ? valid_0_95 : _GEN_222; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_224 = 7'h60 == index[6:0] ? valid_0_96 : _GEN_223; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_225 = 7'h61 == index[6:0] ? valid_0_97 : _GEN_224; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_226 = 7'h62 == index[6:0] ? valid_0_98 : _GEN_225; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_227 = 7'h63 == index[6:0] ? valid_0_99 : _GEN_226; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_228 = 7'h64 == index[6:0] ? valid_0_100 : _GEN_227; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_229 = 7'h65 == index[6:0] ? valid_0_101 : _GEN_228; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_230 = 7'h66 == index[6:0] ? valid_0_102 : _GEN_229; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_231 = 7'h67 == index[6:0] ? valid_0_103 : _GEN_230; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_232 = 7'h68 == index[6:0] ? valid_0_104 : _GEN_231; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_233 = 7'h69 == index[6:0] ? valid_0_105 : _GEN_232; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_234 = 7'h6a == index[6:0] ? valid_0_106 : _GEN_233; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_235 = 7'h6b == index[6:0] ? valid_0_107 : _GEN_234; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_236 = 7'h6c == index[6:0] ? valid_0_108 : _GEN_235; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_237 = 7'h6d == index[6:0] ? valid_0_109 : _GEN_236; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_238 = 7'h6e == index[6:0] ? valid_0_110 : _GEN_237; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_239 = 7'h6f == index[6:0] ? valid_0_111 : _GEN_238; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_240 = 7'h70 == index[6:0] ? valid_0_112 : _GEN_239; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_241 = 7'h71 == index[6:0] ? valid_0_113 : _GEN_240; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_242 = 7'h72 == index[6:0] ? valid_0_114 : _GEN_241; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_243 = 7'h73 == index[6:0] ? valid_0_115 : _GEN_242; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_244 = 7'h74 == index[6:0] ? valid_0_116 : _GEN_243; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_245 = 7'h75 == index[6:0] ? valid_0_117 : _GEN_244; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_246 = 7'h76 == index[6:0] ? valid_0_118 : _GEN_245; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_247 = 7'h77 == index[6:0] ? valid_0_119 : _GEN_246; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_248 = 7'h78 == index[6:0] ? valid_0_120 : _GEN_247; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_249 = 7'h79 == index[6:0] ? valid_0_121 : _GEN_248; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_250 = 7'h7a == index[6:0] ? valid_0_122 : _GEN_249; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_251 = 7'h7b == index[6:0] ? valid_0_123 : _GEN_250; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_252 = 7'h7c == index[6:0] ? valid_0_124 : _GEN_251; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_253 = 7'h7d == index[6:0] ? valid_0_125 : _GEN_252; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_254 = 7'h7e == index[6:0] ? valid_0_126 : _GEN_253; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_255 = 7'h7f == index[6:0] ? valid_0_127 : _GEN_254; // @[d_cache.scala 57:{50,50}]
  wire  _T_6 = _GEN_127 == _GEN_18465 & _GEN_255; // @[d_cache.scala 57:33]
  wire [31:0] _GEN_258 = 7'h1 == index[6:0] ? tag_1_1 : tag_1_0; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_259 = 7'h2 == index[6:0] ? tag_1_2 : _GEN_258; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_260 = 7'h3 == index[6:0] ? tag_1_3 : _GEN_259; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_261 = 7'h4 == index[6:0] ? tag_1_4 : _GEN_260; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_262 = 7'h5 == index[6:0] ? tag_1_5 : _GEN_261; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_263 = 7'h6 == index[6:0] ? tag_1_6 : _GEN_262; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_264 = 7'h7 == index[6:0] ? tag_1_7 : _GEN_263; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_265 = 7'h8 == index[6:0] ? tag_1_8 : _GEN_264; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_266 = 7'h9 == index[6:0] ? tag_1_9 : _GEN_265; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_267 = 7'ha == index[6:0] ? tag_1_10 : _GEN_266; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_268 = 7'hb == index[6:0] ? tag_1_11 : _GEN_267; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_269 = 7'hc == index[6:0] ? tag_1_12 : _GEN_268; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_270 = 7'hd == index[6:0] ? tag_1_13 : _GEN_269; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_271 = 7'he == index[6:0] ? tag_1_14 : _GEN_270; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_272 = 7'hf == index[6:0] ? tag_1_15 : _GEN_271; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_273 = 7'h10 == index[6:0] ? tag_1_16 : _GEN_272; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_274 = 7'h11 == index[6:0] ? tag_1_17 : _GEN_273; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_275 = 7'h12 == index[6:0] ? tag_1_18 : _GEN_274; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_276 = 7'h13 == index[6:0] ? tag_1_19 : _GEN_275; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_277 = 7'h14 == index[6:0] ? tag_1_20 : _GEN_276; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_278 = 7'h15 == index[6:0] ? tag_1_21 : _GEN_277; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_279 = 7'h16 == index[6:0] ? tag_1_22 : _GEN_278; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_280 = 7'h17 == index[6:0] ? tag_1_23 : _GEN_279; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_281 = 7'h18 == index[6:0] ? tag_1_24 : _GEN_280; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_282 = 7'h19 == index[6:0] ? tag_1_25 : _GEN_281; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_283 = 7'h1a == index[6:0] ? tag_1_26 : _GEN_282; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_284 = 7'h1b == index[6:0] ? tag_1_27 : _GEN_283; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_285 = 7'h1c == index[6:0] ? tag_1_28 : _GEN_284; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_286 = 7'h1d == index[6:0] ? tag_1_29 : _GEN_285; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_287 = 7'h1e == index[6:0] ? tag_1_30 : _GEN_286; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_288 = 7'h1f == index[6:0] ? tag_1_31 : _GEN_287; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_289 = 7'h20 == index[6:0] ? tag_1_32 : _GEN_288; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_290 = 7'h21 == index[6:0] ? tag_1_33 : _GEN_289; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_291 = 7'h22 == index[6:0] ? tag_1_34 : _GEN_290; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_292 = 7'h23 == index[6:0] ? tag_1_35 : _GEN_291; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_293 = 7'h24 == index[6:0] ? tag_1_36 : _GEN_292; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_294 = 7'h25 == index[6:0] ? tag_1_37 : _GEN_293; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_295 = 7'h26 == index[6:0] ? tag_1_38 : _GEN_294; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_296 = 7'h27 == index[6:0] ? tag_1_39 : _GEN_295; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_297 = 7'h28 == index[6:0] ? tag_1_40 : _GEN_296; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_298 = 7'h29 == index[6:0] ? tag_1_41 : _GEN_297; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_299 = 7'h2a == index[6:0] ? tag_1_42 : _GEN_298; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_300 = 7'h2b == index[6:0] ? tag_1_43 : _GEN_299; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_301 = 7'h2c == index[6:0] ? tag_1_44 : _GEN_300; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_302 = 7'h2d == index[6:0] ? tag_1_45 : _GEN_301; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_303 = 7'h2e == index[6:0] ? tag_1_46 : _GEN_302; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_304 = 7'h2f == index[6:0] ? tag_1_47 : _GEN_303; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_305 = 7'h30 == index[6:0] ? tag_1_48 : _GEN_304; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_306 = 7'h31 == index[6:0] ? tag_1_49 : _GEN_305; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_307 = 7'h32 == index[6:0] ? tag_1_50 : _GEN_306; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_308 = 7'h33 == index[6:0] ? tag_1_51 : _GEN_307; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_309 = 7'h34 == index[6:0] ? tag_1_52 : _GEN_308; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_310 = 7'h35 == index[6:0] ? tag_1_53 : _GEN_309; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_311 = 7'h36 == index[6:0] ? tag_1_54 : _GEN_310; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_312 = 7'h37 == index[6:0] ? tag_1_55 : _GEN_311; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_313 = 7'h38 == index[6:0] ? tag_1_56 : _GEN_312; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_314 = 7'h39 == index[6:0] ? tag_1_57 : _GEN_313; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_315 = 7'h3a == index[6:0] ? tag_1_58 : _GEN_314; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_316 = 7'h3b == index[6:0] ? tag_1_59 : _GEN_315; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_317 = 7'h3c == index[6:0] ? tag_1_60 : _GEN_316; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_318 = 7'h3d == index[6:0] ? tag_1_61 : _GEN_317; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_319 = 7'h3e == index[6:0] ? tag_1_62 : _GEN_318; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_320 = 7'h3f == index[6:0] ? tag_1_63 : _GEN_319; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_321 = 7'h40 == index[6:0] ? tag_1_64 : _GEN_320; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_322 = 7'h41 == index[6:0] ? tag_1_65 : _GEN_321; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_323 = 7'h42 == index[6:0] ? tag_1_66 : _GEN_322; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_324 = 7'h43 == index[6:0] ? tag_1_67 : _GEN_323; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_325 = 7'h44 == index[6:0] ? tag_1_68 : _GEN_324; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_326 = 7'h45 == index[6:0] ? tag_1_69 : _GEN_325; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_327 = 7'h46 == index[6:0] ? tag_1_70 : _GEN_326; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_328 = 7'h47 == index[6:0] ? tag_1_71 : _GEN_327; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_329 = 7'h48 == index[6:0] ? tag_1_72 : _GEN_328; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_330 = 7'h49 == index[6:0] ? tag_1_73 : _GEN_329; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_331 = 7'h4a == index[6:0] ? tag_1_74 : _GEN_330; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_332 = 7'h4b == index[6:0] ? tag_1_75 : _GEN_331; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_333 = 7'h4c == index[6:0] ? tag_1_76 : _GEN_332; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_334 = 7'h4d == index[6:0] ? tag_1_77 : _GEN_333; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_335 = 7'h4e == index[6:0] ? tag_1_78 : _GEN_334; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_336 = 7'h4f == index[6:0] ? tag_1_79 : _GEN_335; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_337 = 7'h50 == index[6:0] ? tag_1_80 : _GEN_336; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_338 = 7'h51 == index[6:0] ? tag_1_81 : _GEN_337; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_339 = 7'h52 == index[6:0] ? tag_1_82 : _GEN_338; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_340 = 7'h53 == index[6:0] ? tag_1_83 : _GEN_339; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_341 = 7'h54 == index[6:0] ? tag_1_84 : _GEN_340; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_342 = 7'h55 == index[6:0] ? tag_1_85 : _GEN_341; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_343 = 7'h56 == index[6:0] ? tag_1_86 : _GEN_342; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_344 = 7'h57 == index[6:0] ? tag_1_87 : _GEN_343; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_345 = 7'h58 == index[6:0] ? tag_1_88 : _GEN_344; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_346 = 7'h59 == index[6:0] ? tag_1_89 : _GEN_345; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_347 = 7'h5a == index[6:0] ? tag_1_90 : _GEN_346; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_348 = 7'h5b == index[6:0] ? tag_1_91 : _GEN_347; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_349 = 7'h5c == index[6:0] ? tag_1_92 : _GEN_348; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_350 = 7'h5d == index[6:0] ? tag_1_93 : _GEN_349; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_351 = 7'h5e == index[6:0] ? tag_1_94 : _GEN_350; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_352 = 7'h5f == index[6:0] ? tag_1_95 : _GEN_351; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_353 = 7'h60 == index[6:0] ? tag_1_96 : _GEN_352; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_354 = 7'h61 == index[6:0] ? tag_1_97 : _GEN_353; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_355 = 7'h62 == index[6:0] ? tag_1_98 : _GEN_354; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_356 = 7'h63 == index[6:0] ? tag_1_99 : _GEN_355; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_357 = 7'h64 == index[6:0] ? tag_1_100 : _GEN_356; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_358 = 7'h65 == index[6:0] ? tag_1_101 : _GEN_357; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_359 = 7'h66 == index[6:0] ? tag_1_102 : _GEN_358; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_360 = 7'h67 == index[6:0] ? tag_1_103 : _GEN_359; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_361 = 7'h68 == index[6:0] ? tag_1_104 : _GEN_360; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_362 = 7'h69 == index[6:0] ? tag_1_105 : _GEN_361; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_363 = 7'h6a == index[6:0] ? tag_1_106 : _GEN_362; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_364 = 7'h6b == index[6:0] ? tag_1_107 : _GEN_363; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_365 = 7'h6c == index[6:0] ? tag_1_108 : _GEN_364; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_366 = 7'h6d == index[6:0] ? tag_1_109 : _GEN_365; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_367 = 7'h6e == index[6:0] ? tag_1_110 : _GEN_366; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_368 = 7'h6f == index[6:0] ? tag_1_111 : _GEN_367; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_369 = 7'h70 == index[6:0] ? tag_1_112 : _GEN_368; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_370 = 7'h71 == index[6:0] ? tag_1_113 : _GEN_369; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_371 = 7'h72 == index[6:0] ? tag_1_114 : _GEN_370; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_372 = 7'h73 == index[6:0] ? tag_1_115 : _GEN_371; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_373 = 7'h74 == index[6:0] ? tag_1_116 : _GEN_372; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_374 = 7'h75 == index[6:0] ? tag_1_117 : _GEN_373; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_375 = 7'h76 == index[6:0] ? tag_1_118 : _GEN_374; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_376 = 7'h77 == index[6:0] ? tag_1_119 : _GEN_375; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_377 = 7'h78 == index[6:0] ? tag_1_120 : _GEN_376; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_378 = 7'h79 == index[6:0] ? tag_1_121 : _GEN_377; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_379 = 7'h7a == index[6:0] ? tag_1_122 : _GEN_378; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_380 = 7'h7b == index[6:0] ? tag_1_123 : _GEN_379; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_381 = 7'h7c == index[6:0] ? tag_1_124 : _GEN_380; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_382 = 7'h7d == index[6:0] ? tag_1_125 : _GEN_381; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_383 = 7'h7e == index[6:0] ? tag_1_126 : _GEN_382; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_384 = 7'h7f == index[6:0] ? tag_1_127 : _GEN_383; // @[d_cache.scala 62:{24,24}]
  wire  _GEN_386 = 7'h1 == index[6:0] ? valid_1_1 : valid_1_0; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_387 = 7'h2 == index[6:0] ? valid_1_2 : _GEN_386; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_388 = 7'h3 == index[6:0] ? valid_1_3 : _GEN_387; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_389 = 7'h4 == index[6:0] ? valid_1_4 : _GEN_388; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_390 = 7'h5 == index[6:0] ? valid_1_5 : _GEN_389; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_391 = 7'h6 == index[6:0] ? valid_1_6 : _GEN_390; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_392 = 7'h7 == index[6:0] ? valid_1_7 : _GEN_391; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_393 = 7'h8 == index[6:0] ? valid_1_8 : _GEN_392; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_394 = 7'h9 == index[6:0] ? valid_1_9 : _GEN_393; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_395 = 7'ha == index[6:0] ? valid_1_10 : _GEN_394; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_396 = 7'hb == index[6:0] ? valid_1_11 : _GEN_395; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_397 = 7'hc == index[6:0] ? valid_1_12 : _GEN_396; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_398 = 7'hd == index[6:0] ? valid_1_13 : _GEN_397; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_399 = 7'he == index[6:0] ? valid_1_14 : _GEN_398; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_400 = 7'hf == index[6:0] ? valid_1_15 : _GEN_399; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_401 = 7'h10 == index[6:0] ? valid_1_16 : _GEN_400; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_402 = 7'h11 == index[6:0] ? valid_1_17 : _GEN_401; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_403 = 7'h12 == index[6:0] ? valid_1_18 : _GEN_402; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_404 = 7'h13 == index[6:0] ? valid_1_19 : _GEN_403; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_405 = 7'h14 == index[6:0] ? valid_1_20 : _GEN_404; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_406 = 7'h15 == index[6:0] ? valid_1_21 : _GEN_405; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_407 = 7'h16 == index[6:0] ? valid_1_22 : _GEN_406; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_408 = 7'h17 == index[6:0] ? valid_1_23 : _GEN_407; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_409 = 7'h18 == index[6:0] ? valid_1_24 : _GEN_408; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_410 = 7'h19 == index[6:0] ? valid_1_25 : _GEN_409; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_411 = 7'h1a == index[6:0] ? valid_1_26 : _GEN_410; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_412 = 7'h1b == index[6:0] ? valid_1_27 : _GEN_411; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_413 = 7'h1c == index[6:0] ? valid_1_28 : _GEN_412; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_414 = 7'h1d == index[6:0] ? valid_1_29 : _GEN_413; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_415 = 7'h1e == index[6:0] ? valid_1_30 : _GEN_414; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_416 = 7'h1f == index[6:0] ? valid_1_31 : _GEN_415; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_417 = 7'h20 == index[6:0] ? valid_1_32 : _GEN_416; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_418 = 7'h21 == index[6:0] ? valid_1_33 : _GEN_417; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_419 = 7'h22 == index[6:0] ? valid_1_34 : _GEN_418; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_420 = 7'h23 == index[6:0] ? valid_1_35 : _GEN_419; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_421 = 7'h24 == index[6:0] ? valid_1_36 : _GEN_420; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_422 = 7'h25 == index[6:0] ? valid_1_37 : _GEN_421; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_423 = 7'h26 == index[6:0] ? valid_1_38 : _GEN_422; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_424 = 7'h27 == index[6:0] ? valid_1_39 : _GEN_423; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_425 = 7'h28 == index[6:0] ? valid_1_40 : _GEN_424; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_426 = 7'h29 == index[6:0] ? valid_1_41 : _GEN_425; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_427 = 7'h2a == index[6:0] ? valid_1_42 : _GEN_426; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_428 = 7'h2b == index[6:0] ? valid_1_43 : _GEN_427; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_429 = 7'h2c == index[6:0] ? valid_1_44 : _GEN_428; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_430 = 7'h2d == index[6:0] ? valid_1_45 : _GEN_429; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_431 = 7'h2e == index[6:0] ? valid_1_46 : _GEN_430; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_432 = 7'h2f == index[6:0] ? valid_1_47 : _GEN_431; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_433 = 7'h30 == index[6:0] ? valid_1_48 : _GEN_432; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_434 = 7'h31 == index[6:0] ? valid_1_49 : _GEN_433; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_435 = 7'h32 == index[6:0] ? valid_1_50 : _GEN_434; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_436 = 7'h33 == index[6:0] ? valid_1_51 : _GEN_435; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_437 = 7'h34 == index[6:0] ? valid_1_52 : _GEN_436; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_438 = 7'h35 == index[6:0] ? valid_1_53 : _GEN_437; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_439 = 7'h36 == index[6:0] ? valid_1_54 : _GEN_438; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_440 = 7'h37 == index[6:0] ? valid_1_55 : _GEN_439; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_441 = 7'h38 == index[6:0] ? valid_1_56 : _GEN_440; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_442 = 7'h39 == index[6:0] ? valid_1_57 : _GEN_441; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_443 = 7'h3a == index[6:0] ? valid_1_58 : _GEN_442; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_444 = 7'h3b == index[6:0] ? valid_1_59 : _GEN_443; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_445 = 7'h3c == index[6:0] ? valid_1_60 : _GEN_444; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_446 = 7'h3d == index[6:0] ? valid_1_61 : _GEN_445; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_447 = 7'h3e == index[6:0] ? valid_1_62 : _GEN_446; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_448 = 7'h3f == index[6:0] ? valid_1_63 : _GEN_447; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_449 = 7'h40 == index[6:0] ? valid_1_64 : _GEN_448; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_450 = 7'h41 == index[6:0] ? valid_1_65 : _GEN_449; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_451 = 7'h42 == index[6:0] ? valid_1_66 : _GEN_450; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_452 = 7'h43 == index[6:0] ? valid_1_67 : _GEN_451; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_453 = 7'h44 == index[6:0] ? valid_1_68 : _GEN_452; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_454 = 7'h45 == index[6:0] ? valid_1_69 : _GEN_453; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_455 = 7'h46 == index[6:0] ? valid_1_70 : _GEN_454; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_456 = 7'h47 == index[6:0] ? valid_1_71 : _GEN_455; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_457 = 7'h48 == index[6:0] ? valid_1_72 : _GEN_456; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_458 = 7'h49 == index[6:0] ? valid_1_73 : _GEN_457; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_459 = 7'h4a == index[6:0] ? valid_1_74 : _GEN_458; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_460 = 7'h4b == index[6:0] ? valid_1_75 : _GEN_459; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_461 = 7'h4c == index[6:0] ? valid_1_76 : _GEN_460; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_462 = 7'h4d == index[6:0] ? valid_1_77 : _GEN_461; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_463 = 7'h4e == index[6:0] ? valid_1_78 : _GEN_462; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_464 = 7'h4f == index[6:0] ? valid_1_79 : _GEN_463; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_465 = 7'h50 == index[6:0] ? valid_1_80 : _GEN_464; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_466 = 7'h51 == index[6:0] ? valid_1_81 : _GEN_465; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_467 = 7'h52 == index[6:0] ? valid_1_82 : _GEN_466; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_468 = 7'h53 == index[6:0] ? valid_1_83 : _GEN_467; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_469 = 7'h54 == index[6:0] ? valid_1_84 : _GEN_468; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_470 = 7'h55 == index[6:0] ? valid_1_85 : _GEN_469; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_471 = 7'h56 == index[6:0] ? valid_1_86 : _GEN_470; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_472 = 7'h57 == index[6:0] ? valid_1_87 : _GEN_471; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_473 = 7'h58 == index[6:0] ? valid_1_88 : _GEN_472; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_474 = 7'h59 == index[6:0] ? valid_1_89 : _GEN_473; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_475 = 7'h5a == index[6:0] ? valid_1_90 : _GEN_474; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_476 = 7'h5b == index[6:0] ? valid_1_91 : _GEN_475; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_477 = 7'h5c == index[6:0] ? valid_1_92 : _GEN_476; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_478 = 7'h5d == index[6:0] ? valid_1_93 : _GEN_477; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_479 = 7'h5e == index[6:0] ? valid_1_94 : _GEN_478; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_480 = 7'h5f == index[6:0] ? valid_1_95 : _GEN_479; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_481 = 7'h60 == index[6:0] ? valid_1_96 : _GEN_480; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_482 = 7'h61 == index[6:0] ? valid_1_97 : _GEN_481; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_483 = 7'h62 == index[6:0] ? valid_1_98 : _GEN_482; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_484 = 7'h63 == index[6:0] ? valid_1_99 : _GEN_483; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_485 = 7'h64 == index[6:0] ? valid_1_100 : _GEN_484; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_486 = 7'h65 == index[6:0] ? valid_1_101 : _GEN_485; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_487 = 7'h66 == index[6:0] ? valid_1_102 : _GEN_486; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_488 = 7'h67 == index[6:0] ? valid_1_103 : _GEN_487; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_489 = 7'h68 == index[6:0] ? valid_1_104 : _GEN_488; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_490 = 7'h69 == index[6:0] ? valid_1_105 : _GEN_489; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_491 = 7'h6a == index[6:0] ? valid_1_106 : _GEN_490; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_492 = 7'h6b == index[6:0] ? valid_1_107 : _GEN_491; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_493 = 7'h6c == index[6:0] ? valid_1_108 : _GEN_492; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_494 = 7'h6d == index[6:0] ? valid_1_109 : _GEN_493; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_495 = 7'h6e == index[6:0] ? valid_1_110 : _GEN_494; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_496 = 7'h6f == index[6:0] ? valid_1_111 : _GEN_495; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_497 = 7'h70 == index[6:0] ? valid_1_112 : _GEN_496; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_498 = 7'h71 == index[6:0] ? valid_1_113 : _GEN_497; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_499 = 7'h72 == index[6:0] ? valid_1_114 : _GEN_498; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_500 = 7'h73 == index[6:0] ? valid_1_115 : _GEN_499; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_501 = 7'h74 == index[6:0] ? valid_1_116 : _GEN_500; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_502 = 7'h75 == index[6:0] ? valid_1_117 : _GEN_501; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_503 = 7'h76 == index[6:0] ? valid_1_118 : _GEN_502; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_504 = 7'h77 == index[6:0] ? valid_1_119 : _GEN_503; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_505 = 7'h78 == index[6:0] ? valid_1_120 : _GEN_504; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_506 = 7'h79 == index[6:0] ? valid_1_121 : _GEN_505; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_507 = 7'h7a == index[6:0] ? valid_1_122 : _GEN_506; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_508 = 7'h7b == index[6:0] ? valid_1_123 : _GEN_507; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_509 = 7'h7c == index[6:0] ? valid_1_124 : _GEN_508; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_510 = 7'h7d == index[6:0] ? valid_1_125 : _GEN_509; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_511 = 7'h7e == index[6:0] ? valid_1_126 : _GEN_510; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_512 = 7'h7f == index[6:0] ? valid_1_127 : _GEN_511; // @[d_cache.scala 62:{50,50}]
  wire  _T_11 = _GEN_384 == _GEN_18465 & _GEN_512; // @[d_cache.scala 62:33]
  reg [2:0] state; // @[d_cache.scala 76:24]
  wire  _T_20 = 3'h0 == state; // @[d_cache.scala 81:18]
  wire  _T_21 = 3'h1 == state; // @[d_cache.scala 81:18]
  wire  _GEN_775 = 7'h1 == index[6:0] ? dirty_0_1 : dirty_0_0; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_776 = 7'h2 == index[6:0] ? dirty_0_2 : _GEN_775; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_777 = 7'h3 == index[6:0] ? dirty_0_3 : _GEN_776; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_778 = 7'h4 == index[6:0] ? dirty_0_4 : _GEN_777; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_779 = 7'h5 == index[6:0] ? dirty_0_5 : _GEN_778; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_780 = 7'h6 == index[6:0] ? dirty_0_6 : _GEN_779; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_781 = 7'h7 == index[6:0] ? dirty_0_7 : _GEN_780; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_782 = 7'h8 == index[6:0] ? dirty_0_8 : _GEN_781; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_783 = 7'h9 == index[6:0] ? dirty_0_9 : _GEN_782; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_784 = 7'ha == index[6:0] ? dirty_0_10 : _GEN_783; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_785 = 7'hb == index[6:0] ? dirty_0_11 : _GEN_784; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_786 = 7'hc == index[6:0] ? dirty_0_12 : _GEN_785; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_787 = 7'hd == index[6:0] ? dirty_0_13 : _GEN_786; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_788 = 7'he == index[6:0] ? dirty_0_14 : _GEN_787; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_789 = 7'hf == index[6:0] ? dirty_0_15 : _GEN_788; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_790 = 7'h10 == index[6:0] ? dirty_0_16 : _GEN_789; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_791 = 7'h11 == index[6:0] ? dirty_0_17 : _GEN_790; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_792 = 7'h12 == index[6:0] ? dirty_0_18 : _GEN_791; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_793 = 7'h13 == index[6:0] ? dirty_0_19 : _GEN_792; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_794 = 7'h14 == index[6:0] ? dirty_0_20 : _GEN_793; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_795 = 7'h15 == index[6:0] ? dirty_0_21 : _GEN_794; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_796 = 7'h16 == index[6:0] ? dirty_0_22 : _GEN_795; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_797 = 7'h17 == index[6:0] ? dirty_0_23 : _GEN_796; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_798 = 7'h18 == index[6:0] ? dirty_0_24 : _GEN_797; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_799 = 7'h19 == index[6:0] ? dirty_0_25 : _GEN_798; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_800 = 7'h1a == index[6:0] ? dirty_0_26 : _GEN_799; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_801 = 7'h1b == index[6:0] ? dirty_0_27 : _GEN_800; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_802 = 7'h1c == index[6:0] ? dirty_0_28 : _GEN_801; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_803 = 7'h1d == index[6:0] ? dirty_0_29 : _GEN_802; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_804 = 7'h1e == index[6:0] ? dirty_0_30 : _GEN_803; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_805 = 7'h1f == index[6:0] ? dirty_0_31 : _GEN_804; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_806 = 7'h20 == index[6:0] ? dirty_0_32 : _GEN_805; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_807 = 7'h21 == index[6:0] ? dirty_0_33 : _GEN_806; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_808 = 7'h22 == index[6:0] ? dirty_0_34 : _GEN_807; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_809 = 7'h23 == index[6:0] ? dirty_0_35 : _GEN_808; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_810 = 7'h24 == index[6:0] ? dirty_0_36 : _GEN_809; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_811 = 7'h25 == index[6:0] ? dirty_0_37 : _GEN_810; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_812 = 7'h26 == index[6:0] ? dirty_0_38 : _GEN_811; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_813 = 7'h27 == index[6:0] ? dirty_0_39 : _GEN_812; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_814 = 7'h28 == index[6:0] ? dirty_0_40 : _GEN_813; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_815 = 7'h29 == index[6:0] ? dirty_0_41 : _GEN_814; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_816 = 7'h2a == index[6:0] ? dirty_0_42 : _GEN_815; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_817 = 7'h2b == index[6:0] ? dirty_0_43 : _GEN_816; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_818 = 7'h2c == index[6:0] ? dirty_0_44 : _GEN_817; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_819 = 7'h2d == index[6:0] ? dirty_0_45 : _GEN_818; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_820 = 7'h2e == index[6:0] ? dirty_0_46 : _GEN_819; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_821 = 7'h2f == index[6:0] ? dirty_0_47 : _GEN_820; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_822 = 7'h30 == index[6:0] ? dirty_0_48 : _GEN_821; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_823 = 7'h31 == index[6:0] ? dirty_0_49 : _GEN_822; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_824 = 7'h32 == index[6:0] ? dirty_0_50 : _GEN_823; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_825 = 7'h33 == index[6:0] ? dirty_0_51 : _GEN_824; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_826 = 7'h34 == index[6:0] ? dirty_0_52 : _GEN_825; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_827 = 7'h35 == index[6:0] ? dirty_0_53 : _GEN_826; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_828 = 7'h36 == index[6:0] ? dirty_0_54 : _GEN_827; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_829 = 7'h37 == index[6:0] ? dirty_0_55 : _GEN_828; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_830 = 7'h38 == index[6:0] ? dirty_0_56 : _GEN_829; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_831 = 7'h39 == index[6:0] ? dirty_0_57 : _GEN_830; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_832 = 7'h3a == index[6:0] ? dirty_0_58 : _GEN_831; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_833 = 7'h3b == index[6:0] ? dirty_0_59 : _GEN_832; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_834 = 7'h3c == index[6:0] ? dirty_0_60 : _GEN_833; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_835 = 7'h3d == index[6:0] ? dirty_0_61 : _GEN_834; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_836 = 7'h3e == index[6:0] ? dirty_0_62 : _GEN_835; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_837 = 7'h3f == index[6:0] ? dirty_0_63 : _GEN_836; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_838 = 7'h40 == index[6:0] ? dirty_0_64 : _GEN_837; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_839 = 7'h41 == index[6:0] ? dirty_0_65 : _GEN_838; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_840 = 7'h42 == index[6:0] ? dirty_0_66 : _GEN_839; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_841 = 7'h43 == index[6:0] ? dirty_0_67 : _GEN_840; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_842 = 7'h44 == index[6:0] ? dirty_0_68 : _GEN_841; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_843 = 7'h45 == index[6:0] ? dirty_0_69 : _GEN_842; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_844 = 7'h46 == index[6:0] ? dirty_0_70 : _GEN_843; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_845 = 7'h47 == index[6:0] ? dirty_0_71 : _GEN_844; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_846 = 7'h48 == index[6:0] ? dirty_0_72 : _GEN_845; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_847 = 7'h49 == index[6:0] ? dirty_0_73 : _GEN_846; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_848 = 7'h4a == index[6:0] ? dirty_0_74 : _GEN_847; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_849 = 7'h4b == index[6:0] ? dirty_0_75 : _GEN_848; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_850 = 7'h4c == index[6:0] ? dirty_0_76 : _GEN_849; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_851 = 7'h4d == index[6:0] ? dirty_0_77 : _GEN_850; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_852 = 7'h4e == index[6:0] ? dirty_0_78 : _GEN_851; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_853 = 7'h4f == index[6:0] ? dirty_0_79 : _GEN_852; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_854 = 7'h50 == index[6:0] ? dirty_0_80 : _GEN_853; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_855 = 7'h51 == index[6:0] ? dirty_0_81 : _GEN_854; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_856 = 7'h52 == index[6:0] ? dirty_0_82 : _GEN_855; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_857 = 7'h53 == index[6:0] ? dirty_0_83 : _GEN_856; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_858 = 7'h54 == index[6:0] ? dirty_0_84 : _GEN_857; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_859 = 7'h55 == index[6:0] ? dirty_0_85 : _GEN_858; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_860 = 7'h56 == index[6:0] ? dirty_0_86 : _GEN_859; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_861 = 7'h57 == index[6:0] ? dirty_0_87 : _GEN_860; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_862 = 7'h58 == index[6:0] ? dirty_0_88 : _GEN_861; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_863 = 7'h59 == index[6:0] ? dirty_0_89 : _GEN_862; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_864 = 7'h5a == index[6:0] ? dirty_0_90 : _GEN_863; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_865 = 7'h5b == index[6:0] ? dirty_0_91 : _GEN_864; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_866 = 7'h5c == index[6:0] ? dirty_0_92 : _GEN_865; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_867 = 7'h5d == index[6:0] ? dirty_0_93 : _GEN_866; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_868 = 7'h5e == index[6:0] ? dirty_0_94 : _GEN_867; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_869 = 7'h5f == index[6:0] ? dirty_0_95 : _GEN_868; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_870 = 7'h60 == index[6:0] ? dirty_0_96 : _GEN_869; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_871 = 7'h61 == index[6:0] ? dirty_0_97 : _GEN_870; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_872 = 7'h62 == index[6:0] ? dirty_0_98 : _GEN_871; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_873 = 7'h63 == index[6:0] ? dirty_0_99 : _GEN_872; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_874 = 7'h64 == index[6:0] ? dirty_0_100 : _GEN_873; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_875 = 7'h65 == index[6:0] ? dirty_0_101 : _GEN_874; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_876 = 7'h66 == index[6:0] ? dirty_0_102 : _GEN_875; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_877 = 7'h67 == index[6:0] ? dirty_0_103 : _GEN_876; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_878 = 7'h68 == index[6:0] ? dirty_0_104 : _GEN_877; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_879 = 7'h69 == index[6:0] ? dirty_0_105 : _GEN_878; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_880 = 7'h6a == index[6:0] ? dirty_0_106 : _GEN_879; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_881 = 7'h6b == index[6:0] ? dirty_0_107 : _GEN_880; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_882 = 7'h6c == index[6:0] ? dirty_0_108 : _GEN_881; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_883 = 7'h6d == index[6:0] ? dirty_0_109 : _GEN_882; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_884 = 7'h6e == index[6:0] ? dirty_0_110 : _GEN_883; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_885 = 7'h6f == index[6:0] ? dirty_0_111 : _GEN_884; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_886 = 7'h70 == index[6:0] ? dirty_0_112 : _GEN_885; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_887 = 7'h71 == index[6:0] ? dirty_0_113 : _GEN_886; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_888 = 7'h72 == index[6:0] ? dirty_0_114 : _GEN_887; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_889 = 7'h73 == index[6:0] ? dirty_0_115 : _GEN_888; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_890 = 7'h74 == index[6:0] ? dirty_0_116 : _GEN_889; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_891 = 7'h75 == index[6:0] ? dirty_0_117 : _GEN_890; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_892 = 7'h76 == index[6:0] ? dirty_0_118 : _GEN_891; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_893 = 7'h77 == index[6:0] ? dirty_0_119 : _GEN_892; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_894 = 7'h78 == index[6:0] ? dirty_0_120 : _GEN_893; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_895 = 7'h79 == index[6:0] ? dirty_0_121 : _GEN_894; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_896 = 7'h7a == index[6:0] ? dirty_0_122 : _GEN_895; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_897 = 7'h7b == index[6:0] ? dirty_0_123 : _GEN_896; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_898 = 7'h7c == index[6:0] ? dirty_0_124 : _GEN_897; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_899 = 7'h7d == index[6:0] ? dirty_0_125 : _GEN_898; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_900 = 7'h7e == index[6:0] ? dirty_0_126 : _GEN_899; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_901 = 7'h7f == index[6:0] ? dirty_0_127 : _GEN_900; // @[d_cache.scala 93:{27,27}]
  wire [2:0] _GEN_902 = io_from_lsu_rready ? 3'h0 : state; // @[d_cache.scala 76:24 92:41 94:27]
  wire  _GEN_904 = 7'h1 == index[6:0] ? dirty_1_1 : dirty_1_0; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_905 = 7'h2 == index[6:0] ? dirty_1_2 : _GEN_904; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_906 = 7'h3 == index[6:0] ? dirty_1_3 : _GEN_905; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_907 = 7'h4 == index[6:0] ? dirty_1_4 : _GEN_906; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_908 = 7'h5 == index[6:0] ? dirty_1_5 : _GEN_907; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_909 = 7'h6 == index[6:0] ? dirty_1_6 : _GEN_908; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_910 = 7'h7 == index[6:0] ? dirty_1_7 : _GEN_909; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_911 = 7'h8 == index[6:0] ? dirty_1_8 : _GEN_910; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_912 = 7'h9 == index[6:0] ? dirty_1_9 : _GEN_911; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_913 = 7'ha == index[6:0] ? dirty_1_10 : _GEN_912; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_914 = 7'hb == index[6:0] ? dirty_1_11 : _GEN_913; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_915 = 7'hc == index[6:0] ? dirty_1_12 : _GEN_914; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_916 = 7'hd == index[6:0] ? dirty_1_13 : _GEN_915; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_917 = 7'he == index[6:0] ? dirty_1_14 : _GEN_916; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_918 = 7'hf == index[6:0] ? dirty_1_15 : _GEN_917; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_919 = 7'h10 == index[6:0] ? dirty_1_16 : _GEN_918; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_920 = 7'h11 == index[6:0] ? dirty_1_17 : _GEN_919; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_921 = 7'h12 == index[6:0] ? dirty_1_18 : _GEN_920; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_922 = 7'h13 == index[6:0] ? dirty_1_19 : _GEN_921; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_923 = 7'h14 == index[6:0] ? dirty_1_20 : _GEN_922; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_924 = 7'h15 == index[6:0] ? dirty_1_21 : _GEN_923; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_925 = 7'h16 == index[6:0] ? dirty_1_22 : _GEN_924; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_926 = 7'h17 == index[6:0] ? dirty_1_23 : _GEN_925; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_927 = 7'h18 == index[6:0] ? dirty_1_24 : _GEN_926; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_928 = 7'h19 == index[6:0] ? dirty_1_25 : _GEN_927; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_929 = 7'h1a == index[6:0] ? dirty_1_26 : _GEN_928; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_930 = 7'h1b == index[6:0] ? dirty_1_27 : _GEN_929; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_931 = 7'h1c == index[6:0] ? dirty_1_28 : _GEN_930; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_932 = 7'h1d == index[6:0] ? dirty_1_29 : _GEN_931; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_933 = 7'h1e == index[6:0] ? dirty_1_30 : _GEN_932; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_934 = 7'h1f == index[6:0] ? dirty_1_31 : _GEN_933; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_935 = 7'h20 == index[6:0] ? dirty_1_32 : _GEN_934; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_936 = 7'h21 == index[6:0] ? dirty_1_33 : _GEN_935; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_937 = 7'h22 == index[6:0] ? dirty_1_34 : _GEN_936; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_938 = 7'h23 == index[6:0] ? dirty_1_35 : _GEN_937; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_939 = 7'h24 == index[6:0] ? dirty_1_36 : _GEN_938; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_940 = 7'h25 == index[6:0] ? dirty_1_37 : _GEN_939; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_941 = 7'h26 == index[6:0] ? dirty_1_38 : _GEN_940; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_942 = 7'h27 == index[6:0] ? dirty_1_39 : _GEN_941; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_943 = 7'h28 == index[6:0] ? dirty_1_40 : _GEN_942; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_944 = 7'h29 == index[6:0] ? dirty_1_41 : _GEN_943; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_945 = 7'h2a == index[6:0] ? dirty_1_42 : _GEN_944; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_946 = 7'h2b == index[6:0] ? dirty_1_43 : _GEN_945; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_947 = 7'h2c == index[6:0] ? dirty_1_44 : _GEN_946; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_948 = 7'h2d == index[6:0] ? dirty_1_45 : _GEN_947; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_949 = 7'h2e == index[6:0] ? dirty_1_46 : _GEN_948; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_950 = 7'h2f == index[6:0] ? dirty_1_47 : _GEN_949; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_951 = 7'h30 == index[6:0] ? dirty_1_48 : _GEN_950; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_952 = 7'h31 == index[6:0] ? dirty_1_49 : _GEN_951; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_953 = 7'h32 == index[6:0] ? dirty_1_50 : _GEN_952; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_954 = 7'h33 == index[6:0] ? dirty_1_51 : _GEN_953; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_955 = 7'h34 == index[6:0] ? dirty_1_52 : _GEN_954; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_956 = 7'h35 == index[6:0] ? dirty_1_53 : _GEN_955; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_957 = 7'h36 == index[6:0] ? dirty_1_54 : _GEN_956; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_958 = 7'h37 == index[6:0] ? dirty_1_55 : _GEN_957; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_959 = 7'h38 == index[6:0] ? dirty_1_56 : _GEN_958; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_960 = 7'h39 == index[6:0] ? dirty_1_57 : _GEN_959; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_961 = 7'h3a == index[6:0] ? dirty_1_58 : _GEN_960; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_962 = 7'h3b == index[6:0] ? dirty_1_59 : _GEN_961; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_963 = 7'h3c == index[6:0] ? dirty_1_60 : _GEN_962; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_964 = 7'h3d == index[6:0] ? dirty_1_61 : _GEN_963; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_965 = 7'h3e == index[6:0] ? dirty_1_62 : _GEN_964; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_966 = 7'h3f == index[6:0] ? dirty_1_63 : _GEN_965; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_967 = 7'h40 == index[6:0] ? dirty_1_64 : _GEN_966; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_968 = 7'h41 == index[6:0] ? dirty_1_65 : _GEN_967; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_969 = 7'h42 == index[6:0] ? dirty_1_66 : _GEN_968; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_970 = 7'h43 == index[6:0] ? dirty_1_67 : _GEN_969; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_971 = 7'h44 == index[6:0] ? dirty_1_68 : _GEN_970; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_972 = 7'h45 == index[6:0] ? dirty_1_69 : _GEN_971; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_973 = 7'h46 == index[6:0] ? dirty_1_70 : _GEN_972; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_974 = 7'h47 == index[6:0] ? dirty_1_71 : _GEN_973; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_975 = 7'h48 == index[6:0] ? dirty_1_72 : _GEN_974; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_976 = 7'h49 == index[6:0] ? dirty_1_73 : _GEN_975; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_977 = 7'h4a == index[6:0] ? dirty_1_74 : _GEN_976; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_978 = 7'h4b == index[6:0] ? dirty_1_75 : _GEN_977; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_979 = 7'h4c == index[6:0] ? dirty_1_76 : _GEN_978; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_980 = 7'h4d == index[6:0] ? dirty_1_77 : _GEN_979; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_981 = 7'h4e == index[6:0] ? dirty_1_78 : _GEN_980; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_982 = 7'h4f == index[6:0] ? dirty_1_79 : _GEN_981; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_983 = 7'h50 == index[6:0] ? dirty_1_80 : _GEN_982; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_984 = 7'h51 == index[6:0] ? dirty_1_81 : _GEN_983; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_985 = 7'h52 == index[6:0] ? dirty_1_82 : _GEN_984; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_986 = 7'h53 == index[6:0] ? dirty_1_83 : _GEN_985; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_987 = 7'h54 == index[6:0] ? dirty_1_84 : _GEN_986; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_988 = 7'h55 == index[6:0] ? dirty_1_85 : _GEN_987; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_989 = 7'h56 == index[6:0] ? dirty_1_86 : _GEN_988; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_990 = 7'h57 == index[6:0] ? dirty_1_87 : _GEN_989; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_991 = 7'h58 == index[6:0] ? dirty_1_88 : _GEN_990; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_992 = 7'h59 == index[6:0] ? dirty_1_89 : _GEN_991; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_993 = 7'h5a == index[6:0] ? dirty_1_90 : _GEN_992; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_994 = 7'h5b == index[6:0] ? dirty_1_91 : _GEN_993; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_995 = 7'h5c == index[6:0] ? dirty_1_92 : _GEN_994; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_996 = 7'h5d == index[6:0] ? dirty_1_93 : _GEN_995; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_997 = 7'h5e == index[6:0] ? dirty_1_94 : _GEN_996; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_998 = 7'h5f == index[6:0] ? dirty_1_95 : _GEN_997; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_999 = 7'h60 == index[6:0] ? dirty_1_96 : _GEN_998; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1000 = 7'h61 == index[6:0] ? dirty_1_97 : _GEN_999; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1001 = 7'h62 == index[6:0] ? dirty_1_98 : _GEN_1000; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1002 = 7'h63 == index[6:0] ? dirty_1_99 : _GEN_1001; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1003 = 7'h64 == index[6:0] ? dirty_1_100 : _GEN_1002; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1004 = 7'h65 == index[6:0] ? dirty_1_101 : _GEN_1003; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1005 = 7'h66 == index[6:0] ? dirty_1_102 : _GEN_1004; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1006 = 7'h67 == index[6:0] ? dirty_1_103 : _GEN_1005; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1007 = 7'h68 == index[6:0] ? dirty_1_104 : _GEN_1006; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1008 = 7'h69 == index[6:0] ? dirty_1_105 : _GEN_1007; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1009 = 7'h6a == index[6:0] ? dirty_1_106 : _GEN_1008; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1010 = 7'h6b == index[6:0] ? dirty_1_107 : _GEN_1009; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1011 = 7'h6c == index[6:0] ? dirty_1_108 : _GEN_1010; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1012 = 7'h6d == index[6:0] ? dirty_1_109 : _GEN_1011; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1013 = 7'h6e == index[6:0] ? dirty_1_110 : _GEN_1012; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1014 = 7'h6f == index[6:0] ? dirty_1_111 : _GEN_1013; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1015 = 7'h70 == index[6:0] ? dirty_1_112 : _GEN_1014; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1016 = 7'h71 == index[6:0] ? dirty_1_113 : _GEN_1015; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1017 = 7'h72 == index[6:0] ? dirty_1_114 : _GEN_1016; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1018 = 7'h73 == index[6:0] ? dirty_1_115 : _GEN_1017; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1019 = 7'h74 == index[6:0] ? dirty_1_116 : _GEN_1018; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1020 = 7'h75 == index[6:0] ? dirty_1_117 : _GEN_1019; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1021 = 7'h76 == index[6:0] ? dirty_1_118 : _GEN_1020; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1022 = 7'h77 == index[6:0] ? dirty_1_119 : _GEN_1021; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1023 = 7'h78 == index[6:0] ? dirty_1_120 : _GEN_1022; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1024 = 7'h79 == index[6:0] ? dirty_1_121 : _GEN_1023; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1025 = 7'h7a == index[6:0] ? dirty_1_122 : _GEN_1024; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1026 = 7'h7b == index[6:0] ? dirty_1_123 : _GEN_1025; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1027 = 7'h7c == index[6:0] ? dirty_1_124 : _GEN_1026; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1028 = 7'h7d == index[6:0] ? dirty_1_125 : _GEN_1027; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1029 = 7'h7e == index[6:0] ? dirty_1_126 : _GEN_1028; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_1030 = 7'h7f == index[6:0] ? dirty_1_127 : _GEN_1029; // @[d_cache.scala 99:{27,27}]
  wire [2:0] _GEN_1031 = way1_hit ? _GEN_902 : 3'h3; // @[d_cache.scala 103:23 97:33]
  wire [63:0] _GEN_18467 = {{32'd0}, io_from_lsu_wdata}; // @[d_cache.scala 109:53]
  wire [63:0] _ram_0_T = _GEN_18467 & wmask; // @[d_cache.scala 109:53]
  wire [126:0] _GEN_19511 = {{63'd0}, _ram_0_T}; // @[d_cache.scala 109:62]
  wire [126:0] _ram_0_T_1 = _GEN_19511 << shift_bit; // @[d_cache.scala 109:62]
  wire [126:0] _GEN_19512 = {{63'd0}, wmask}; // @[d_cache.scala 109:102]
  wire [126:0] _ram_0_T_3 = _GEN_19512 << shift_bit; // @[d_cache.scala 109:102]
  wire [126:0] _ram_0_T_4 = ~_ram_0_T_3; // @[d_cache.scala 109:94]
  wire [63:0] _GEN_1034 = 7'h1 == index[6:0] ? ram_0_1 : ram_0_0; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1035 = 7'h2 == index[6:0] ? ram_0_2 : _GEN_1034; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1036 = 7'h3 == index[6:0] ? ram_0_3 : _GEN_1035; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1037 = 7'h4 == index[6:0] ? ram_0_4 : _GEN_1036; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1038 = 7'h5 == index[6:0] ? ram_0_5 : _GEN_1037; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1039 = 7'h6 == index[6:0] ? ram_0_6 : _GEN_1038; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1040 = 7'h7 == index[6:0] ? ram_0_7 : _GEN_1039; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1041 = 7'h8 == index[6:0] ? ram_0_8 : _GEN_1040; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1042 = 7'h9 == index[6:0] ? ram_0_9 : _GEN_1041; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1043 = 7'ha == index[6:0] ? ram_0_10 : _GEN_1042; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1044 = 7'hb == index[6:0] ? ram_0_11 : _GEN_1043; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1045 = 7'hc == index[6:0] ? ram_0_12 : _GEN_1044; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1046 = 7'hd == index[6:0] ? ram_0_13 : _GEN_1045; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1047 = 7'he == index[6:0] ? ram_0_14 : _GEN_1046; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1048 = 7'hf == index[6:0] ? ram_0_15 : _GEN_1047; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1049 = 7'h10 == index[6:0] ? ram_0_16 : _GEN_1048; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1050 = 7'h11 == index[6:0] ? ram_0_17 : _GEN_1049; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1051 = 7'h12 == index[6:0] ? ram_0_18 : _GEN_1050; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1052 = 7'h13 == index[6:0] ? ram_0_19 : _GEN_1051; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1053 = 7'h14 == index[6:0] ? ram_0_20 : _GEN_1052; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1054 = 7'h15 == index[6:0] ? ram_0_21 : _GEN_1053; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1055 = 7'h16 == index[6:0] ? ram_0_22 : _GEN_1054; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1056 = 7'h17 == index[6:0] ? ram_0_23 : _GEN_1055; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1057 = 7'h18 == index[6:0] ? ram_0_24 : _GEN_1056; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1058 = 7'h19 == index[6:0] ? ram_0_25 : _GEN_1057; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1059 = 7'h1a == index[6:0] ? ram_0_26 : _GEN_1058; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1060 = 7'h1b == index[6:0] ? ram_0_27 : _GEN_1059; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1061 = 7'h1c == index[6:0] ? ram_0_28 : _GEN_1060; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1062 = 7'h1d == index[6:0] ? ram_0_29 : _GEN_1061; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1063 = 7'h1e == index[6:0] ? ram_0_30 : _GEN_1062; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1064 = 7'h1f == index[6:0] ? ram_0_31 : _GEN_1063; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1065 = 7'h20 == index[6:0] ? ram_0_32 : _GEN_1064; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1066 = 7'h21 == index[6:0] ? ram_0_33 : _GEN_1065; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1067 = 7'h22 == index[6:0] ? ram_0_34 : _GEN_1066; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1068 = 7'h23 == index[6:0] ? ram_0_35 : _GEN_1067; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1069 = 7'h24 == index[6:0] ? ram_0_36 : _GEN_1068; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1070 = 7'h25 == index[6:0] ? ram_0_37 : _GEN_1069; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1071 = 7'h26 == index[6:0] ? ram_0_38 : _GEN_1070; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1072 = 7'h27 == index[6:0] ? ram_0_39 : _GEN_1071; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1073 = 7'h28 == index[6:0] ? ram_0_40 : _GEN_1072; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1074 = 7'h29 == index[6:0] ? ram_0_41 : _GEN_1073; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1075 = 7'h2a == index[6:0] ? ram_0_42 : _GEN_1074; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1076 = 7'h2b == index[6:0] ? ram_0_43 : _GEN_1075; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1077 = 7'h2c == index[6:0] ? ram_0_44 : _GEN_1076; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1078 = 7'h2d == index[6:0] ? ram_0_45 : _GEN_1077; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1079 = 7'h2e == index[6:0] ? ram_0_46 : _GEN_1078; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1080 = 7'h2f == index[6:0] ? ram_0_47 : _GEN_1079; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1081 = 7'h30 == index[6:0] ? ram_0_48 : _GEN_1080; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1082 = 7'h31 == index[6:0] ? ram_0_49 : _GEN_1081; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1083 = 7'h32 == index[6:0] ? ram_0_50 : _GEN_1082; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1084 = 7'h33 == index[6:0] ? ram_0_51 : _GEN_1083; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1085 = 7'h34 == index[6:0] ? ram_0_52 : _GEN_1084; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1086 = 7'h35 == index[6:0] ? ram_0_53 : _GEN_1085; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1087 = 7'h36 == index[6:0] ? ram_0_54 : _GEN_1086; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1088 = 7'h37 == index[6:0] ? ram_0_55 : _GEN_1087; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1089 = 7'h38 == index[6:0] ? ram_0_56 : _GEN_1088; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1090 = 7'h39 == index[6:0] ? ram_0_57 : _GEN_1089; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1091 = 7'h3a == index[6:0] ? ram_0_58 : _GEN_1090; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1092 = 7'h3b == index[6:0] ? ram_0_59 : _GEN_1091; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1093 = 7'h3c == index[6:0] ? ram_0_60 : _GEN_1092; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1094 = 7'h3d == index[6:0] ? ram_0_61 : _GEN_1093; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1095 = 7'h3e == index[6:0] ? ram_0_62 : _GEN_1094; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1096 = 7'h3f == index[6:0] ? ram_0_63 : _GEN_1095; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1097 = 7'h40 == index[6:0] ? ram_0_64 : _GEN_1096; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1098 = 7'h41 == index[6:0] ? ram_0_65 : _GEN_1097; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1099 = 7'h42 == index[6:0] ? ram_0_66 : _GEN_1098; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1100 = 7'h43 == index[6:0] ? ram_0_67 : _GEN_1099; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1101 = 7'h44 == index[6:0] ? ram_0_68 : _GEN_1100; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1102 = 7'h45 == index[6:0] ? ram_0_69 : _GEN_1101; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1103 = 7'h46 == index[6:0] ? ram_0_70 : _GEN_1102; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1104 = 7'h47 == index[6:0] ? ram_0_71 : _GEN_1103; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1105 = 7'h48 == index[6:0] ? ram_0_72 : _GEN_1104; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1106 = 7'h49 == index[6:0] ? ram_0_73 : _GEN_1105; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1107 = 7'h4a == index[6:0] ? ram_0_74 : _GEN_1106; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1108 = 7'h4b == index[6:0] ? ram_0_75 : _GEN_1107; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1109 = 7'h4c == index[6:0] ? ram_0_76 : _GEN_1108; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1110 = 7'h4d == index[6:0] ? ram_0_77 : _GEN_1109; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1111 = 7'h4e == index[6:0] ? ram_0_78 : _GEN_1110; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1112 = 7'h4f == index[6:0] ? ram_0_79 : _GEN_1111; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1113 = 7'h50 == index[6:0] ? ram_0_80 : _GEN_1112; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1114 = 7'h51 == index[6:0] ? ram_0_81 : _GEN_1113; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1115 = 7'h52 == index[6:0] ? ram_0_82 : _GEN_1114; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1116 = 7'h53 == index[6:0] ? ram_0_83 : _GEN_1115; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1117 = 7'h54 == index[6:0] ? ram_0_84 : _GEN_1116; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1118 = 7'h55 == index[6:0] ? ram_0_85 : _GEN_1117; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1119 = 7'h56 == index[6:0] ? ram_0_86 : _GEN_1118; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1120 = 7'h57 == index[6:0] ? ram_0_87 : _GEN_1119; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1121 = 7'h58 == index[6:0] ? ram_0_88 : _GEN_1120; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1122 = 7'h59 == index[6:0] ? ram_0_89 : _GEN_1121; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1123 = 7'h5a == index[6:0] ? ram_0_90 : _GEN_1122; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1124 = 7'h5b == index[6:0] ? ram_0_91 : _GEN_1123; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1125 = 7'h5c == index[6:0] ? ram_0_92 : _GEN_1124; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1126 = 7'h5d == index[6:0] ? ram_0_93 : _GEN_1125; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1127 = 7'h5e == index[6:0] ? ram_0_94 : _GEN_1126; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1128 = 7'h5f == index[6:0] ? ram_0_95 : _GEN_1127; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1129 = 7'h60 == index[6:0] ? ram_0_96 : _GEN_1128; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1130 = 7'h61 == index[6:0] ? ram_0_97 : _GEN_1129; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1131 = 7'h62 == index[6:0] ? ram_0_98 : _GEN_1130; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1132 = 7'h63 == index[6:0] ? ram_0_99 : _GEN_1131; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1133 = 7'h64 == index[6:0] ? ram_0_100 : _GEN_1132; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1134 = 7'h65 == index[6:0] ? ram_0_101 : _GEN_1133; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1135 = 7'h66 == index[6:0] ? ram_0_102 : _GEN_1134; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1136 = 7'h67 == index[6:0] ? ram_0_103 : _GEN_1135; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1137 = 7'h68 == index[6:0] ? ram_0_104 : _GEN_1136; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1138 = 7'h69 == index[6:0] ? ram_0_105 : _GEN_1137; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1139 = 7'h6a == index[6:0] ? ram_0_106 : _GEN_1138; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1140 = 7'h6b == index[6:0] ? ram_0_107 : _GEN_1139; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1141 = 7'h6c == index[6:0] ? ram_0_108 : _GEN_1140; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1142 = 7'h6d == index[6:0] ? ram_0_109 : _GEN_1141; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1143 = 7'h6e == index[6:0] ? ram_0_110 : _GEN_1142; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1144 = 7'h6f == index[6:0] ? ram_0_111 : _GEN_1143; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1145 = 7'h70 == index[6:0] ? ram_0_112 : _GEN_1144; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1146 = 7'h71 == index[6:0] ? ram_0_113 : _GEN_1145; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1147 = 7'h72 == index[6:0] ? ram_0_114 : _GEN_1146; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1148 = 7'h73 == index[6:0] ? ram_0_115 : _GEN_1147; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1149 = 7'h74 == index[6:0] ? ram_0_116 : _GEN_1148; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1150 = 7'h75 == index[6:0] ? ram_0_117 : _GEN_1149; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1151 = 7'h76 == index[6:0] ? ram_0_118 : _GEN_1150; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1152 = 7'h77 == index[6:0] ? ram_0_119 : _GEN_1151; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1153 = 7'h78 == index[6:0] ? ram_0_120 : _GEN_1152; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1154 = 7'h79 == index[6:0] ? ram_0_121 : _GEN_1153; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1155 = 7'h7a == index[6:0] ? ram_0_122 : _GEN_1154; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1156 = 7'h7b == index[6:0] ? ram_0_123 : _GEN_1155; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1157 = 7'h7c == index[6:0] ? ram_0_124 : _GEN_1156; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1158 = 7'h7d == index[6:0] ? ram_0_125 : _GEN_1157; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1159 = 7'h7e == index[6:0] ? ram_0_126 : _GEN_1158; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_1160 = 7'h7f == index[6:0] ? ram_0_127 : _GEN_1159; // @[d_cache.scala 109:{92,92}]
  wire [126:0] _GEN_18468 = {{63'd0}, _GEN_1160}; // @[d_cache.scala 109:92]
  wire [126:0] _ram_0_T_5 = _GEN_18468 & _ram_0_T_4; // @[d_cache.scala 109:92]
  wire [126:0] _ram_0_T_6 = _ram_0_T_1 | _ram_0_T_5; // @[d_cache.scala 109:76]
  wire [63:0] _GEN_1161 = 7'h0 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_0; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1162 = 7'h1 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_1; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1163 = 7'h2 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_2; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1164 = 7'h3 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_3; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1165 = 7'h4 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_4; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1166 = 7'h5 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_5; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1167 = 7'h6 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_6; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1168 = 7'h7 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_7; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1169 = 7'h8 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_8; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1170 = 7'h9 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_9; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1171 = 7'ha == index[6:0] ? _ram_0_T_6[63:0] : ram_0_10; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1172 = 7'hb == index[6:0] ? _ram_0_T_6[63:0] : ram_0_11; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1173 = 7'hc == index[6:0] ? _ram_0_T_6[63:0] : ram_0_12; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1174 = 7'hd == index[6:0] ? _ram_0_T_6[63:0] : ram_0_13; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1175 = 7'he == index[6:0] ? _ram_0_T_6[63:0] : ram_0_14; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1176 = 7'hf == index[6:0] ? _ram_0_T_6[63:0] : ram_0_15; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1177 = 7'h10 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_16; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1178 = 7'h11 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_17; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1179 = 7'h12 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_18; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1180 = 7'h13 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_19; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1181 = 7'h14 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_20; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1182 = 7'h15 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_21; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1183 = 7'h16 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_22; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1184 = 7'h17 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_23; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1185 = 7'h18 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_24; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1186 = 7'h19 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_25; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1187 = 7'h1a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_26; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1188 = 7'h1b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_27; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1189 = 7'h1c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_28; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1190 = 7'h1d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_29; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1191 = 7'h1e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_30; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1192 = 7'h1f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_31; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1193 = 7'h20 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_32; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1194 = 7'h21 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_33; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1195 = 7'h22 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_34; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1196 = 7'h23 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_35; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1197 = 7'h24 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_36; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1198 = 7'h25 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_37; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1199 = 7'h26 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_38; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1200 = 7'h27 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_39; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1201 = 7'h28 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_40; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1202 = 7'h29 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_41; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1203 = 7'h2a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_42; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1204 = 7'h2b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_43; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1205 = 7'h2c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_44; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1206 = 7'h2d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_45; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1207 = 7'h2e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_46; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1208 = 7'h2f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_47; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1209 = 7'h30 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_48; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1210 = 7'h31 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_49; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1211 = 7'h32 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_50; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1212 = 7'h33 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_51; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1213 = 7'h34 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_52; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1214 = 7'h35 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_53; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1215 = 7'h36 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_54; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1216 = 7'h37 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_55; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1217 = 7'h38 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_56; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1218 = 7'h39 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_57; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1219 = 7'h3a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_58; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1220 = 7'h3b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_59; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1221 = 7'h3c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_60; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1222 = 7'h3d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_61; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1223 = 7'h3e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_62; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1224 = 7'h3f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_63; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1225 = 7'h40 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_64; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1226 = 7'h41 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_65; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1227 = 7'h42 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_66; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1228 = 7'h43 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_67; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1229 = 7'h44 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_68; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1230 = 7'h45 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_69; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1231 = 7'h46 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_70; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1232 = 7'h47 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_71; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1233 = 7'h48 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_72; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1234 = 7'h49 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_73; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1235 = 7'h4a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_74; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1236 = 7'h4b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_75; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1237 = 7'h4c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_76; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1238 = 7'h4d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_77; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1239 = 7'h4e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_78; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1240 = 7'h4f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_79; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1241 = 7'h50 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_80; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1242 = 7'h51 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_81; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1243 = 7'h52 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_82; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1244 = 7'h53 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_83; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1245 = 7'h54 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_84; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1246 = 7'h55 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_85; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1247 = 7'h56 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_86; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1248 = 7'h57 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_87; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1249 = 7'h58 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_88; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1250 = 7'h59 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_89; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1251 = 7'h5a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_90; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1252 = 7'h5b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_91; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1253 = 7'h5c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_92; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1254 = 7'h5d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_93; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1255 = 7'h5e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_94; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1256 = 7'h5f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_95; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1257 = 7'h60 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_96; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1258 = 7'h61 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_97; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1259 = 7'h62 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_98; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1260 = 7'h63 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_99; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1261 = 7'h64 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_100; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1262 = 7'h65 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_101; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1263 = 7'h66 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_102; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1264 = 7'h67 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_103; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1265 = 7'h68 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_104; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1266 = 7'h69 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_105; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1267 = 7'h6a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_106; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1268 = 7'h6b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_107; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1269 = 7'h6c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_108; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1270 = 7'h6d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_109; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1271 = 7'h6e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_110; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1272 = 7'h6f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_111; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1273 = 7'h70 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_112; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1274 = 7'h71 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_113; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1275 = 7'h72 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_114; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1276 = 7'h73 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_115; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1277 = 7'h74 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_116; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1278 = 7'h75 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_117; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1279 = 7'h76 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_118; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1280 = 7'h77 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_119; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1281 = 7'h78 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_120; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1282 = 7'h79 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_121; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1283 = 7'h7a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_122; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1284 = 7'h7b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_123; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1285 = 7'h7c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_124; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1286 = 7'h7d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_125; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1287 = 7'h7e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_126; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1288 = 7'h7f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_127; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_1289 = 7'h0 == index[6:0] ? _ram_0_T : recent_wdata0_0; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1290 = 7'h1 == index[6:0] ? _ram_0_T : recent_wdata0_1; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1291 = 7'h2 == index[6:0] ? _ram_0_T : recent_wdata0_2; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1292 = 7'h3 == index[6:0] ? _ram_0_T : recent_wdata0_3; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1293 = 7'h4 == index[6:0] ? _ram_0_T : recent_wdata0_4; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1294 = 7'h5 == index[6:0] ? _ram_0_T : recent_wdata0_5; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1295 = 7'h6 == index[6:0] ? _ram_0_T : recent_wdata0_6; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1296 = 7'h7 == index[6:0] ? _ram_0_T : recent_wdata0_7; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1297 = 7'h8 == index[6:0] ? _ram_0_T : recent_wdata0_8; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1298 = 7'h9 == index[6:0] ? _ram_0_T : recent_wdata0_9; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1299 = 7'ha == index[6:0] ? _ram_0_T : recent_wdata0_10; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1300 = 7'hb == index[6:0] ? _ram_0_T : recent_wdata0_11; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1301 = 7'hc == index[6:0] ? _ram_0_T : recent_wdata0_12; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1302 = 7'hd == index[6:0] ? _ram_0_T : recent_wdata0_13; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1303 = 7'he == index[6:0] ? _ram_0_T : recent_wdata0_14; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1304 = 7'hf == index[6:0] ? _ram_0_T : recent_wdata0_15; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1305 = 7'h10 == index[6:0] ? _ram_0_T : recent_wdata0_16; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1306 = 7'h11 == index[6:0] ? _ram_0_T : recent_wdata0_17; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1307 = 7'h12 == index[6:0] ? _ram_0_T : recent_wdata0_18; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1308 = 7'h13 == index[6:0] ? _ram_0_T : recent_wdata0_19; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1309 = 7'h14 == index[6:0] ? _ram_0_T : recent_wdata0_20; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1310 = 7'h15 == index[6:0] ? _ram_0_T : recent_wdata0_21; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1311 = 7'h16 == index[6:0] ? _ram_0_T : recent_wdata0_22; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1312 = 7'h17 == index[6:0] ? _ram_0_T : recent_wdata0_23; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1313 = 7'h18 == index[6:0] ? _ram_0_T : recent_wdata0_24; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1314 = 7'h19 == index[6:0] ? _ram_0_T : recent_wdata0_25; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1315 = 7'h1a == index[6:0] ? _ram_0_T : recent_wdata0_26; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1316 = 7'h1b == index[6:0] ? _ram_0_T : recent_wdata0_27; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1317 = 7'h1c == index[6:0] ? _ram_0_T : recent_wdata0_28; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1318 = 7'h1d == index[6:0] ? _ram_0_T : recent_wdata0_29; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1319 = 7'h1e == index[6:0] ? _ram_0_T : recent_wdata0_30; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1320 = 7'h1f == index[6:0] ? _ram_0_T : recent_wdata0_31; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1321 = 7'h20 == index[6:0] ? _ram_0_T : recent_wdata0_32; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1322 = 7'h21 == index[6:0] ? _ram_0_T : recent_wdata0_33; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1323 = 7'h22 == index[6:0] ? _ram_0_T : recent_wdata0_34; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1324 = 7'h23 == index[6:0] ? _ram_0_T : recent_wdata0_35; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1325 = 7'h24 == index[6:0] ? _ram_0_T : recent_wdata0_36; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1326 = 7'h25 == index[6:0] ? _ram_0_T : recent_wdata0_37; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1327 = 7'h26 == index[6:0] ? _ram_0_T : recent_wdata0_38; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1328 = 7'h27 == index[6:0] ? _ram_0_T : recent_wdata0_39; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1329 = 7'h28 == index[6:0] ? _ram_0_T : recent_wdata0_40; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1330 = 7'h29 == index[6:0] ? _ram_0_T : recent_wdata0_41; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1331 = 7'h2a == index[6:0] ? _ram_0_T : recent_wdata0_42; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1332 = 7'h2b == index[6:0] ? _ram_0_T : recent_wdata0_43; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1333 = 7'h2c == index[6:0] ? _ram_0_T : recent_wdata0_44; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1334 = 7'h2d == index[6:0] ? _ram_0_T : recent_wdata0_45; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1335 = 7'h2e == index[6:0] ? _ram_0_T : recent_wdata0_46; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1336 = 7'h2f == index[6:0] ? _ram_0_T : recent_wdata0_47; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1337 = 7'h30 == index[6:0] ? _ram_0_T : recent_wdata0_48; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1338 = 7'h31 == index[6:0] ? _ram_0_T : recent_wdata0_49; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1339 = 7'h32 == index[6:0] ? _ram_0_T : recent_wdata0_50; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1340 = 7'h33 == index[6:0] ? _ram_0_T : recent_wdata0_51; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1341 = 7'h34 == index[6:0] ? _ram_0_T : recent_wdata0_52; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1342 = 7'h35 == index[6:0] ? _ram_0_T : recent_wdata0_53; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1343 = 7'h36 == index[6:0] ? _ram_0_T : recent_wdata0_54; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1344 = 7'h37 == index[6:0] ? _ram_0_T : recent_wdata0_55; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1345 = 7'h38 == index[6:0] ? _ram_0_T : recent_wdata0_56; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1346 = 7'h39 == index[6:0] ? _ram_0_T : recent_wdata0_57; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1347 = 7'h3a == index[6:0] ? _ram_0_T : recent_wdata0_58; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1348 = 7'h3b == index[6:0] ? _ram_0_T : recent_wdata0_59; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1349 = 7'h3c == index[6:0] ? _ram_0_T : recent_wdata0_60; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1350 = 7'h3d == index[6:0] ? _ram_0_T : recent_wdata0_61; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1351 = 7'h3e == index[6:0] ? _ram_0_T : recent_wdata0_62; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1352 = 7'h3f == index[6:0] ? _ram_0_T : recent_wdata0_63; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1353 = 7'h40 == index[6:0] ? _ram_0_T : recent_wdata0_64; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1354 = 7'h41 == index[6:0] ? _ram_0_T : recent_wdata0_65; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1355 = 7'h42 == index[6:0] ? _ram_0_T : recent_wdata0_66; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1356 = 7'h43 == index[6:0] ? _ram_0_T : recent_wdata0_67; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1357 = 7'h44 == index[6:0] ? _ram_0_T : recent_wdata0_68; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1358 = 7'h45 == index[6:0] ? _ram_0_T : recent_wdata0_69; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1359 = 7'h46 == index[6:0] ? _ram_0_T : recent_wdata0_70; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1360 = 7'h47 == index[6:0] ? _ram_0_T : recent_wdata0_71; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1361 = 7'h48 == index[6:0] ? _ram_0_T : recent_wdata0_72; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1362 = 7'h49 == index[6:0] ? _ram_0_T : recent_wdata0_73; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1363 = 7'h4a == index[6:0] ? _ram_0_T : recent_wdata0_74; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1364 = 7'h4b == index[6:0] ? _ram_0_T : recent_wdata0_75; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1365 = 7'h4c == index[6:0] ? _ram_0_T : recent_wdata0_76; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1366 = 7'h4d == index[6:0] ? _ram_0_T : recent_wdata0_77; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1367 = 7'h4e == index[6:0] ? _ram_0_T : recent_wdata0_78; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1368 = 7'h4f == index[6:0] ? _ram_0_T : recent_wdata0_79; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1369 = 7'h50 == index[6:0] ? _ram_0_T : recent_wdata0_80; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1370 = 7'h51 == index[6:0] ? _ram_0_T : recent_wdata0_81; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1371 = 7'h52 == index[6:0] ? _ram_0_T : recent_wdata0_82; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1372 = 7'h53 == index[6:0] ? _ram_0_T : recent_wdata0_83; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1373 = 7'h54 == index[6:0] ? _ram_0_T : recent_wdata0_84; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1374 = 7'h55 == index[6:0] ? _ram_0_T : recent_wdata0_85; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1375 = 7'h56 == index[6:0] ? _ram_0_T : recent_wdata0_86; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1376 = 7'h57 == index[6:0] ? _ram_0_T : recent_wdata0_87; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1377 = 7'h58 == index[6:0] ? _ram_0_T : recent_wdata0_88; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1378 = 7'h59 == index[6:0] ? _ram_0_T : recent_wdata0_89; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1379 = 7'h5a == index[6:0] ? _ram_0_T : recent_wdata0_90; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1380 = 7'h5b == index[6:0] ? _ram_0_T : recent_wdata0_91; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1381 = 7'h5c == index[6:0] ? _ram_0_T : recent_wdata0_92; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1382 = 7'h5d == index[6:0] ? _ram_0_T : recent_wdata0_93; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1383 = 7'h5e == index[6:0] ? _ram_0_T : recent_wdata0_94; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1384 = 7'h5f == index[6:0] ? _ram_0_T : recent_wdata0_95; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1385 = 7'h60 == index[6:0] ? _ram_0_T : recent_wdata0_96; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1386 = 7'h61 == index[6:0] ? _ram_0_T : recent_wdata0_97; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1387 = 7'h62 == index[6:0] ? _ram_0_T : recent_wdata0_98; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1388 = 7'h63 == index[6:0] ? _ram_0_T : recent_wdata0_99; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1389 = 7'h64 == index[6:0] ? _ram_0_T : recent_wdata0_100; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1390 = 7'h65 == index[6:0] ? _ram_0_T : recent_wdata0_101; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1391 = 7'h66 == index[6:0] ? _ram_0_T : recent_wdata0_102; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1392 = 7'h67 == index[6:0] ? _ram_0_T : recent_wdata0_103; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1393 = 7'h68 == index[6:0] ? _ram_0_T : recent_wdata0_104; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1394 = 7'h69 == index[6:0] ? _ram_0_T : recent_wdata0_105; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1395 = 7'h6a == index[6:0] ? _ram_0_T : recent_wdata0_106; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1396 = 7'h6b == index[6:0] ? _ram_0_T : recent_wdata0_107; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1397 = 7'h6c == index[6:0] ? _ram_0_T : recent_wdata0_108; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1398 = 7'h6d == index[6:0] ? _ram_0_T : recent_wdata0_109; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1399 = 7'h6e == index[6:0] ? _ram_0_T : recent_wdata0_110; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1400 = 7'h6f == index[6:0] ? _ram_0_T : recent_wdata0_111; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1401 = 7'h70 == index[6:0] ? _ram_0_T : recent_wdata0_112; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1402 = 7'h71 == index[6:0] ? _ram_0_T : recent_wdata0_113; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1403 = 7'h72 == index[6:0] ? _ram_0_T : recent_wdata0_114; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1404 = 7'h73 == index[6:0] ? _ram_0_T : recent_wdata0_115; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1405 = 7'h74 == index[6:0] ? _ram_0_T : recent_wdata0_116; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1406 = 7'h75 == index[6:0] ? _ram_0_T : recent_wdata0_117; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1407 = 7'h76 == index[6:0] ? _ram_0_T : recent_wdata0_118; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1408 = 7'h77 == index[6:0] ? _ram_0_T : recent_wdata0_119; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1409 = 7'h78 == index[6:0] ? _ram_0_T : recent_wdata0_120; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1410 = 7'h79 == index[6:0] ? _ram_0_T : recent_wdata0_121; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1411 = 7'h7a == index[6:0] ? _ram_0_T : recent_wdata0_122; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1412 = 7'h7b == index[6:0] ? _ram_0_T : recent_wdata0_123; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1413 = 7'h7c == index[6:0] ? _ram_0_T : recent_wdata0_124; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1414 = 7'h7d == index[6:0] ? _ram_0_T : recent_wdata0_125; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1415 = 7'h7e == index[6:0] ? _ram_0_T : recent_wdata0_126; // @[d_cache.scala 110:{38,38} 20:32]
  wire [63:0] _GEN_1416 = 7'h7f == index[6:0] ? _ram_0_T : recent_wdata0_127; // @[d_cache.scala 110:{38,38} 20:32]
  wire  _GEN_18470 = 7'h0 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1417 = 7'h0 == index[6:0] | dirty_0_0; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18471 = 7'h1 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1418 = 7'h1 == index[6:0] | dirty_0_1; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18472 = 7'h2 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1419 = 7'h2 == index[6:0] | dirty_0_2; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18473 = 7'h3 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1420 = 7'h3 == index[6:0] | dirty_0_3; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18474 = 7'h4 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1421 = 7'h4 == index[6:0] | dirty_0_4; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18475 = 7'h5 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1422 = 7'h5 == index[6:0] | dirty_0_5; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18476 = 7'h6 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1423 = 7'h6 == index[6:0] | dirty_0_6; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18477 = 7'h7 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1424 = 7'h7 == index[6:0] | dirty_0_7; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18478 = 7'h8 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1425 = 7'h8 == index[6:0] | dirty_0_8; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18479 = 7'h9 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1426 = 7'h9 == index[6:0] | dirty_0_9; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18480 = 7'ha == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1427 = 7'ha == index[6:0] | dirty_0_10; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18481 = 7'hb == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1428 = 7'hb == index[6:0] | dirty_0_11; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18482 = 7'hc == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1429 = 7'hc == index[6:0] | dirty_0_12; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18483 = 7'hd == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1430 = 7'hd == index[6:0] | dirty_0_13; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18484 = 7'he == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1431 = 7'he == index[6:0] | dirty_0_14; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18485 = 7'hf == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1432 = 7'hf == index[6:0] | dirty_0_15; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18486 = 7'h10 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1433 = 7'h10 == index[6:0] | dirty_0_16; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18487 = 7'h11 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1434 = 7'h11 == index[6:0] | dirty_0_17; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18488 = 7'h12 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1435 = 7'h12 == index[6:0] | dirty_0_18; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18489 = 7'h13 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1436 = 7'h13 == index[6:0] | dirty_0_19; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18490 = 7'h14 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1437 = 7'h14 == index[6:0] | dirty_0_20; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18491 = 7'h15 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1438 = 7'h15 == index[6:0] | dirty_0_21; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18492 = 7'h16 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1439 = 7'h16 == index[6:0] | dirty_0_22; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18493 = 7'h17 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1440 = 7'h17 == index[6:0] | dirty_0_23; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18494 = 7'h18 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1441 = 7'h18 == index[6:0] | dirty_0_24; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18495 = 7'h19 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1442 = 7'h19 == index[6:0] | dirty_0_25; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18496 = 7'h1a == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1443 = 7'h1a == index[6:0] | dirty_0_26; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18497 = 7'h1b == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1444 = 7'h1b == index[6:0] | dirty_0_27; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18498 = 7'h1c == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1445 = 7'h1c == index[6:0] | dirty_0_28; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18499 = 7'h1d == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1446 = 7'h1d == index[6:0] | dirty_0_29; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18500 = 7'h1e == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1447 = 7'h1e == index[6:0] | dirty_0_30; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18501 = 7'h1f == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1448 = 7'h1f == index[6:0] | dirty_0_31; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18502 = 7'h20 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1449 = 7'h20 == index[6:0] | dirty_0_32; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18503 = 7'h21 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1450 = 7'h21 == index[6:0] | dirty_0_33; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18504 = 7'h22 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1451 = 7'h22 == index[6:0] | dirty_0_34; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18505 = 7'h23 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1452 = 7'h23 == index[6:0] | dirty_0_35; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18506 = 7'h24 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1453 = 7'h24 == index[6:0] | dirty_0_36; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18507 = 7'h25 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1454 = 7'h25 == index[6:0] | dirty_0_37; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18508 = 7'h26 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1455 = 7'h26 == index[6:0] | dirty_0_38; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18509 = 7'h27 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1456 = 7'h27 == index[6:0] | dirty_0_39; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18510 = 7'h28 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1457 = 7'h28 == index[6:0] | dirty_0_40; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18511 = 7'h29 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1458 = 7'h29 == index[6:0] | dirty_0_41; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18512 = 7'h2a == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1459 = 7'h2a == index[6:0] | dirty_0_42; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18513 = 7'h2b == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1460 = 7'h2b == index[6:0] | dirty_0_43; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18514 = 7'h2c == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1461 = 7'h2c == index[6:0] | dirty_0_44; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18515 = 7'h2d == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1462 = 7'h2d == index[6:0] | dirty_0_45; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18516 = 7'h2e == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1463 = 7'h2e == index[6:0] | dirty_0_46; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18517 = 7'h2f == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1464 = 7'h2f == index[6:0] | dirty_0_47; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18518 = 7'h30 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1465 = 7'h30 == index[6:0] | dirty_0_48; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18519 = 7'h31 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1466 = 7'h31 == index[6:0] | dirty_0_49; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18520 = 7'h32 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1467 = 7'h32 == index[6:0] | dirty_0_50; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18521 = 7'h33 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1468 = 7'h33 == index[6:0] | dirty_0_51; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18522 = 7'h34 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1469 = 7'h34 == index[6:0] | dirty_0_52; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18523 = 7'h35 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1470 = 7'h35 == index[6:0] | dirty_0_53; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18524 = 7'h36 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1471 = 7'h36 == index[6:0] | dirty_0_54; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18525 = 7'h37 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1472 = 7'h37 == index[6:0] | dirty_0_55; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18526 = 7'h38 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1473 = 7'h38 == index[6:0] | dirty_0_56; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18527 = 7'h39 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1474 = 7'h39 == index[6:0] | dirty_0_57; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18528 = 7'h3a == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1475 = 7'h3a == index[6:0] | dirty_0_58; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18529 = 7'h3b == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1476 = 7'h3b == index[6:0] | dirty_0_59; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18530 = 7'h3c == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1477 = 7'h3c == index[6:0] | dirty_0_60; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18531 = 7'h3d == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1478 = 7'h3d == index[6:0] | dirty_0_61; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18532 = 7'h3e == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1479 = 7'h3e == index[6:0] | dirty_0_62; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18533 = 7'h3f == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1480 = 7'h3f == index[6:0] | dirty_0_63; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18534 = 7'h40 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1481 = 7'h40 == index[6:0] | dirty_0_64; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18535 = 7'h41 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1482 = 7'h41 == index[6:0] | dirty_0_65; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18536 = 7'h42 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1483 = 7'h42 == index[6:0] | dirty_0_66; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18537 = 7'h43 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1484 = 7'h43 == index[6:0] | dirty_0_67; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18538 = 7'h44 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1485 = 7'h44 == index[6:0] | dirty_0_68; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18539 = 7'h45 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1486 = 7'h45 == index[6:0] | dirty_0_69; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18540 = 7'h46 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1487 = 7'h46 == index[6:0] | dirty_0_70; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18541 = 7'h47 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1488 = 7'h47 == index[6:0] | dirty_0_71; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18542 = 7'h48 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1489 = 7'h48 == index[6:0] | dirty_0_72; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18543 = 7'h49 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1490 = 7'h49 == index[6:0] | dirty_0_73; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18544 = 7'h4a == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1491 = 7'h4a == index[6:0] | dirty_0_74; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18545 = 7'h4b == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1492 = 7'h4b == index[6:0] | dirty_0_75; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18546 = 7'h4c == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1493 = 7'h4c == index[6:0] | dirty_0_76; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18547 = 7'h4d == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1494 = 7'h4d == index[6:0] | dirty_0_77; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18548 = 7'h4e == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1495 = 7'h4e == index[6:0] | dirty_0_78; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18549 = 7'h4f == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1496 = 7'h4f == index[6:0] | dirty_0_79; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18550 = 7'h50 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1497 = 7'h50 == index[6:0] | dirty_0_80; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18551 = 7'h51 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1498 = 7'h51 == index[6:0] | dirty_0_81; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18552 = 7'h52 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1499 = 7'h52 == index[6:0] | dirty_0_82; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18553 = 7'h53 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1500 = 7'h53 == index[6:0] | dirty_0_83; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18554 = 7'h54 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1501 = 7'h54 == index[6:0] | dirty_0_84; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18555 = 7'h55 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1502 = 7'h55 == index[6:0] | dirty_0_85; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18556 = 7'h56 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1503 = 7'h56 == index[6:0] | dirty_0_86; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18557 = 7'h57 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1504 = 7'h57 == index[6:0] | dirty_0_87; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18558 = 7'h58 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1505 = 7'h58 == index[6:0] | dirty_0_88; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18559 = 7'h59 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1506 = 7'h59 == index[6:0] | dirty_0_89; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18560 = 7'h5a == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1507 = 7'h5a == index[6:0] | dirty_0_90; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18561 = 7'h5b == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1508 = 7'h5b == index[6:0] | dirty_0_91; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18562 = 7'h5c == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1509 = 7'h5c == index[6:0] | dirty_0_92; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18563 = 7'h5d == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1510 = 7'h5d == index[6:0] | dirty_0_93; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18564 = 7'h5e == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1511 = 7'h5e == index[6:0] | dirty_0_94; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18565 = 7'h5f == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1512 = 7'h5f == index[6:0] | dirty_0_95; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18566 = 7'h60 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1513 = 7'h60 == index[6:0] | dirty_0_96; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18567 = 7'h61 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1514 = 7'h61 == index[6:0] | dirty_0_97; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18568 = 7'h62 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1515 = 7'h62 == index[6:0] | dirty_0_98; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18569 = 7'h63 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1516 = 7'h63 == index[6:0] | dirty_0_99; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18570 = 7'h64 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1517 = 7'h64 == index[6:0] | dirty_0_100; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18571 = 7'h65 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1518 = 7'h65 == index[6:0] | dirty_0_101; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18572 = 7'h66 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1519 = 7'h66 == index[6:0] | dirty_0_102; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18573 = 7'h67 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1520 = 7'h67 == index[6:0] | dirty_0_103; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18574 = 7'h68 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1521 = 7'h68 == index[6:0] | dirty_0_104; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18575 = 7'h69 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1522 = 7'h69 == index[6:0] | dirty_0_105; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18576 = 7'h6a == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1523 = 7'h6a == index[6:0] | dirty_0_106; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18577 = 7'h6b == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1524 = 7'h6b == index[6:0] | dirty_0_107; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18578 = 7'h6c == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1525 = 7'h6c == index[6:0] | dirty_0_108; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18579 = 7'h6d == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1526 = 7'h6d == index[6:0] | dirty_0_109; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18580 = 7'h6e == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1527 = 7'h6e == index[6:0] | dirty_0_110; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18581 = 7'h6f == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1528 = 7'h6f == index[6:0] | dirty_0_111; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18582 = 7'h70 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1529 = 7'h70 == index[6:0] | dirty_0_112; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18583 = 7'h71 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1530 = 7'h71 == index[6:0] | dirty_0_113; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18584 = 7'h72 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1531 = 7'h72 == index[6:0] | dirty_0_114; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18585 = 7'h73 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1532 = 7'h73 == index[6:0] | dirty_0_115; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18586 = 7'h74 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1533 = 7'h74 == index[6:0] | dirty_0_116; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18587 = 7'h75 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1534 = 7'h75 == index[6:0] | dirty_0_117; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18588 = 7'h76 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1535 = 7'h76 == index[6:0] | dirty_0_118; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18589 = 7'h77 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1536 = 7'h77 == index[6:0] | dirty_0_119; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18590 = 7'h78 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1537 = 7'h78 == index[6:0] | dirty_0_120; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18591 = 7'h79 == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1538 = 7'h79 == index[6:0] | dirty_0_121; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18592 = 7'h7a == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1539 = 7'h7a == index[6:0] | dirty_0_122; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18593 = 7'h7b == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1540 = 7'h7b == index[6:0] | dirty_0_123; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18594 = 7'h7c == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1541 = 7'h7c == index[6:0] | dirty_0_124; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18595 = 7'h7d == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1542 = 7'h7d == index[6:0] | dirty_0_125; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18596 = 7'h7e == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1543 = 7'h7e == index[6:0] | dirty_0_126; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_18597 = 7'h7f == index[6:0]; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_1544 = 7'h7f == index[6:0] | dirty_0_127; // @[d_cache.scala 113:{32,32} 26:26]
  wire [63:0] _GEN_1546 = 7'h1 == index[6:0] ? ram_1_1 : ram_1_0; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1547 = 7'h2 == index[6:0] ? ram_1_2 : _GEN_1546; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1548 = 7'h3 == index[6:0] ? ram_1_3 : _GEN_1547; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1549 = 7'h4 == index[6:0] ? ram_1_4 : _GEN_1548; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1550 = 7'h5 == index[6:0] ? ram_1_5 : _GEN_1549; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1551 = 7'h6 == index[6:0] ? ram_1_6 : _GEN_1550; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1552 = 7'h7 == index[6:0] ? ram_1_7 : _GEN_1551; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1553 = 7'h8 == index[6:0] ? ram_1_8 : _GEN_1552; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1554 = 7'h9 == index[6:0] ? ram_1_9 : _GEN_1553; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1555 = 7'ha == index[6:0] ? ram_1_10 : _GEN_1554; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1556 = 7'hb == index[6:0] ? ram_1_11 : _GEN_1555; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1557 = 7'hc == index[6:0] ? ram_1_12 : _GEN_1556; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1558 = 7'hd == index[6:0] ? ram_1_13 : _GEN_1557; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1559 = 7'he == index[6:0] ? ram_1_14 : _GEN_1558; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1560 = 7'hf == index[6:0] ? ram_1_15 : _GEN_1559; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1561 = 7'h10 == index[6:0] ? ram_1_16 : _GEN_1560; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1562 = 7'h11 == index[6:0] ? ram_1_17 : _GEN_1561; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1563 = 7'h12 == index[6:0] ? ram_1_18 : _GEN_1562; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1564 = 7'h13 == index[6:0] ? ram_1_19 : _GEN_1563; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1565 = 7'h14 == index[6:0] ? ram_1_20 : _GEN_1564; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1566 = 7'h15 == index[6:0] ? ram_1_21 : _GEN_1565; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1567 = 7'h16 == index[6:0] ? ram_1_22 : _GEN_1566; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1568 = 7'h17 == index[6:0] ? ram_1_23 : _GEN_1567; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1569 = 7'h18 == index[6:0] ? ram_1_24 : _GEN_1568; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1570 = 7'h19 == index[6:0] ? ram_1_25 : _GEN_1569; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1571 = 7'h1a == index[6:0] ? ram_1_26 : _GEN_1570; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1572 = 7'h1b == index[6:0] ? ram_1_27 : _GEN_1571; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1573 = 7'h1c == index[6:0] ? ram_1_28 : _GEN_1572; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1574 = 7'h1d == index[6:0] ? ram_1_29 : _GEN_1573; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1575 = 7'h1e == index[6:0] ? ram_1_30 : _GEN_1574; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1576 = 7'h1f == index[6:0] ? ram_1_31 : _GEN_1575; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1577 = 7'h20 == index[6:0] ? ram_1_32 : _GEN_1576; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1578 = 7'h21 == index[6:0] ? ram_1_33 : _GEN_1577; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1579 = 7'h22 == index[6:0] ? ram_1_34 : _GEN_1578; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1580 = 7'h23 == index[6:0] ? ram_1_35 : _GEN_1579; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1581 = 7'h24 == index[6:0] ? ram_1_36 : _GEN_1580; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1582 = 7'h25 == index[6:0] ? ram_1_37 : _GEN_1581; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1583 = 7'h26 == index[6:0] ? ram_1_38 : _GEN_1582; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1584 = 7'h27 == index[6:0] ? ram_1_39 : _GEN_1583; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1585 = 7'h28 == index[6:0] ? ram_1_40 : _GEN_1584; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1586 = 7'h29 == index[6:0] ? ram_1_41 : _GEN_1585; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1587 = 7'h2a == index[6:0] ? ram_1_42 : _GEN_1586; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1588 = 7'h2b == index[6:0] ? ram_1_43 : _GEN_1587; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1589 = 7'h2c == index[6:0] ? ram_1_44 : _GEN_1588; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1590 = 7'h2d == index[6:0] ? ram_1_45 : _GEN_1589; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1591 = 7'h2e == index[6:0] ? ram_1_46 : _GEN_1590; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1592 = 7'h2f == index[6:0] ? ram_1_47 : _GEN_1591; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1593 = 7'h30 == index[6:0] ? ram_1_48 : _GEN_1592; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1594 = 7'h31 == index[6:0] ? ram_1_49 : _GEN_1593; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1595 = 7'h32 == index[6:0] ? ram_1_50 : _GEN_1594; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1596 = 7'h33 == index[6:0] ? ram_1_51 : _GEN_1595; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1597 = 7'h34 == index[6:0] ? ram_1_52 : _GEN_1596; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1598 = 7'h35 == index[6:0] ? ram_1_53 : _GEN_1597; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1599 = 7'h36 == index[6:0] ? ram_1_54 : _GEN_1598; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1600 = 7'h37 == index[6:0] ? ram_1_55 : _GEN_1599; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1601 = 7'h38 == index[6:0] ? ram_1_56 : _GEN_1600; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1602 = 7'h39 == index[6:0] ? ram_1_57 : _GEN_1601; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1603 = 7'h3a == index[6:0] ? ram_1_58 : _GEN_1602; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1604 = 7'h3b == index[6:0] ? ram_1_59 : _GEN_1603; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1605 = 7'h3c == index[6:0] ? ram_1_60 : _GEN_1604; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1606 = 7'h3d == index[6:0] ? ram_1_61 : _GEN_1605; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1607 = 7'h3e == index[6:0] ? ram_1_62 : _GEN_1606; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1608 = 7'h3f == index[6:0] ? ram_1_63 : _GEN_1607; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1609 = 7'h40 == index[6:0] ? ram_1_64 : _GEN_1608; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1610 = 7'h41 == index[6:0] ? ram_1_65 : _GEN_1609; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1611 = 7'h42 == index[6:0] ? ram_1_66 : _GEN_1610; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1612 = 7'h43 == index[6:0] ? ram_1_67 : _GEN_1611; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1613 = 7'h44 == index[6:0] ? ram_1_68 : _GEN_1612; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1614 = 7'h45 == index[6:0] ? ram_1_69 : _GEN_1613; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1615 = 7'h46 == index[6:0] ? ram_1_70 : _GEN_1614; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1616 = 7'h47 == index[6:0] ? ram_1_71 : _GEN_1615; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1617 = 7'h48 == index[6:0] ? ram_1_72 : _GEN_1616; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1618 = 7'h49 == index[6:0] ? ram_1_73 : _GEN_1617; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1619 = 7'h4a == index[6:0] ? ram_1_74 : _GEN_1618; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1620 = 7'h4b == index[6:0] ? ram_1_75 : _GEN_1619; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1621 = 7'h4c == index[6:0] ? ram_1_76 : _GEN_1620; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1622 = 7'h4d == index[6:0] ? ram_1_77 : _GEN_1621; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1623 = 7'h4e == index[6:0] ? ram_1_78 : _GEN_1622; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1624 = 7'h4f == index[6:0] ? ram_1_79 : _GEN_1623; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1625 = 7'h50 == index[6:0] ? ram_1_80 : _GEN_1624; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1626 = 7'h51 == index[6:0] ? ram_1_81 : _GEN_1625; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1627 = 7'h52 == index[6:0] ? ram_1_82 : _GEN_1626; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1628 = 7'h53 == index[6:0] ? ram_1_83 : _GEN_1627; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1629 = 7'h54 == index[6:0] ? ram_1_84 : _GEN_1628; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1630 = 7'h55 == index[6:0] ? ram_1_85 : _GEN_1629; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1631 = 7'h56 == index[6:0] ? ram_1_86 : _GEN_1630; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1632 = 7'h57 == index[6:0] ? ram_1_87 : _GEN_1631; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1633 = 7'h58 == index[6:0] ? ram_1_88 : _GEN_1632; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1634 = 7'h59 == index[6:0] ? ram_1_89 : _GEN_1633; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1635 = 7'h5a == index[6:0] ? ram_1_90 : _GEN_1634; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1636 = 7'h5b == index[6:0] ? ram_1_91 : _GEN_1635; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1637 = 7'h5c == index[6:0] ? ram_1_92 : _GEN_1636; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1638 = 7'h5d == index[6:0] ? ram_1_93 : _GEN_1637; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1639 = 7'h5e == index[6:0] ? ram_1_94 : _GEN_1638; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1640 = 7'h5f == index[6:0] ? ram_1_95 : _GEN_1639; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1641 = 7'h60 == index[6:0] ? ram_1_96 : _GEN_1640; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1642 = 7'h61 == index[6:0] ? ram_1_97 : _GEN_1641; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1643 = 7'h62 == index[6:0] ? ram_1_98 : _GEN_1642; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1644 = 7'h63 == index[6:0] ? ram_1_99 : _GEN_1643; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1645 = 7'h64 == index[6:0] ? ram_1_100 : _GEN_1644; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1646 = 7'h65 == index[6:0] ? ram_1_101 : _GEN_1645; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1647 = 7'h66 == index[6:0] ? ram_1_102 : _GEN_1646; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1648 = 7'h67 == index[6:0] ? ram_1_103 : _GEN_1647; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1649 = 7'h68 == index[6:0] ? ram_1_104 : _GEN_1648; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1650 = 7'h69 == index[6:0] ? ram_1_105 : _GEN_1649; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1651 = 7'h6a == index[6:0] ? ram_1_106 : _GEN_1650; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1652 = 7'h6b == index[6:0] ? ram_1_107 : _GEN_1651; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1653 = 7'h6c == index[6:0] ? ram_1_108 : _GEN_1652; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1654 = 7'h6d == index[6:0] ? ram_1_109 : _GEN_1653; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1655 = 7'h6e == index[6:0] ? ram_1_110 : _GEN_1654; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1656 = 7'h6f == index[6:0] ? ram_1_111 : _GEN_1655; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1657 = 7'h70 == index[6:0] ? ram_1_112 : _GEN_1656; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1658 = 7'h71 == index[6:0] ? ram_1_113 : _GEN_1657; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1659 = 7'h72 == index[6:0] ? ram_1_114 : _GEN_1658; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1660 = 7'h73 == index[6:0] ? ram_1_115 : _GEN_1659; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1661 = 7'h74 == index[6:0] ? ram_1_116 : _GEN_1660; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1662 = 7'h75 == index[6:0] ? ram_1_117 : _GEN_1661; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1663 = 7'h76 == index[6:0] ? ram_1_118 : _GEN_1662; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1664 = 7'h77 == index[6:0] ? ram_1_119 : _GEN_1663; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1665 = 7'h78 == index[6:0] ? ram_1_120 : _GEN_1664; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1666 = 7'h79 == index[6:0] ? ram_1_121 : _GEN_1665; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1667 = 7'h7a == index[6:0] ? ram_1_122 : _GEN_1666; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1668 = 7'h7b == index[6:0] ? ram_1_123 : _GEN_1667; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1669 = 7'h7c == index[6:0] ? ram_1_124 : _GEN_1668; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1670 = 7'h7d == index[6:0] ? ram_1_125 : _GEN_1669; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1671 = 7'h7e == index[6:0] ? ram_1_126 : _GEN_1670; // @[d_cache.scala 117:{92,92}]
  wire [63:0] _GEN_1672 = 7'h7f == index[6:0] ? ram_1_127 : _GEN_1671; // @[d_cache.scala 117:{92,92}]
  wire [126:0] _GEN_18599 = {{63'd0}, _GEN_1672}; // @[d_cache.scala 117:92]
  wire [126:0] _ram_1_T_5 = _GEN_18599 & _ram_0_T_4; // @[d_cache.scala 117:92]
  wire [126:0] _ram_1_T_6 = _ram_0_T_1 | _ram_1_T_5; // @[d_cache.scala 117:76]
  wire [63:0] _GEN_1673 = 7'h0 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_0; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1674 = 7'h1 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_1; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1675 = 7'h2 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_2; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1676 = 7'h3 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_3; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1677 = 7'h4 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_4; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1678 = 7'h5 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_5; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1679 = 7'h6 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_6; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1680 = 7'h7 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_7; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1681 = 7'h8 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_8; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1682 = 7'h9 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_9; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1683 = 7'ha == index[6:0] ? _ram_1_T_6[63:0] : ram_1_10; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1684 = 7'hb == index[6:0] ? _ram_1_T_6[63:0] : ram_1_11; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1685 = 7'hc == index[6:0] ? _ram_1_T_6[63:0] : ram_1_12; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1686 = 7'hd == index[6:0] ? _ram_1_T_6[63:0] : ram_1_13; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1687 = 7'he == index[6:0] ? _ram_1_T_6[63:0] : ram_1_14; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1688 = 7'hf == index[6:0] ? _ram_1_T_6[63:0] : ram_1_15; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1689 = 7'h10 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_16; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1690 = 7'h11 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_17; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1691 = 7'h12 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_18; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1692 = 7'h13 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_19; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1693 = 7'h14 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_20; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1694 = 7'h15 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_21; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1695 = 7'h16 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_22; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1696 = 7'h17 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_23; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1697 = 7'h18 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_24; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1698 = 7'h19 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_25; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1699 = 7'h1a == index[6:0] ? _ram_1_T_6[63:0] : ram_1_26; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1700 = 7'h1b == index[6:0] ? _ram_1_T_6[63:0] : ram_1_27; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1701 = 7'h1c == index[6:0] ? _ram_1_T_6[63:0] : ram_1_28; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1702 = 7'h1d == index[6:0] ? _ram_1_T_6[63:0] : ram_1_29; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1703 = 7'h1e == index[6:0] ? _ram_1_T_6[63:0] : ram_1_30; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1704 = 7'h1f == index[6:0] ? _ram_1_T_6[63:0] : ram_1_31; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1705 = 7'h20 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_32; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1706 = 7'h21 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_33; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1707 = 7'h22 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_34; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1708 = 7'h23 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_35; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1709 = 7'h24 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_36; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1710 = 7'h25 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_37; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1711 = 7'h26 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_38; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1712 = 7'h27 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_39; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1713 = 7'h28 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_40; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1714 = 7'h29 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_41; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1715 = 7'h2a == index[6:0] ? _ram_1_T_6[63:0] : ram_1_42; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1716 = 7'h2b == index[6:0] ? _ram_1_T_6[63:0] : ram_1_43; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1717 = 7'h2c == index[6:0] ? _ram_1_T_6[63:0] : ram_1_44; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1718 = 7'h2d == index[6:0] ? _ram_1_T_6[63:0] : ram_1_45; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1719 = 7'h2e == index[6:0] ? _ram_1_T_6[63:0] : ram_1_46; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1720 = 7'h2f == index[6:0] ? _ram_1_T_6[63:0] : ram_1_47; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1721 = 7'h30 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_48; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1722 = 7'h31 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_49; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1723 = 7'h32 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_50; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1724 = 7'h33 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_51; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1725 = 7'h34 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_52; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1726 = 7'h35 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_53; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1727 = 7'h36 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_54; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1728 = 7'h37 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_55; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1729 = 7'h38 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_56; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1730 = 7'h39 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_57; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1731 = 7'h3a == index[6:0] ? _ram_1_T_6[63:0] : ram_1_58; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1732 = 7'h3b == index[6:0] ? _ram_1_T_6[63:0] : ram_1_59; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1733 = 7'h3c == index[6:0] ? _ram_1_T_6[63:0] : ram_1_60; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1734 = 7'h3d == index[6:0] ? _ram_1_T_6[63:0] : ram_1_61; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1735 = 7'h3e == index[6:0] ? _ram_1_T_6[63:0] : ram_1_62; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1736 = 7'h3f == index[6:0] ? _ram_1_T_6[63:0] : ram_1_63; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1737 = 7'h40 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_64; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1738 = 7'h41 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_65; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1739 = 7'h42 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_66; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1740 = 7'h43 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_67; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1741 = 7'h44 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_68; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1742 = 7'h45 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_69; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1743 = 7'h46 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_70; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1744 = 7'h47 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_71; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1745 = 7'h48 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_72; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1746 = 7'h49 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_73; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1747 = 7'h4a == index[6:0] ? _ram_1_T_6[63:0] : ram_1_74; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1748 = 7'h4b == index[6:0] ? _ram_1_T_6[63:0] : ram_1_75; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1749 = 7'h4c == index[6:0] ? _ram_1_T_6[63:0] : ram_1_76; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1750 = 7'h4d == index[6:0] ? _ram_1_T_6[63:0] : ram_1_77; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1751 = 7'h4e == index[6:0] ? _ram_1_T_6[63:0] : ram_1_78; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1752 = 7'h4f == index[6:0] ? _ram_1_T_6[63:0] : ram_1_79; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1753 = 7'h50 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_80; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1754 = 7'h51 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_81; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1755 = 7'h52 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_82; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1756 = 7'h53 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_83; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1757 = 7'h54 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_84; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1758 = 7'h55 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_85; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1759 = 7'h56 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_86; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1760 = 7'h57 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_87; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1761 = 7'h58 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_88; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1762 = 7'h59 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_89; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1763 = 7'h5a == index[6:0] ? _ram_1_T_6[63:0] : ram_1_90; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1764 = 7'h5b == index[6:0] ? _ram_1_T_6[63:0] : ram_1_91; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1765 = 7'h5c == index[6:0] ? _ram_1_T_6[63:0] : ram_1_92; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1766 = 7'h5d == index[6:0] ? _ram_1_T_6[63:0] : ram_1_93; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1767 = 7'h5e == index[6:0] ? _ram_1_T_6[63:0] : ram_1_94; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1768 = 7'h5f == index[6:0] ? _ram_1_T_6[63:0] : ram_1_95; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1769 = 7'h60 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_96; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1770 = 7'h61 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_97; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1771 = 7'h62 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_98; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1772 = 7'h63 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_99; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1773 = 7'h64 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_100; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1774 = 7'h65 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_101; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1775 = 7'h66 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_102; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1776 = 7'h67 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_103; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1777 = 7'h68 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_104; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1778 = 7'h69 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_105; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1779 = 7'h6a == index[6:0] ? _ram_1_T_6[63:0] : ram_1_106; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1780 = 7'h6b == index[6:0] ? _ram_1_T_6[63:0] : ram_1_107; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1781 = 7'h6c == index[6:0] ? _ram_1_T_6[63:0] : ram_1_108; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1782 = 7'h6d == index[6:0] ? _ram_1_T_6[63:0] : ram_1_109; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1783 = 7'h6e == index[6:0] ? _ram_1_T_6[63:0] : ram_1_110; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1784 = 7'h6f == index[6:0] ? _ram_1_T_6[63:0] : ram_1_111; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1785 = 7'h70 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_112; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1786 = 7'h71 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_113; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1787 = 7'h72 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_114; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1788 = 7'h73 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_115; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1789 = 7'h74 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_116; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1790 = 7'h75 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_117; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1791 = 7'h76 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_118; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1792 = 7'h77 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_119; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1793 = 7'h78 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_120; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1794 = 7'h79 == index[6:0] ? _ram_1_T_6[63:0] : ram_1_121; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1795 = 7'h7a == index[6:0] ? _ram_1_T_6[63:0] : ram_1_122; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1796 = 7'h7b == index[6:0] ? _ram_1_T_6[63:0] : ram_1_123; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1797 = 7'h7c == index[6:0] ? _ram_1_T_6[63:0] : ram_1_124; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1798 = 7'h7d == index[6:0] ? _ram_1_T_6[63:0] : ram_1_125; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1799 = 7'h7e == index[6:0] ? _ram_1_T_6[63:0] : ram_1_126; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1800 = 7'h7f == index[6:0] ? _ram_1_T_6[63:0] : ram_1_127; // @[d_cache.scala 117:{30,30} 19:24]
  wire [63:0] _GEN_1801 = 7'h0 == index[6:0] ? _ram_0_T : recent_wdata1_0; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1802 = 7'h1 == index[6:0] ? _ram_0_T : recent_wdata1_1; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1803 = 7'h2 == index[6:0] ? _ram_0_T : recent_wdata1_2; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1804 = 7'h3 == index[6:0] ? _ram_0_T : recent_wdata1_3; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1805 = 7'h4 == index[6:0] ? _ram_0_T : recent_wdata1_4; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1806 = 7'h5 == index[6:0] ? _ram_0_T : recent_wdata1_5; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1807 = 7'h6 == index[6:0] ? _ram_0_T : recent_wdata1_6; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1808 = 7'h7 == index[6:0] ? _ram_0_T : recent_wdata1_7; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1809 = 7'h8 == index[6:0] ? _ram_0_T : recent_wdata1_8; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1810 = 7'h9 == index[6:0] ? _ram_0_T : recent_wdata1_9; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1811 = 7'ha == index[6:0] ? _ram_0_T : recent_wdata1_10; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1812 = 7'hb == index[6:0] ? _ram_0_T : recent_wdata1_11; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1813 = 7'hc == index[6:0] ? _ram_0_T : recent_wdata1_12; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1814 = 7'hd == index[6:0] ? _ram_0_T : recent_wdata1_13; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1815 = 7'he == index[6:0] ? _ram_0_T : recent_wdata1_14; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1816 = 7'hf == index[6:0] ? _ram_0_T : recent_wdata1_15; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1817 = 7'h10 == index[6:0] ? _ram_0_T : recent_wdata1_16; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1818 = 7'h11 == index[6:0] ? _ram_0_T : recent_wdata1_17; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1819 = 7'h12 == index[6:0] ? _ram_0_T : recent_wdata1_18; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1820 = 7'h13 == index[6:0] ? _ram_0_T : recent_wdata1_19; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1821 = 7'h14 == index[6:0] ? _ram_0_T : recent_wdata1_20; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1822 = 7'h15 == index[6:0] ? _ram_0_T : recent_wdata1_21; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1823 = 7'h16 == index[6:0] ? _ram_0_T : recent_wdata1_22; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1824 = 7'h17 == index[6:0] ? _ram_0_T : recent_wdata1_23; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1825 = 7'h18 == index[6:0] ? _ram_0_T : recent_wdata1_24; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1826 = 7'h19 == index[6:0] ? _ram_0_T : recent_wdata1_25; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1827 = 7'h1a == index[6:0] ? _ram_0_T : recent_wdata1_26; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1828 = 7'h1b == index[6:0] ? _ram_0_T : recent_wdata1_27; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1829 = 7'h1c == index[6:0] ? _ram_0_T : recent_wdata1_28; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1830 = 7'h1d == index[6:0] ? _ram_0_T : recent_wdata1_29; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1831 = 7'h1e == index[6:0] ? _ram_0_T : recent_wdata1_30; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1832 = 7'h1f == index[6:0] ? _ram_0_T : recent_wdata1_31; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1833 = 7'h20 == index[6:0] ? _ram_0_T : recent_wdata1_32; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1834 = 7'h21 == index[6:0] ? _ram_0_T : recent_wdata1_33; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1835 = 7'h22 == index[6:0] ? _ram_0_T : recent_wdata1_34; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1836 = 7'h23 == index[6:0] ? _ram_0_T : recent_wdata1_35; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1837 = 7'h24 == index[6:0] ? _ram_0_T : recent_wdata1_36; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1838 = 7'h25 == index[6:0] ? _ram_0_T : recent_wdata1_37; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1839 = 7'h26 == index[6:0] ? _ram_0_T : recent_wdata1_38; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1840 = 7'h27 == index[6:0] ? _ram_0_T : recent_wdata1_39; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1841 = 7'h28 == index[6:0] ? _ram_0_T : recent_wdata1_40; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1842 = 7'h29 == index[6:0] ? _ram_0_T : recent_wdata1_41; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1843 = 7'h2a == index[6:0] ? _ram_0_T : recent_wdata1_42; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1844 = 7'h2b == index[6:0] ? _ram_0_T : recent_wdata1_43; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1845 = 7'h2c == index[6:0] ? _ram_0_T : recent_wdata1_44; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1846 = 7'h2d == index[6:0] ? _ram_0_T : recent_wdata1_45; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1847 = 7'h2e == index[6:0] ? _ram_0_T : recent_wdata1_46; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1848 = 7'h2f == index[6:0] ? _ram_0_T : recent_wdata1_47; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1849 = 7'h30 == index[6:0] ? _ram_0_T : recent_wdata1_48; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1850 = 7'h31 == index[6:0] ? _ram_0_T : recent_wdata1_49; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1851 = 7'h32 == index[6:0] ? _ram_0_T : recent_wdata1_50; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1852 = 7'h33 == index[6:0] ? _ram_0_T : recent_wdata1_51; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1853 = 7'h34 == index[6:0] ? _ram_0_T : recent_wdata1_52; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1854 = 7'h35 == index[6:0] ? _ram_0_T : recent_wdata1_53; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1855 = 7'h36 == index[6:0] ? _ram_0_T : recent_wdata1_54; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1856 = 7'h37 == index[6:0] ? _ram_0_T : recent_wdata1_55; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1857 = 7'h38 == index[6:0] ? _ram_0_T : recent_wdata1_56; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1858 = 7'h39 == index[6:0] ? _ram_0_T : recent_wdata1_57; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1859 = 7'h3a == index[6:0] ? _ram_0_T : recent_wdata1_58; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1860 = 7'h3b == index[6:0] ? _ram_0_T : recent_wdata1_59; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1861 = 7'h3c == index[6:0] ? _ram_0_T : recent_wdata1_60; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1862 = 7'h3d == index[6:0] ? _ram_0_T : recent_wdata1_61; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1863 = 7'h3e == index[6:0] ? _ram_0_T : recent_wdata1_62; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1864 = 7'h3f == index[6:0] ? _ram_0_T : recent_wdata1_63; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1865 = 7'h40 == index[6:0] ? _ram_0_T : recent_wdata1_64; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1866 = 7'h41 == index[6:0] ? _ram_0_T : recent_wdata1_65; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1867 = 7'h42 == index[6:0] ? _ram_0_T : recent_wdata1_66; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1868 = 7'h43 == index[6:0] ? _ram_0_T : recent_wdata1_67; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1869 = 7'h44 == index[6:0] ? _ram_0_T : recent_wdata1_68; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1870 = 7'h45 == index[6:0] ? _ram_0_T : recent_wdata1_69; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1871 = 7'h46 == index[6:0] ? _ram_0_T : recent_wdata1_70; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1872 = 7'h47 == index[6:0] ? _ram_0_T : recent_wdata1_71; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1873 = 7'h48 == index[6:0] ? _ram_0_T : recent_wdata1_72; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1874 = 7'h49 == index[6:0] ? _ram_0_T : recent_wdata1_73; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1875 = 7'h4a == index[6:0] ? _ram_0_T : recent_wdata1_74; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1876 = 7'h4b == index[6:0] ? _ram_0_T : recent_wdata1_75; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1877 = 7'h4c == index[6:0] ? _ram_0_T : recent_wdata1_76; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1878 = 7'h4d == index[6:0] ? _ram_0_T : recent_wdata1_77; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1879 = 7'h4e == index[6:0] ? _ram_0_T : recent_wdata1_78; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1880 = 7'h4f == index[6:0] ? _ram_0_T : recent_wdata1_79; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1881 = 7'h50 == index[6:0] ? _ram_0_T : recent_wdata1_80; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1882 = 7'h51 == index[6:0] ? _ram_0_T : recent_wdata1_81; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1883 = 7'h52 == index[6:0] ? _ram_0_T : recent_wdata1_82; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1884 = 7'h53 == index[6:0] ? _ram_0_T : recent_wdata1_83; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1885 = 7'h54 == index[6:0] ? _ram_0_T : recent_wdata1_84; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1886 = 7'h55 == index[6:0] ? _ram_0_T : recent_wdata1_85; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1887 = 7'h56 == index[6:0] ? _ram_0_T : recent_wdata1_86; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1888 = 7'h57 == index[6:0] ? _ram_0_T : recent_wdata1_87; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1889 = 7'h58 == index[6:0] ? _ram_0_T : recent_wdata1_88; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1890 = 7'h59 == index[6:0] ? _ram_0_T : recent_wdata1_89; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1891 = 7'h5a == index[6:0] ? _ram_0_T : recent_wdata1_90; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1892 = 7'h5b == index[6:0] ? _ram_0_T : recent_wdata1_91; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1893 = 7'h5c == index[6:0] ? _ram_0_T : recent_wdata1_92; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1894 = 7'h5d == index[6:0] ? _ram_0_T : recent_wdata1_93; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1895 = 7'h5e == index[6:0] ? _ram_0_T : recent_wdata1_94; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1896 = 7'h5f == index[6:0] ? _ram_0_T : recent_wdata1_95; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1897 = 7'h60 == index[6:0] ? _ram_0_T : recent_wdata1_96; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1898 = 7'h61 == index[6:0] ? _ram_0_T : recent_wdata1_97; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1899 = 7'h62 == index[6:0] ? _ram_0_T : recent_wdata1_98; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1900 = 7'h63 == index[6:0] ? _ram_0_T : recent_wdata1_99; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1901 = 7'h64 == index[6:0] ? _ram_0_T : recent_wdata1_100; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1902 = 7'h65 == index[6:0] ? _ram_0_T : recent_wdata1_101; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1903 = 7'h66 == index[6:0] ? _ram_0_T : recent_wdata1_102; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1904 = 7'h67 == index[6:0] ? _ram_0_T : recent_wdata1_103; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1905 = 7'h68 == index[6:0] ? _ram_0_T : recent_wdata1_104; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1906 = 7'h69 == index[6:0] ? _ram_0_T : recent_wdata1_105; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1907 = 7'h6a == index[6:0] ? _ram_0_T : recent_wdata1_106; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1908 = 7'h6b == index[6:0] ? _ram_0_T : recent_wdata1_107; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1909 = 7'h6c == index[6:0] ? _ram_0_T : recent_wdata1_108; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1910 = 7'h6d == index[6:0] ? _ram_0_T : recent_wdata1_109; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1911 = 7'h6e == index[6:0] ? _ram_0_T : recent_wdata1_110; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1912 = 7'h6f == index[6:0] ? _ram_0_T : recent_wdata1_111; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1913 = 7'h70 == index[6:0] ? _ram_0_T : recent_wdata1_112; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1914 = 7'h71 == index[6:0] ? _ram_0_T : recent_wdata1_113; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1915 = 7'h72 == index[6:0] ? _ram_0_T : recent_wdata1_114; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1916 = 7'h73 == index[6:0] ? _ram_0_T : recent_wdata1_115; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1917 = 7'h74 == index[6:0] ? _ram_0_T : recent_wdata1_116; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1918 = 7'h75 == index[6:0] ? _ram_0_T : recent_wdata1_117; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1919 = 7'h76 == index[6:0] ? _ram_0_T : recent_wdata1_118; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1920 = 7'h77 == index[6:0] ? _ram_0_T : recent_wdata1_119; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1921 = 7'h78 == index[6:0] ? _ram_0_T : recent_wdata1_120; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1922 = 7'h79 == index[6:0] ? _ram_0_T : recent_wdata1_121; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1923 = 7'h7a == index[6:0] ? _ram_0_T : recent_wdata1_122; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1924 = 7'h7b == index[6:0] ? _ram_0_T : recent_wdata1_123; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1925 = 7'h7c == index[6:0] ? _ram_0_T : recent_wdata1_124; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1926 = 7'h7d == index[6:0] ? _ram_0_T : recent_wdata1_125; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1927 = 7'h7e == index[6:0] ? _ram_0_T : recent_wdata1_126; // @[d_cache.scala 119:{38,38} 21:32]
  wire [63:0] _GEN_1928 = 7'h7f == index[6:0] ? _ram_0_T : recent_wdata1_127; // @[d_cache.scala 119:{38,38} 21:32]
  wire  _GEN_1929 = _GEN_18470 | dirty_1_0; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1930 = _GEN_18471 | dirty_1_1; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1931 = _GEN_18472 | dirty_1_2; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1932 = _GEN_18473 | dirty_1_3; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1933 = _GEN_18474 | dirty_1_4; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1934 = _GEN_18475 | dirty_1_5; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1935 = _GEN_18476 | dirty_1_6; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1936 = _GEN_18477 | dirty_1_7; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1937 = _GEN_18478 | dirty_1_8; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1938 = _GEN_18479 | dirty_1_9; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1939 = _GEN_18480 | dirty_1_10; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1940 = _GEN_18481 | dirty_1_11; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1941 = _GEN_18482 | dirty_1_12; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1942 = _GEN_18483 | dirty_1_13; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1943 = _GEN_18484 | dirty_1_14; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1944 = _GEN_18485 | dirty_1_15; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1945 = _GEN_18486 | dirty_1_16; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1946 = _GEN_18487 | dirty_1_17; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1947 = _GEN_18488 | dirty_1_18; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1948 = _GEN_18489 | dirty_1_19; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1949 = _GEN_18490 | dirty_1_20; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1950 = _GEN_18491 | dirty_1_21; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1951 = _GEN_18492 | dirty_1_22; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1952 = _GEN_18493 | dirty_1_23; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1953 = _GEN_18494 | dirty_1_24; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1954 = _GEN_18495 | dirty_1_25; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1955 = _GEN_18496 | dirty_1_26; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1956 = _GEN_18497 | dirty_1_27; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1957 = _GEN_18498 | dirty_1_28; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1958 = _GEN_18499 | dirty_1_29; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1959 = _GEN_18500 | dirty_1_30; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1960 = _GEN_18501 | dirty_1_31; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1961 = _GEN_18502 | dirty_1_32; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1962 = _GEN_18503 | dirty_1_33; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1963 = _GEN_18504 | dirty_1_34; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1964 = _GEN_18505 | dirty_1_35; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1965 = _GEN_18506 | dirty_1_36; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1966 = _GEN_18507 | dirty_1_37; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1967 = _GEN_18508 | dirty_1_38; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1968 = _GEN_18509 | dirty_1_39; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1969 = _GEN_18510 | dirty_1_40; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1970 = _GEN_18511 | dirty_1_41; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1971 = _GEN_18512 | dirty_1_42; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1972 = _GEN_18513 | dirty_1_43; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1973 = _GEN_18514 | dirty_1_44; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1974 = _GEN_18515 | dirty_1_45; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1975 = _GEN_18516 | dirty_1_46; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1976 = _GEN_18517 | dirty_1_47; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1977 = _GEN_18518 | dirty_1_48; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1978 = _GEN_18519 | dirty_1_49; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1979 = _GEN_18520 | dirty_1_50; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1980 = _GEN_18521 | dirty_1_51; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1981 = _GEN_18522 | dirty_1_52; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1982 = _GEN_18523 | dirty_1_53; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1983 = _GEN_18524 | dirty_1_54; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1984 = _GEN_18525 | dirty_1_55; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1985 = _GEN_18526 | dirty_1_56; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1986 = _GEN_18527 | dirty_1_57; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1987 = _GEN_18528 | dirty_1_58; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1988 = _GEN_18529 | dirty_1_59; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1989 = _GEN_18530 | dirty_1_60; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1990 = _GEN_18531 | dirty_1_61; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1991 = _GEN_18532 | dirty_1_62; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1992 = _GEN_18533 | dirty_1_63; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1993 = _GEN_18534 | dirty_1_64; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1994 = _GEN_18535 | dirty_1_65; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1995 = _GEN_18536 | dirty_1_66; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1996 = _GEN_18537 | dirty_1_67; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1997 = _GEN_18538 | dirty_1_68; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1998 = _GEN_18539 | dirty_1_69; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_1999 = _GEN_18540 | dirty_1_70; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2000 = _GEN_18541 | dirty_1_71; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2001 = _GEN_18542 | dirty_1_72; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2002 = _GEN_18543 | dirty_1_73; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2003 = _GEN_18544 | dirty_1_74; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2004 = _GEN_18545 | dirty_1_75; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2005 = _GEN_18546 | dirty_1_76; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2006 = _GEN_18547 | dirty_1_77; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2007 = _GEN_18548 | dirty_1_78; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2008 = _GEN_18549 | dirty_1_79; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2009 = _GEN_18550 | dirty_1_80; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2010 = _GEN_18551 | dirty_1_81; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2011 = _GEN_18552 | dirty_1_82; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2012 = _GEN_18553 | dirty_1_83; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2013 = _GEN_18554 | dirty_1_84; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2014 = _GEN_18555 | dirty_1_85; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2015 = _GEN_18556 | dirty_1_86; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2016 = _GEN_18557 | dirty_1_87; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2017 = _GEN_18558 | dirty_1_88; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2018 = _GEN_18559 | dirty_1_89; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2019 = _GEN_18560 | dirty_1_90; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2020 = _GEN_18561 | dirty_1_91; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2021 = _GEN_18562 | dirty_1_92; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2022 = _GEN_18563 | dirty_1_93; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2023 = _GEN_18564 | dirty_1_94; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2024 = _GEN_18565 | dirty_1_95; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2025 = _GEN_18566 | dirty_1_96; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2026 = _GEN_18567 | dirty_1_97; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2027 = _GEN_18568 | dirty_1_98; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2028 = _GEN_18569 | dirty_1_99; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2029 = _GEN_18570 | dirty_1_100; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2030 = _GEN_18571 | dirty_1_101; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2031 = _GEN_18572 | dirty_1_102; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2032 = _GEN_18573 | dirty_1_103; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2033 = _GEN_18574 | dirty_1_104; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2034 = _GEN_18575 | dirty_1_105; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2035 = _GEN_18576 | dirty_1_106; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2036 = _GEN_18577 | dirty_1_107; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2037 = _GEN_18578 | dirty_1_108; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2038 = _GEN_18579 | dirty_1_109; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2039 = _GEN_18580 | dirty_1_110; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2040 = _GEN_18581 | dirty_1_111; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2041 = _GEN_18582 | dirty_1_112; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2042 = _GEN_18583 | dirty_1_113; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2043 = _GEN_18584 | dirty_1_114; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2044 = _GEN_18585 | dirty_1_115; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2045 = _GEN_18586 | dirty_1_116; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2046 = _GEN_18587 | dirty_1_117; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2047 = _GEN_18588 | dirty_1_118; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2048 = _GEN_18589 | dirty_1_119; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2049 = _GEN_18590 | dirty_1_120; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2050 = _GEN_18591 | dirty_1_121; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2051 = _GEN_18592 | dirty_1_122; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2052 = _GEN_18593 | dirty_1_123; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2053 = _GEN_18594 | dirty_1_124; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2054 = _GEN_18595 | dirty_1_125; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2055 = _GEN_18596 | dirty_1_126; // @[d_cache.scala 120:{32,32} 27:26]
  wire  _GEN_2056 = _GEN_18597 | dirty_1_127; // @[d_cache.scala 120:{32,32} 27:26]
  wire [2:0] _GEN_2057 = way1_hit ? 3'h0 : 3'h4; // @[d_cache.scala 115:33 116:23 122:23]
  wire [63:0] _GEN_2058 = way1_hit ? _GEN_1673 : ram_1_0; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2059 = way1_hit ? _GEN_1674 : ram_1_1; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2060 = way1_hit ? _GEN_1675 : ram_1_2; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2061 = way1_hit ? _GEN_1676 : ram_1_3; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2062 = way1_hit ? _GEN_1677 : ram_1_4; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2063 = way1_hit ? _GEN_1678 : ram_1_5; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2064 = way1_hit ? _GEN_1679 : ram_1_6; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2065 = way1_hit ? _GEN_1680 : ram_1_7; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2066 = way1_hit ? _GEN_1681 : ram_1_8; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2067 = way1_hit ? _GEN_1682 : ram_1_9; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2068 = way1_hit ? _GEN_1683 : ram_1_10; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2069 = way1_hit ? _GEN_1684 : ram_1_11; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2070 = way1_hit ? _GEN_1685 : ram_1_12; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2071 = way1_hit ? _GEN_1686 : ram_1_13; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2072 = way1_hit ? _GEN_1687 : ram_1_14; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2073 = way1_hit ? _GEN_1688 : ram_1_15; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2074 = way1_hit ? _GEN_1689 : ram_1_16; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2075 = way1_hit ? _GEN_1690 : ram_1_17; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2076 = way1_hit ? _GEN_1691 : ram_1_18; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2077 = way1_hit ? _GEN_1692 : ram_1_19; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2078 = way1_hit ? _GEN_1693 : ram_1_20; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2079 = way1_hit ? _GEN_1694 : ram_1_21; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2080 = way1_hit ? _GEN_1695 : ram_1_22; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2081 = way1_hit ? _GEN_1696 : ram_1_23; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2082 = way1_hit ? _GEN_1697 : ram_1_24; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2083 = way1_hit ? _GEN_1698 : ram_1_25; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2084 = way1_hit ? _GEN_1699 : ram_1_26; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2085 = way1_hit ? _GEN_1700 : ram_1_27; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2086 = way1_hit ? _GEN_1701 : ram_1_28; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2087 = way1_hit ? _GEN_1702 : ram_1_29; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2088 = way1_hit ? _GEN_1703 : ram_1_30; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2089 = way1_hit ? _GEN_1704 : ram_1_31; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2090 = way1_hit ? _GEN_1705 : ram_1_32; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2091 = way1_hit ? _GEN_1706 : ram_1_33; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2092 = way1_hit ? _GEN_1707 : ram_1_34; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2093 = way1_hit ? _GEN_1708 : ram_1_35; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2094 = way1_hit ? _GEN_1709 : ram_1_36; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2095 = way1_hit ? _GEN_1710 : ram_1_37; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2096 = way1_hit ? _GEN_1711 : ram_1_38; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2097 = way1_hit ? _GEN_1712 : ram_1_39; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2098 = way1_hit ? _GEN_1713 : ram_1_40; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2099 = way1_hit ? _GEN_1714 : ram_1_41; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2100 = way1_hit ? _GEN_1715 : ram_1_42; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2101 = way1_hit ? _GEN_1716 : ram_1_43; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2102 = way1_hit ? _GEN_1717 : ram_1_44; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2103 = way1_hit ? _GEN_1718 : ram_1_45; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2104 = way1_hit ? _GEN_1719 : ram_1_46; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2105 = way1_hit ? _GEN_1720 : ram_1_47; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2106 = way1_hit ? _GEN_1721 : ram_1_48; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2107 = way1_hit ? _GEN_1722 : ram_1_49; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2108 = way1_hit ? _GEN_1723 : ram_1_50; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2109 = way1_hit ? _GEN_1724 : ram_1_51; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2110 = way1_hit ? _GEN_1725 : ram_1_52; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2111 = way1_hit ? _GEN_1726 : ram_1_53; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2112 = way1_hit ? _GEN_1727 : ram_1_54; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2113 = way1_hit ? _GEN_1728 : ram_1_55; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2114 = way1_hit ? _GEN_1729 : ram_1_56; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2115 = way1_hit ? _GEN_1730 : ram_1_57; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2116 = way1_hit ? _GEN_1731 : ram_1_58; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2117 = way1_hit ? _GEN_1732 : ram_1_59; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2118 = way1_hit ? _GEN_1733 : ram_1_60; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2119 = way1_hit ? _GEN_1734 : ram_1_61; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2120 = way1_hit ? _GEN_1735 : ram_1_62; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2121 = way1_hit ? _GEN_1736 : ram_1_63; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2122 = way1_hit ? _GEN_1737 : ram_1_64; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2123 = way1_hit ? _GEN_1738 : ram_1_65; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2124 = way1_hit ? _GEN_1739 : ram_1_66; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2125 = way1_hit ? _GEN_1740 : ram_1_67; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2126 = way1_hit ? _GEN_1741 : ram_1_68; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2127 = way1_hit ? _GEN_1742 : ram_1_69; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2128 = way1_hit ? _GEN_1743 : ram_1_70; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2129 = way1_hit ? _GEN_1744 : ram_1_71; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2130 = way1_hit ? _GEN_1745 : ram_1_72; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2131 = way1_hit ? _GEN_1746 : ram_1_73; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2132 = way1_hit ? _GEN_1747 : ram_1_74; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2133 = way1_hit ? _GEN_1748 : ram_1_75; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2134 = way1_hit ? _GEN_1749 : ram_1_76; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2135 = way1_hit ? _GEN_1750 : ram_1_77; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2136 = way1_hit ? _GEN_1751 : ram_1_78; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2137 = way1_hit ? _GEN_1752 : ram_1_79; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2138 = way1_hit ? _GEN_1753 : ram_1_80; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2139 = way1_hit ? _GEN_1754 : ram_1_81; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2140 = way1_hit ? _GEN_1755 : ram_1_82; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2141 = way1_hit ? _GEN_1756 : ram_1_83; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2142 = way1_hit ? _GEN_1757 : ram_1_84; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2143 = way1_hit ? _GEN_1758 : ram_1_85; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2144 = way1_hit ? _GEN_1759 : ram_1_86; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2145 = way1_hit ? _GEN_1760 : ram_1_87; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2146 = way1_hit ? _GEN_1761 : ram_1_88; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2147 = way1_hit ? _GEN_1762 : ram_1_89; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2148 = way1_hit ? _GEN_1763 : ram_1_90; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2149 = way1_hit ? _GEN_1764 : ram_1_91; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2150 = way1_hit ? _GEN_1765 : ram_1_92; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2151 = way1_hit ? _GEN_1766 : ram_1_93; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2152 = way1_hit ? _GEN_1767 : ram_1_94; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2153 = way1_hit ? _GEN_1768 : ram_1_95; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2154 = way1_hit ? _GEN_1769 : ram_1_96; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2155 = way1_hit ? _GEN_1770 : ram_1_97; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2156 = way1_hit ? _GEN_1771 : ram_1_98; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2157 = way1_hit ? _GEN_1772 : ram_1_99; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2158 = way1_hit ? _GEN_1773 : ram_1_100; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2159 = way1_hit ? _GEN_1774 : ram_1_101; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2160 = way1_hit ? _GEN_1775 : ram_1_102; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2161 = way1_hit ? _GEN_1776 : ram_1_103; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2162 = way1_hit ? _GEN_1777 : ram_1_104; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2163 = way1_hit ? _GEN_1778 : ram_1_105; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2164 = way1_hit ? _GEN_1779 : ram_1_106; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2165 = way1_hit ? _GEN_1780 : ram_1_107; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2166 = way1_hit ? _GEN_1781 : ram_1_108; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2167 = way1_hit ? _GEN_1782 : ram_1_109; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2168 = way1_hit ? _GEN_1783 : ram_1_110; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2169 = way1_hit ? _GEN_1784 : ram_1_111; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2170 = way1_hit ? _GEN_1785 : ram_1_112; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2171 = way1_hit ? _GEN_1786 : ram_1_113; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2172 = way1_hit ? _GEN_1787 : ram_1_114; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2173 = way1_hit ? _GEN_1788 : ram_1_115; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2174 = way1_hit ? _GEN_1789 : ram_1_116; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2175 = way1_hit ? _GEN_1790 : ram_1_117; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2176 = way1_hit ? _GEN_1791 : ram_1_118; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2177 = way1_hit ? _GEN_1792 : ram_1_119; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2178 = way1_hit ? _GEN_1793 : ram_1_120; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2179 = way1_hit ? _GEN_1794 : ram_1_121; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2180 = way1_hit ? _GEN_1795 : ram_1_122; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2181 = way1_hit ? _GEN_1796 : ram_1_123; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2182 = way1_hit ? _GEN_1797 : ram_1_124; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2183 = way1_hit ? _GEN_1798 : ram_1_125; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2184 = way1_hit ? _GEN_1799 : ram_1_126; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2185 = way1_hit ? _GEN_1800 : ram_1_127; // @[d_cache.scala 115:33 19:24]
  wire [63:0] _GEN_2186 = way1_hit ? _GEN_1801 : recent_wdata1_0; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2187 = way1_hit ? _GEN_1802 : recent_wdata1_1; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2188 = way1_hit ? _GEN_1803 : recent_wdata1_2; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2189 = way1_hit ? _GEN_1804 : recent_wdata1_3; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2190 = way1_hit ? _GEN_1805 : recent_wdata1_4; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2191 = way1_hit ? _GEN_1806 : recent_wdata1_5; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2192 = way1_hit ? _GEN_1807 : recent_wdata1_6; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2193 = way1_hit ? _GEN_1808 : recent_wdata1_7; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2194 = way1_hit ? _GEN_1809 : recent_wdata1_8; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2195 = way1_hit ? _GEN_1810 : recent_wdata1_9; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2196 = way1_hit ? _GEN_1811 : recent_wdata1_10; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2197 = way1_hit ? _GEN_1812 : recent_wdata1_11; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2198 = way1_hit ? _GEN_1813 : recent_wdata1_12; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2199 = way1_hit ? _GEN_1814 : recent_wdata1_13; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2200 = way1_hit ? _GEN_1815 : recent_wdata1_14; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2201 = way1_hit ? _GEN_1816 : recent_wdata1_15; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2202 = way1_hit ? _GEN_1817 : recent_wdata1_16; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2203 = way1_hit ? _GEN_1818 : recent_wdata1_17; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2204 = way1_hit ? _GEN_1819 : recent_wdata1_18; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2205 = way1_hit ? _GEN_1820 : recent_wdata1_19; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2206 = way1_hit ? _GEN_1821 : recent_wdata1_20; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2207 = way1_hit ? _GEN_1822 : recent_wdata1_21; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2208 = way1_hit ? _GEN_1823 : recent_wdata1_22; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2209 = way1_hit ? _GEN_1824 : recent_wdata1_23; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2210 = way1_hit ? _GEN_1825 : recent_wdata1_24; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2211 = way1_hit ? _GEN_1826 : recent_wdata1_25; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2212 = way1_hit ? _GEN_1827 : recent_wdata1_26; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2213 = way1_hit ? _GEN_1828 : recent_wdata1_27; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2214 = way1_hit ? _GEN_1829 : recent_wdata1_28; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2215 = way1_hit ? _GEN_1830 : recent_wdata1_29; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2216 = way1_hit ? _GEN_1831 : recent_wdata1_30; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2217 = way1_hit ? _GEN_1832 : recent_wdata1_31; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2218 = way1_hit ? _GEN_1833 : recent_wdata1_32; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2219 = way1_hit ? _GEN_1834 : recent_wdata1_33; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2220 = way1_hit ? _GEN_1835 : recent_wdata1_34; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2221 = way1_hit ? _GEN_1836 : recent_wdata1_35; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2222 = way1_hit ? _GEN_1837 : recent_wdata1_36; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2223 = way1_hit ? _GEN_1838 : recent_wdata1_37; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2224 = way1_hit ? _GEN_1839 : recent_wdata1_38; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2225 = way1_hit ? _GEN_1840 : recent_wdata1_39; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2226 = way1_hit ? _GEN_1841 : recent_wdata1_40; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2227 = way1_hit ? _GEN_1842 : recent_wdata1_41; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2228 = way1_hit ? _GEN_1843 : recent_wdata1_42; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2229 = way1_hit ? _GEN_1844 : recent_wdata1_43; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2230 = way1_hit ? _GEN_1845 : recent_wdata1_44; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2231 = way1_hit ? _GEN_1846 : recent_wdata1_45; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2232 = way1_hit ? _GEN_1847 : recent_wdata1_46; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2233 = way1_hit ? _GEN_1848 : recent_wdata1_47; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2234 = way1_hit ? _GEN_1849 : recent_wdata1_48; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2235 = way1_hit ? _GEN_1850 : recent_wdata1_49; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2236 = way1_hit ? _GEN_1851 : recent_wdata1_50; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2237 = way1_hit ? _GEN_1852 : recent_wdata1_51; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2238 = way1_hit ? _GEN_1853 : recent_wdata1_52; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2239 = way1_hit ? _GEN_1854 : recent_wdata1_53; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2240 = way1_hit ? _GEN_1855 : recent_wdata1_54; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2241 = way1_hit ? _GEN_1856 : recent_wdata1_55; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2242 = way1_hit ? _GEN_1857 : recent_wdata1_56; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2243 = way1_hit ? _GEN_1858 : recent_wdata1_57; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2244 = way1_hit ? _GEN_1859 : recent_wdata1_58; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2245 = way1_hit ? _GEN_1860 : recent_wdata1_59; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2246 = way1_hit ? _GEN_1861 : recent_wdata1_60; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2247 = way1_hit ? _GEN_1862 : recent_wdata1_61; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2248 = way1_hit ? _GEN_1863 : recent_wdata1_62; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2249 = way1_hit ? _GEN_1864 : recent_wdata1_63; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2250 = way1_hit ? _GEN_1865 : recent_wdata1_64; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2251 = way1_hit ? _GEN_1866 : recent_wdata1_65; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2252 = way1_hit ? _GEN_1867 : recent_wdata1_66; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2253 = way1_hit ? _GEN_1868 : recent_wdata1_67; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2254 = way1_hit ? _GEN_1869 : recent_wdata1_68; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2255 = way1_hit ? _GEN_1870 : recent_wdata1_69; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2256 = way1_hit ? _GEN_1871 : recent_wdata1_70; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2257 = way1_hit ? _GEN_1872 : recent_wdata1_71; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2258 = way1_hit ? _GEN_1873 : recent_wdata1_72; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2259 = way1_hit ? _GEN_1874 : recent_wdata1_73; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2260 = way1_hit ? _GEN_1875 : recent_wdata1_74; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2261 = way1_hit ? _GEN_1876 : recent_wdata1_75; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2262 = way1_hit ? _GEN_1877 : recent_wdata1_76; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2263 = way1_hit ? _GEN_1878 : recent_wdata1_77; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2264 = way1_hit ? _GEN_1879 : recent_wdata1_78; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2265 = way1_hit ? _GEN_1880 : recent_wdata1_79; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2266 = way1_hit ? _GEN_1881 : recent_wdata1_80; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2267 = way1_hit ? _GEN_1882 : recent_wdata1_81; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2268 = way1_hit ? _GEN_1883 : recent_wdata1_82; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2269 = way1_hit ? _GEN_1884 : recent_wdata1_83; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2270 = way1_hit ? _GEN_1885 : recent_wdata1_84; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2271 = way1_hit ? _GEN_1886 : recent_wdata1_85; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2272 = way1_hit ? _GEN_1887 : recent_wdata1_86; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2273 = way1_hit ? _GEN_1888 : recent_wdata1_87; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2274 = way1_hit ? _GEN_1889 : recent_wdata1_88; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2275 = way1_hit ? _GEN_1890 : recent_wdata1_89; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2276 = way1_hit ? _GEN_1891 : recent_wdata1_90; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2277 = way1_hit ? _GEN_1892 : recent_wdata1_91; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2278 = way1_hit ? _GEN_1893 : recent_wdata1_92; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2279 = way1_hit ? _GEN_1894 : recent_wdata1_93; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2280 = way1_hit ? _GEN_1895 : recent_wdata1_94; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2281 = way1_hit ? _GEN_1896 : recent_wdata1_95; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2282 = way1_hit ? _GEN_1897 : recent_wdata1_96; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2283 = way1_hit ? _GEN_1898 : recent_wdata1_97; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2284 = way1_hit ? _GEN_1899 : recent_wdata1_98; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2285 = way1_hit ? _GEN_1900 : recent_wdata1_99; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2286 = way1_hit ? _GEN_1901 : recent_wdata1_100; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2287 = way1_hit ? _GEN_1902 : recent_wdata1_101; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2288 = way1_hit ? _GEN_1903 : recent_wdata1_102; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2289 = way1_hit ? _GEN_1904 : recent_wdata1_103; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2290 = way1_hit ? _GEN_1905 : recent_wdata1_104; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2291 = way1_hit ? _GEN_1906 : recent_wdata1_105; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2292 = way1_hit ? _GEN_1907 : recent_wdata1_106; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2293 = way1_hit ? _GEN_1908 : recent_wdata1_107; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2294 = way1_hit ? _GEN_1909 : recent_wdata1_108; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2295 = way1_hit ? _GEN_1910 : recent_wdata1_109; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2296 = way1_hit ? _GEN_1911 : recent_wdata1_110; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2297 = way1_hit ? _GEN_1912 : recent_wdata1_111; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2298 = way1_hit ? _GEN_1913 : recent_wdata1_112; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2299 = way1_hit ? _GEN_1914 : recent_wdata1_113; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2300 = way1_hit ? _GEN_1915 : recent_wdata1_114; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2301 = way1_hit ? _GEN_1916 : recent_wdata1_115; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2302 = way1_hit ? _GEN_1917 : recent_wdata1_116; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2303 = way1_hit ? _GEN_1918 : recent_wdata1_117; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2304 = way1_hit ? _GEN_1919 : recent_wdata1_118; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2305 = way1_hit ? _GEN_1920 : recent_wdata1_119; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2306 = way1_hit ? _GEN_1921 : recent_wdata1_120; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2307 = way1_hit ? _GEN_1922 : recent_wdata1_121; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2308 = way1_hit ? _GEN_1923 : recent_wdata1_122; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2309 = way1_hit ? _GEN_1924 : recent_wdata1_123; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2310 = way1_hit ? _GEN_1925 : recent_wdata1_124; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2311 = way1_hit ? _GEN_1926 : recent_wdata1_125; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2312 = way1_hit ? _GEN_1927 : recent_wdata1_126; // @[d_cache.scala 115:33 21:32]
  wire [63:0] _GEN_2313 = way1_hit ? _GEN_1928 : recent_wdata1_127; // @[d_cache.scala 115:33 21:32]
  wire  _GEN_2314 = way1_hit ? _GEN_1929 : dirty_1_0; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2315 = way1_hit ? _GEN_1930 : dirty_1_1; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2316 = way1_hit ? _GEN_1931 : dirty_1_2; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2317 = way1_hit ? _GEN_1932 : dirty_1_3; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2318 = way1_hit ? _GEN_1933 : dirty_1_4; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2319 = way1_hit ? _GEN_1934 : dirty_1_5; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2320 = way1_hit ? _GEN_1935 : dirty_1_6; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2321 = way1_hit ? _GEN_1936 : dirty_1_7; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2322 = way1_hit ? _GEN_1937 : dirty_1_8; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2323 = way1_hit ? _GEN_1938 : dirty_1_9; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2324 = way1_hit ? _GEN_1939 : dirty_1_10; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2325 = way1_hit ? _GEN_1940 : dirty_1_11; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2326 = way1_hit ? _GEN_1941 : dirty_1_12; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2327 = way1_hit ? _GEN_1942 : dirty_1_13; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2328 = way1_hit ? _GEN_1943 : dirty_1_14; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2329 = way1_hit ? _GEN_1944 : dirty_1_15; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2330 = way1_hit ? _GEN_1945 : dirty_1_16; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2331 = way1_hit ? _GEN_1946 : dirty_1_17; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2332 = way1_hit ? _GEN_1947 : dirty_1_18; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2333 = way1_hit ? _GEN_1948 : dirty_1_19; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2334 = way1_hit ? _GEN_1949 : dirty_1_20; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2335 = way1_hit ? _GEN_1950 : dirty_1_21; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2336 = way1_hit ? _GEN_1951 : dirty_1_22; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2337 = way1_hit ? _GEN_1952 : dirty_1_23; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2338 = way1_hit ? _GEN_1953 : dirty_1_24; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2339 = way1_hit ? _GEN_1954 : dirty_1_25; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2340 = way1_hit ? _GEN_1955 : dirty_1_26; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2341 = way1_hit ? _GEN_1956 : dirty_1_27; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2342 = way1_hit ? _GEN_1957 : dirty_1_28; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2343 = way1_hit ? _GEN_1958 : dirty_1_29; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2344 = way1_hit ? _GEN_1959 : dirty_1_30; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2345 = way1_hit ? _GEN_1960 : dirty_1_31; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2346 = way1_hit ? _GEN_1961 : dirty_1_32; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2347 = way1_hit ? _GEN_1962 : dirty_1_33; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2348 = way1_hit ? _GEN_1963 : dirty_1_34; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2349 = way1_hit ? _GEN_1964 : dirty_1_35; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2350 = way1_hit ? _GEN_1965 : dirty_1_36; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2351 = way1_hit ? _GEN_1966 : dirty_1_37; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2352 = way1_hit ? _GEN_1967 : dirty_1_38; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2353 = way1_hit ? _GEN_1968 : dirty_1_39; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2354 = way1_hit ? _GEN_1969 : dirty_1_40; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2355 = way1_hit ? _GEN_1970 : dirty_1_41; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2356 = way1_hit ? _GEN_1971 : dirty_1_42; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2357 = way1_hit ? _GEN_1972 : dirty_1_43; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2358 = way1_hit ? _GEN_1973 : dirty_1_44; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2359 = way1_hit ? _GEN_1974 : dirty_1_45; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2360 = way1_hit ? _GEN_1975 : dirty_1_46; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2361 = way1_hit ? _GEN_1976 : dirty_1_47; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2362 = way1_hit ? _GEN_1977 : dirty_1_48; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2363 = way1_hit ? _GEN_1978 : dirty_1_49; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2364 = way1_hit ? _GEN_1979 : dirty_1_50; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2365 = way1_hit ? _GEN_1980 : dirty_1_51; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2366 = way1_hit ? _GEN_1981 : dirty_1_52; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2367 = way1_hit ? _GEN_1982 : dirty_1_53; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2368 = way1_hit ? _GEN_1983 : dirty_1_54; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2369 = way1_hit ? _GEN_1984 : dirty_1_55; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2370 = way1_hit ? _GEN_1985 : dirty_1_56; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2371 = way1_hit ? _GEN_1986 : dirty_1_57; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2372 = way1_hit ? _GEN_1987 : dirty_1_58; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2373 = way1_hit ? _GEN_1988 : dirty_1_59; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2374 = way1_hit ? _GEN_1989 : dirty_1_60; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2375 = way1_hit ? _GEN_1990 : dirty_1_61; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2376 = way1_hit ? _GEN_1991 : dirty_1_62; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2377 = way1_hit ? _GEN_1992 : dirty_1_63; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2378 = way1_hit ? _GEN_1993 : dirty_1_64; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2379 = way1_hit ? _GEN_1994 : dirty_1_65; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2380 = way1_hit ? _GEN_1995 : dirty_1_66; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2381 = way1_hit ? _GEN_1996 : dirty_1_67; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2382 = way1_hit ? _GEN_1997 : dirty_1_68; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2383 = way1_hit ? _GEN_1998 : dirty_1_69; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2384 = way1_hit ? _GEN_1999 : dirty_1_70; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2385 = way1_hit ? _GEN_2000 : dirty_1_71; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2386 = way1_hit ? _GEN_2001 : dirty_1_72; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2387 = way1_hit ? _GEN_2002 : dirty_1_73; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2388 = way1_hit ? _GEN_2003 : dirty_1_74; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2389 = way1_hit ? _GEN_2004 : dirty_1_75; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2390 = way1_hit ? _GEN_2005 : dirty_1_76; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2391 = way1_hit ? _GEN_2006 : dirty_1_77; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2392 = way1_hit ? _GEN_2007 : dirty_1_78; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2393 = way1_hit ? _GEN_2008 : dirty_1_79; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2394 = way1_hit ? _GEN_2009 : dirty_1_80; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2395 = way1_hit ? _GEN_2010 : dirty_1_81; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2396 = way1_hit ? _GEN_2011 : dirty_1_82; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2397 = way1_hit ? _GEN_2012 : dirty_1_83; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2398 = way1_hit ? _GEN_2013 : dirty_1_84; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2399 = way1_hit ? _GEN_2014 : dirty_1_85; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2400 = way1_hit ? _GEN_2015 : dirty_1_86; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2401 = way1_hit ? _GEN_2016 : dirty_1_87; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2402 = way1_hit ? _GEN_2017 : dirty_1_88; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2403 = way1_hit ? _GEN_2018 : dirty_1_89; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2404 = way1_hit ? _GEN_2019 : dirty_1_90; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2405 = way1_hit ? _GEN_2020 : dirty_1_91; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2406 = way1_hit ? _GEN_2021 : dirty_1_92; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2407 = way1_hit ? _GEN_2022 : dirty_1_93; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2408 = way1_hit ? _GEN_2023 : dirty_1_94; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2409 = way1_hit ? _GEN_2024 : dirty_1_95; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2410 = way1_hit ? _GEN_2025 : dirty_1_96; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2411 = way1_hit ? _GEN_2026 : dirty_1_97; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2412 = way1_hit ? _GEN_2027 : dirty_1_98; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2413 = way1_hit ? _GEN_2028 : dirty_1_99; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2414 = way1_hit ? _GEN_2029 : dirty_1_100; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2415 = way1_hit ? _GEN_2030 : dirty_1_101; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2416 = way1_hit ? _GEN_2031 : dirty_1_102; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2417 = way1_hit ? _GEN_2032 : dirty_1_103; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2418 = way1_hit ? _GEN_2033 : dirty_1_104; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2419 = way1_hit ? _GEN_2034 : dirty_1_105; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2420 = way1_hit ? _GEN_2035 : dirty_1_106; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2421 = way1_hit ? _GEN_2036 : dirty_1_107; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2422 = way1_hit ? _GEN_2037 : dirty_1_108; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2423 = way1_hit ? _GEN_2038 : dirty_1_109; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2424 = way1_hit ? _GEN_2039 : dirty_1_110; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2425 = way1_hit ? _GEN_2040 : dirty_1_111; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2426 = way1_hit ? _GEN_2041 : dirty_1_112; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2427 = way1_hit ? _GEN_2042 : dirty_1_113; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2428 = way1_hit ? _GEN_2043 : dirty_1_114; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2429 = way1_hit ? _GEN_2044 : dirty_1_115; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2430 = way1_hit ? _GEN_2045 : dirty_1_116; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2431 = way1_hit ? _GEN_2046 : dirty_1_117; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2432 = way1_hit ? _GEN_2047 : dirty_1_118; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2433 = way1_hit ? _GEN_2048 : dirty_1_119; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2434 = way1_hit ? _GEN_2049 : dirty_1_120; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2435 = way1_hit ? _GEN_2050 : dirty_1_121; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2436 = way1_hit ? _GEN_2051 : dirty_1_122; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2437 = way1_hit ? _GEN_2052 : dirty_1_123; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2438 = way1_hit ? _GEN_2053 : dirty_1_124; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2439 = way1_hit ? _GEN_2054 : dirty_1_125; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2440 = way1_hit ? _GEN_2055 : dirty_1_126; // @[d_cache.scala 115:33 27:26]
  wire  _GEN_2441 = way1_hit ? _GEN_2056 : dirty_1_127; // @[d_cache.scala 115:33 27:26]
  wire [2:0] _GEN_2442 = way0_hit ? 3'h0 : _GEN_2057; // @[d_cache.scala 107:27 108:23]
  wire [63:0] _GEN_2443 = way0_hit ? _GEN_1161 : ram_0_0; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2444 = way0_hit ? _GEN_1162 : ram_0_1; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2445 = way0_hit ? _GEN_1163 : ram_0_2; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2446 = way0_hit ? _GEN_1164 : ram_0_3; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2447 = way0_hit ? _GEN_1165 : ram_0_4; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2448 = way0_hit ? _GEN_1166 : ram_0_5; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2449 = way0_hit ? _GEN_1167 : ram_0_6; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2450 = way0_hit ? _GEN_1168 : ram_0_7; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2451 = way0_hit ? _GEN_1169 : ram_0_8; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2452 = way0_hit ? _GEN_1170 : ram_0_9; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2453 = way0_hit ? _GEN_1171 : ram_0_10; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2454 = way0_hit ? _GEN_1172 : ram_0_11; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2455 = way0_hit ? _GEN_1173 : ram_0_12; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2456 = way0_hit ? _GEN_1174 : ram_0_13; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2457 = way0_hit ? _GEN_1175 : ram_0_14; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2458 = way0_hit ? _GEN_1176 : ram_0_15; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2459 = way0_hit ? _GEN_1177 : ram_0_16; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2460 = way0_hit ? _GEN_1178 : ram_0_17; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2461 = way0_hit ? _GEN_1179 : ram_0_18; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2462 = way0_hit ? _GEN_1180 : ram_0_19; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2463 = way0_hit ? _GEN_1181 : ram_0_20; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2464 = way0_hit ? _GEN_1182 : ram_0_21; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2465 = way0_hit ? _GEN_1183 : ram_0_22; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2466 = way0_hit ? _GEN_1184 : ram_0_23; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2467 = way0_hit ? _GEN_1185 : ram_0_24; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2468 = way0_hit ? _GEN_1186 : ram_0_25; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2469 = way0_hit ? _GEN_1187 : ram_0_26; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2470 = way0_hit ? _GEN_1188 : ram_0_27; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2471 = way0_hit ? _GEN_1189 : ram_0_28; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2472 = way0_hit ? _GEN_1190 : ram_0_29; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2473 = way0_hit ? _GEN_1191 : ram_0_30; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2474 = way0_hit ? _GEN_1192 : ram_0_31; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2475 = way0_hit ? _GEN_1193 : ram_0_32; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2476 = way0_hit ? _GEN_1194 : ram_0_33; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2477 = way0_hit ? _GEN_1195 : ram_0_34; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2478 = way0_hit ? _GEN_1196 : ram_0_35; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2479 = way0_hit ? _GEN_1197 : ram_0_36; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2480 = way0_hit ? _GEN_1198 : ram_0_37; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2481 = way0_hit ? _GEN_1199 : ram_0_38; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2482 = way0_hit ? _GEN_1200 : ram_0_39; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2483 = way0_hit ? _GEN_1201 : ram_0_40; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2484 = way0_hit ? _GEN_1202 : ram_0_41; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2485 = way0_hit ? _GEN_1203 : ram_0_42; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2486 = way0_hit ? _GEN_1204 : ram_0_43; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2487 = way0_hit ? _GEN_1205 : ram_0_44; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2488 = way0_hit ? _GEN_1206 : ram_0_45; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2489 = way0_hit ? _GEN_1207 : ram_0_46; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2490 = way0_hit ? _GEN_1208 : ram_0_47; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2491 = way0_hit ? _GEN_1209 : ram_0_48; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2492 = way0_hit ? _GEN_1210 : ram_0_49; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2493 = way0_hit ? _GEN_1211 : ram_0_50; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2494 = way0_hit ? _GEN_1212 : ram_0_51; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2495 = way0_hit ? _GEN_1213 : ram_0_52; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2496 = way0_hit ? _GEN_1214 : ram_0_53; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2497 = way0_hit ? _GEN_1215 : ram_0_54; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2498 = way0_hit ? _GEN_1216 : ram_0_55; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2499 = way0_hit ? _GEN_1217 : ram_0_56; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2500 = way0_hit ? _GEN_1218 : ram_0_57; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2501 = way0_hit ? _GEN_1219 : ram_0_58; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2502 = way0_hit ? _GEN_1220 : ram_0_59; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2503 = way0_hit ? _GEN_1221 : ram_0_60; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2504 = way0_hit ? _GEN_1222 : ram_0_61; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2505 = way0_hit ? _GEN_1223 : ram_0_62; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2506 = way0_hit ? _GEN_1224 : ram_0_63; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2507 = way0_hit ? _GEN_1225 : ram_0_64; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2508 = way0_hit ? _GEN_1226 : ram_0_65; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2509 = way0_hit ? _GEN_1227 : ram_0_66; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2510 = way0_hit ? _GEN_1228 : ram_0_67; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2511 = way0_hit ? _GEN_1229 : ram_0_68; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2512 = way0_hit ? _GEN_1230 : ram_0_69; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2513 = way0_hit ? _GEN_1231 : ram_0_70; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2514 = way0_hit ? _GEN_1232 : ram_0_71; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2515 = way0_hit ? _GEN_1233 : ram_0_72; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2516 = way0_hit ? _GEN_1234 : ram_0_73; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2517 = way0_hit ? _GEN_1235 : ram_0_74; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2518 = way0_hit ? _GEN_1236 : ram_0_75; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2519 = way0_hit ? _GEN_1237 : ram_0_76; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2520 = way0_hit ? _GEN_1238 : ram_0_77; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2521 = way0_hit ? _GEN_1239 : ram_0_78; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2522 = way0_hit ? _GEN_1240 : ram_0_79; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2523 = way0_hit ? _GEN_1241 : ram_0_80; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2524 = way0_hit ? _GEN_1242 : ram_0_81; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2525 = way0_hit ? _GEN_1243 : ram_0_82; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2526 = way0_hit ? _GEN_1244 : ram_0_83; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2527 = way0_hit ? _GEN_1245 : ram_0_84; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2528 = way0_hit ? _GEN_1246 : ram_0_85; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2529 = way0_hit ? _GEN_1247 : ram_0_86; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2530 = way0_hit ? _GEN_1248 : ram_0_87; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2531 = way0_hit ? _GEN_1249 : ram_0_88; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2532 = way0_hit ? _GEN_1250 : ram_0_89; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2533 = way0_hit ? _GEN_1251 : ram_0_90; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2534 = way0_hit ? _GEN_1252 : ram_0_91; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2535 = way0_hit ? _GEN_1253 : ram_0_92; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2536 = way0_hit ? _GEN_1254 : ram_0_93; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2537 = way0_hit ? _GEN_1255 : ram_0_94; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2538 = way0_hit ? _GEN_1256 : ram_0_95; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2539 = way0_hit ? _GEN_1257 : ram_0_96; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2540 = way0_hit ? _GEN_1258 : ram_0_97; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2541 = way0_hit ? _GEN_1259 : ram_0_98; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2542 = way0_hit ? _GEN_1260 : ram_0_99; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2543 = way0_hit ? _GEN_1261 : ram_0_100; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2544 = way0_hit ? _GEN_1262 : ram_0_101; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2545 = way0_hit ? _GEN_1263 : ram_0_102; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2546 = way0_hit ? _GEN_1264 : ram_0_103; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2547 = way0_hit ? _GEN_1265 : ram_0_104; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2548 = way0_hit ? _GEN_1266 : ram_0_105; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2549 = way0_hit ? _GEN_1267 : ram_0_106; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2550 = way0_hit ? _GEN_1268 : ram_0_107; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2551 = way0_hit ? _GEN_1269 : ram_0_108; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2552 = way0_hit ? _GEN_1270 : ram_0_109; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2553 = way0_hit ? _GEN_1271 : ram_0_110; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2554 = way0_hit ? _GEN_1272 : ram_0_111; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2555 = way0_hit ? _GEN_1273 : ram_0_112; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2556 = way0_hit ? _GEN_1274 : ram_0_113; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2557 = way0_hit ? _GEN_1275 : ram_0_114; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2558 = way0_hit ? _GEN_1276 : ram_0_115; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2559 = way0_hit ? _GEN_1277 : ram_0_116; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2560 = way0_hit ? _GEN_1278 : ram_0_117; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2561 = way0_hit ? _GEN_1279 : ram_0_118; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2562 = way0_hit ? _GEN_1280 : ram_0_119; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2563 = way0_hit ? _GEN_1281 : ram_0_120; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2564 = way0_hit ? _GEN_1282 : ram_0_121; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2565 = way0_hit ? _GEN_1283 : ram_0_122; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2566 = way0_hit ? _GEN_1284 : ram_0_123; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2567 = way0_hit ? _GEN_1285 : ram_0_124; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2568 = way0_hit ? _GEN_1286 : ram_0_125; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2569 = way0_hit ? _GEN_1287 : ram_0_126; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2570 = way0_hit ? _GEN_1288 : ram_0_127; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_2571 = way0_hit ? _GEN_1289 : recent_wdata0_0; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2572 = way0_hit ? _GEN_1290 : recent_wdata0_1; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2573 = way0_hit ? _GEN_1291 : recent_wdata0_2; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2574 = way0_hit ? _GEN_1292 : recent_wdata0_3; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2575 = way0_hit ? _GEN_1293 : recent_wdata0_4; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2576 = way0_hit ? _GEN_1294 : recent_wdata0_5; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2577 = way0_hit ? _GEN_1295 : recent_wdata0_6; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2578 = way0_hit ? _GEN_1296 : recent_wdata0_7; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2579 = way0_hit ? _GEN_1297 : recent_wdata0_8; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2580 = way0_hit ? _GEN_1298 : recent_wdata0_9; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2581 = way0_hit ? _GEN_1299 : recent_wdata0_10; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2582 = way0_hit ? _GEN_1300 : recent_wdata0_11; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2583 = way0_hit ? _GEN_1301 : recent_wdata0_12; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2584 = way0_hit ? _GEN_1302 : recent_wdata0_13; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2585 = way0_hit ? _GEN_1303 : recent_wdata0_14; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2586 = way0_hit ? _GEN_1304 : recent_wdata0_15; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2587 = way0_hit ? _GEN_1305 : recent_wdata0_16; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2588 = way0_hit ? _GEN_1306 : recent_wdata0_17; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2589 = way0_hit ? _GEN_1307 : recent_wdata0_18; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2590 = way0_hit ? _GEN_1308 : recent_wdata0_19; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2591 = way0_hit ? _GEN_1309 : recent_wdata0_20; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2592 = way0_hit ? _GEN_1310 : recent_wdata0_21; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2593 = way0_hit ? _GEN_1311 : recent_wdata0_22; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2594 = way0_hit ? _GEN_1312 : recent_wdata0_23; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2595 = way0_hit ? _GEN_1313 : recent_wdata0_24; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2596 = way0_hit ? _GEN_1314 : recent_wdata0_25; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2597 = way0_hit ? _GEN_1315 : recent_wdata0_26; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2598 = way0_hit ? _GEN_1316 : recent_wdata0_27; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2599 = way0_hit ? _GEN_1317 : recent_wdata0_28; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2600 = way0_hit ? _GEN_1318 : recent_wdata0_29; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2601 = way0_hit ? _GEN_1319 : recent_wdata0_30; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2602 = way0_hit ? _GEN_1320 : recent_wdata0_31; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2603 = way0_hit ? _GEN_1321 : recent_wdata0_32; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2604 = way0_hit ? _GEN_1322 : recent_wdata0_33; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2605 = way0_hit ? _GEN_1323 : recent_wdata0_34; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2606 = way0_hit ? _GEN_1324 : recent_wdata0_35; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2607 = way0_hit ? _GEN_1325 : recent_wdata0_36; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2608 = way0_hit ? _GEN_1326 : recent_wdata0_37; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2609 = way0_hit ? _GEN_1327 : recent_wdata0_38; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2610 = way0_hit ? _GEN_1328 : recent_wdata0_39; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2611 = way0_hit ? _GEN_1329 : recent_wdata0_40; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2612 = way0_hit ? _GEN_1330 : recent_wdata0_41; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2613 = way0_hit ? _GEN_1331 : recent_wdata0_42; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2614 = way0_hit ? _GEN_1332 : recent_wdata0_43; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2615 = way0_hit ? _GEN_1333 : recent_wdata0_44; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2616 = way0_hit ? _GEN_1334 : recent_wdata0_45; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2617 = way0_hit ? _GEN_1335 : recent_wdata0_46; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2618 = way0_hit ? _GEN_1336 : recent_wdata0_47; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2619 = way0_hit ? _GEN_1337 : recent_wdata0_48; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2620 = way0_hit ? _GEN_1338 : recent_wdata0_49; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2621 = way0_hit ? _GEN_1339 : recent_wdata0_50; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2622 = way0_hit ? _GEN_1340 : recent_wdata0_51; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2623 = way0_hit ? _GEN_1341 : recent_wdata0_52; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2624 = way0_hit ? _GEN_1342 : recent_wdata0_53; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2625 = way0_hit ? _GEN_1343 : recent_wdata0_54; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2626 = way0_hit ? _GEN_1344 : recent_wdata0_55; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2627 = way0_hit ? _GEN_1345 : recent_wdata0_56; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2628 = way0_hit ? _GEN_1346 : recent_wdata0_57; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2629 = way0_hit ? _GEN_1347 : recent_wdata0_58; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2630 = way0_hit ? _GEN_1348 : recent_wdata0_59; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2631 = way0_hit ? _GEN_1349 : recent_wdata0_60; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2632 = way0_hit ? _GEN_1350 : recent_wdata0_61; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2633 = way0_hit ? _GEN_1351 : recent_wdata0_62; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2634 = way0_hit ? _GEN_1352 : recent_wdata0_63; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2635 = way0_hit ? _GEN_1353 : recent_wdata0_64; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2636 = way0_hit ? _GEN_1354 : recent_wdata0_65; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2637 = way0_hit ? _GEN_1355 : recent_wdata0_66; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2638 = way0_hit ? _GEN_1356 : recent_wdata0_67; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2639 = way0_hit ? _GEN_1357 : recent_wdata0_68; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2640 = way0_hit ? _GEN_1358 : recent_wdata0_69; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2641 = way0_hit ? _GEN_1359 : recent_wdata0_70; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2642 = way0_hit ? _GEN_1360 : recent_wdata0_71; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2643 = way0_hit ? _GEN_1361 : recent_wdata0_72; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2644 = way0_hit ? _GEN_1362 : recent_wdata0_73; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2645 = way0_hit ? _GEN_1363 : recent_wdata0_74; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2646 = way0_hit ? _GEN_1364 : recent_wdata0_75; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2647 = way0_hit ? _GEN_1365 : recent_wdata0_76; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2648 = way0_hit ? _GEN_1366 : recent_wdata0_77; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2649 = way0_hit ? _GEN_1367 : recent_wdata0_78; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2650 = way0_hit ? _GEN_1368 : recent_wdata0_79; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2651 = way0_hit ? _GEN_1369 : recent_wdata0_80; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2652 = way0_hit ? _GEN_1370 : recent_wdata0_81; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2653 = way0_hit ? _GEN_1371 : recent_wdata0_82; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2654 = way0_hit ? _GEN_1372 : recent_wdata0_83; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2655 = way0_hit ? _GEN_1373 : recent_wdata0_84; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2656 = way0_hit ? _GEN_1374 : recent_wdata0_85; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2657 = way0_hit ? _GEN_1375 : recent_wdata0_86; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2658 = way0_hit ? _GEN_1376 : recent_wdata0_87; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2659 = way0_hit ? _GEN_1377 : recent_wdata0_88; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2660 = way0_hit ? _GEN_1378 : recent_wdata0_89; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2661 = way0_hit ? _GEN_1379 : recent_wdata0_90; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2662 = way0_hit ? _GEN_1380 : recent_wdata0_91; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2663 = way0_hit ? _GEN_1381 : recent_wdata0_92; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2664 = way0_hit ? _GEN_1382 : recent_wdata0_93; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2665 = way0_hit ? _GEN_1383 : recent_wdata0_94; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2666 = way0_hit ? _GEN_1384 : recent_wdata0_95; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2667 = way0_hit ? _GEN_1385 : recent_wdata0_96; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2668 = way0_hit ? _GEN_1386 : recent_wdata0_97; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2669 = way0_hit ? _GEN_1387 : recent_wdata0_98; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2670 = way0_hit ? _GEN_1388 : recent_wdata0_99; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2671 = way0_hit ? _GEN_1389 : recent_wdata0_100; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2672 = way0_hit ? _GEN_1390 : recent_wdata0_101; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2673 = way0_hit ? _GEN_1391 : recent_wdata0_102; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2674 = way0_hit ? _GEN_1392 : recent_wdata0_103; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2675 = way0_hit ? _GEN_1393 : recent_wdata0_104; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2676 = way0_hit ? _GEN_1394 : recent_wdata0_105; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2677 = way0_hit ? _GEN_1395 : recent_wdata0_106; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2678 = way0_hit ? _GEN_1396 : recent_wdata0_107; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2679 = way0_hit ? _GEN_1397 : recent_wdata0_108; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2680 = way0_hit ? _GEN_1398 : recent_wdata0_109; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2681 = way0_hit ? _GEN_1399 : recent_wdata0_110; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2682 = way0_hit ? _GEN_1400 : recent_wdata0_111; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2683 = way0_hit ? _GEN_1401 : recent_wdata0_112; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2684 = way0_hit ? _GEN_1402 : recent_wdata0_113; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2685 = way0_hit ? _GEN_1403 : recent_wdata0_114; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2686 = way0_hit ? _GEN_1404 : recent_wdata0_115; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2687 = way0_hit ? _GEN_1405 : recent_wdata0_116; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2688 = way0_hit ? _GEN_1406 : recent_wdata0_117; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2689 = way0_hit ? _GEN_1407 : recent_wdata0_118; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2690 = way0_hit ? _GEN_1408 : recent_wdata0_119; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2691 = way0_hit ? _GEN_1409 : recent_wdata0_120; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2692 = way0_hit ? _GEN_1410 : recent_wdata0_121; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2693 = way0_hit ? _GEN_1411 : recent_wdata0_122; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2694 = way0_hit ? _GEN_1412 : recent_wdata0_123; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2695 = way0_hit ? _GEN_1413 : recent_wdata0_124; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2696 = way0_hit ? _GEN_1414 : recent_wdata0_125; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2697 = way0_hit ? _GEN_1415 : recent_wdata0_126; // @[d_cache.scala 107:27 20:32]
  wire [63:0] _GEN_2698 = way0_hit ? _GEN_1416 : recent_wdata0_127; // @[d_cache.scala 107:27 20:32]
  wire  _GEN_2699 = way0_hit ? _GEN_1417 : dirty_0_0; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2700 = way0_hit ? _GEN_1418 : dirty_0_1; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2701 = way0_hit ? _GEN_1419 : dirty_0_2; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2702 = way0_hit ? _GEN_1420 : dirty_0_3; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2703 = way0_hit ? _GEN_1421 : dirty_0_4; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2704 = way0_hit ? _GEN_1422 : dirty_0_5; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2705 = way0_hit ? _GEN_1423 : dirty_0_6; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2706 = way0_hit ? _GEN_1424 : dirty_0_7; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2707 = way0_hit ? _GEN_1425 : dirty_0_8; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2708 = way0_hit ? _GEN_1426 : dirty_0_9; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2709 = way0_hit ? _GEN_1427 : dirty_0_10; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2710 = way0_hit ? _GEN_1428 : dirty_0_11; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2711 = way0_hit ? _GEN_1429 : dirty_0_12; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2712 = way0_hit ? _GEN_1430 : dirty_0_13; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2713 = way0_hit ? _GEN_1431 : dirty_0_14; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2714 = way0_hit ? _GEN_1432 : dirty_0_15; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2715 = way0_hit ? _GEN_1433 : dirty_0_16; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2716 = way0_hit ? _GEN_1434 : dirty_0_17; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2717 = way0_hit ? _GEN_1435 : dirty_0_18; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2718 = way0_hit ? _GEN_1436 : dirty_0_19; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2719 = way0_hit ? _GEN_1437 : dirty_0_20; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2720 = way0_hit ? _GEN_1438 : dirty_0_21; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2721 = way0_hit ? _GEN_1439 : dirty_0_22; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2722 = way0_hit ? _GEN_1440 : dirty_0_23; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2723 = way0_hit ? _GEN_1441 : dirty_0_24; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2724 = way0_hit ? _GEN_1442 : dirty_0_25; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2725 = way0_hit ? _GEN_1443 : dirty_0_26; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2726 = way0_hit ? _GEN_1444 : dirty_0_27; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2727 = way0_hit ? _GEN_1445 : dirty_0_28; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2728 = way0_hit ? _GEN_1446 : dirty_0_29; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2729 = way0_hit ? _GEN_1447 : dirty_0_30; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2730 = way0_hit ? _GEN_1448 : dirty_0_31; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2731 = way0_hit ? _GEN_1449 : dirty_0_32; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2732 = way0_hit ? _GEN_1450 : dirty_0_33; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2733 = way0_hit ? _GEN_1451 : dirty_0_34; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2734 = way0_hit ? _GEN_1452 : dirty_0_35; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2735 = way0_hit ? _GEN_1453 : dirty_0_36; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2736 = way0_hit ? _GEN_1454 : dirty_0_37; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2737 = way0_hit ? _GEN_1455 : dirty_0_38; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2738 = way0_hit ? _GEN_1456 : dirty_0_39; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2739 = way0_hit ? _GEN_1457 : dirty_0_40; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2740 = way0_hit ? _GEN_1458 : dirty_0_41; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2741 = way0_hit ? _GEN_1459 : dirty_0_42; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2742 = way0_hit ? _GEN_1460 : dirty_0_43; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2743 = way0_hit ? _GEN_1461 : dirty_0_44; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2744 = way0_hit ? _GEN_1462 : dirty_0_45; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2745 = way0_hit ? _GEN_1463 : dirty_0_46; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2746 = way0_hit ? _GEN_1464 : dirty_0_47; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2747 = way0_hit ? _GEN_1465 : dirty_0_48; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2748 = way0_hit ? _GEN_1466 : dirty_0_49; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2749 = way0_hit ? _GEN_1467 : dirty_0_50; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2750 = way0_hit ? _GEN_1468 : dirty_0_51; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2751 = way0_hit ? _GEN_1469 : dirty_0_52; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2752 = way0_hit ? _GEN_1470 : dirty_0_53; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2753 = way0_hit ? _GEN_1471 : dirty_0_54; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2754 = way0_hit ? _GEN_1472 : dirty_0_55; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2755 = way0_hit ? _GEN_1473 : dirty_0_56; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2756 = way0_hit ? _GEN_1474 : dirty_0_57; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2757 = way0_hit ? _GEN_1475 : dirty_0_58; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2758 = way0_hit ? _GEN_1476 : dirty_0_59; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2759 = way0_hit ? _GEN_1477 : dirty_0_60; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2760 = way0_hit ? _GEN_1478 : dirty_0_61; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2761 = way0_hit ? _GEN_1479 : dirty_0_62; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2762 = way0_hit ? _GEN_1480 : dirty_0_63; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2763 = way0_hit ? _GEN_1481 : dirty_0_64; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2764 = way0_hit ? _GEN_1482 : dirty_0_65; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2765 = way0_hit ? _GEN_1483 : dirty_0_66; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2766 = way0_hit ? _GEN_1484 : dirty_0_67; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2767 = way0_hit ? _GEN_1485 : dirty_0_68; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2768 = way0_hit ? _GEN_1486 : dirty_0_69; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2769 = way0_hit ? _GEN_1487 : dirty_0_70; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2770 = way0_hit ? _GEN_1488 : dirty_0_71; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2771 = way0_hit ? _GEN_1489 : dirty_0_72; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2772 = way0_hit ? _GEN_1490 : dirty_0_73; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2773 = way0_hit ? _GEN_1491 : dirty_0_74; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2774 = way0_hit ? _GEN_1492 : dirty_0_75; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2775 = way0_hit ? _GEN_1493 : dirty_0_76; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2776 = way0_hit ? _GEN_1494 : dirty_0_77; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2777 = way0_hit ? _GEN_1495 : dirty_0_78; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2778 = way0_hit ? _GEN_1496 : dirty_0_79; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2779 = way0_hit ? _GEN_1497 : dirty_0_80; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2780 = way0_hit ? _GEN_1498 : dirty_0_81; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2781 = way0_hit ? _GEN_1499 : dirty_0_82; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2782 = way0_hit ? _GEN_1500 : dirty_0_83; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2783 = way0_hit ? _GEN_1501 : dirty_0_84; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2784 = way0_hit ? _GEN_1502 : dirty_0_85; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2785 = way0_hit ? _GEN_1503 : dirty_0_86; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2786 = way0_hit ? _GEN_1504 : dirty_0_87; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2787 = way0_hit ? _GEN_1505 : dirty_0_88; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2788 = way0_hit ? _GEN_1506 : dirty_0_89; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2789 = way0_hit ? _GEN_1507 : dirty_0_90; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2790 = way0_hit ? _GEN_1508 : dirty_0_91; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2791 = way0_hit ? _GEN_1509 : dirty_0_92; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2792 = way0_hit ? _GEN_1510 : dirty_0_93; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2793 = way0_hit ? _GEN_1511 : dirty_0_94; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2794 = way0_hit ? _GEN_1512 : dirty_0_95; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2795 = way0_hit ? _GEN_1513 : dirty_0_96; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2796 = way0_hit ? _GEN_1514 : dirty_0_97; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2797 = way0_hit ? _GEN_1515 : dirty_0_98; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2798 = way0_hit ? _GEN_1516 : dirty_0_99; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2799 = way0_hit ? _GEN_1517 : dirty_0_100; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2800 = way0_hit ? _GEN_1518 : dirty_0_101; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2801 = way0_hit ? _GEN_1519 : dirty_0_102; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2802 = way0_hit ? _GEN_1520 : dirty_0_103; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2803 = way0_hit ? _GEN_1521 : dirty_0_104; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2804 = way0_hit ? _GEN_1522 : dirty_0_105; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2805 = way0_hit ? _GEN_1523 : dirty_0_106; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2806 = way0_hit ? _GEN_1524 : dirty_0_107; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2807 = way0_hit ? _GEN_1525 : dirty_0_108; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2808 = way0_hit ? _GEN_1526 : dirty_0_109; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2809 = way0_hit ? _GEN_1527 : dirty_0_110; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2810 = way0_hit ? _GEN_1528 : dirty_0_111; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2811 = way0_hit ? _GEN_1529 : dirty_0_112; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2812 = way0_hit ? _GEN_1530 : dirty_0_113; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2813 = way0_hit ? _GEN_1531 : dirty_0_114; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2814 = way0_hit ? _GEN_1532 : dirty_0_115; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2815 = way0_hit ? _GEN_1533 : dirty_0_116; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2816 = way0_hit ? _GEN_1534 : dirty_0_117; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2817 = way0_hit ? _GEN_1535 : dirty_0_118; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2818 = way0_hit ? _GEN_1536 : dirty_0_119; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2819 = way0_hit ? _GEN_1537 : dirty_0_120; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2820 = way0_hit ? _GEN_1538 : dirty_0_121; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2821 = way0_hit ? _GEN_1539 : dirty_0_122; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2822 = way0_hit ? _GEN_1540 : dirty_0_123; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2823 = way0_hit ? _GEN_1541 : dirty_0_124; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2824 = way0_hit ? _GEN_1542 : dirty_0_125; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2825 = way0_hit ? _GEN_1543 : dirty_0_126; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_2826 = way0_hit ? _GEN_1544 : dirty_0_127; // @[d_cache.scala 107:27 26:26]
  wire [63:0] _GEN_2827 = way0_hit ? ram_1_0 : _GEN_2058; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2828 = way0_hit ? ram_1_1 : _GEN_2059; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2829 = way0_hit ? ram_1_2 : _GEN_2060; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2830 = way0_hit ? ram_1_3 : _GEN_2061; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2831 = way0_hit ? ram_1_4 : _GEN_2062; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2832 = way0_hit ? ram_1_5 : _GEN_2063; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2833 = way0_hit ? ram_1_6 : _GEN_2064; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2834 = way0_hit ? ram_1_7 : _GEN_2065; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2835 = way0_hit ? ram_1_8 : _GEN_2066; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2836 = way0_hit ? ram_1_9 : _GEN_2067; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2837 = way0_hit ? ram_1_10 : _GEN_2068; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2838 = way0_hit ? ram_1_11 : _GEN_2069; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2839 = way0_hit ? ram_1_12 : _GEN_2070; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2840 = way0_hit ? ram_1_13 : _GEN_2071; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2841 = way0_hit ? ram_1_14 : _GEN_2072; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2842 = way0_hit ? ram_1_15 : _GEN_2073; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2843 = way0_hit ? ram_1_16 : _GEN_2074; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2844 = way0_hit ? ram_1_17 : _GEN_2075; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2845 = way0_hit ? ram_1_18 : _GEN_2076; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2846 = way0_hit ? ram_1_19 : _GEN_2077; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2847 = way0_hit ? ram_1_20 : _GEN_2078; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2848 = way0_hit ? ram_1_21 : _GEN_2079; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2849 = way0_hit ? ram_1_22 : _GEN_2080; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2850 = way0_hit ? ram_1_23 : _GEN_2081; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2851 = way0_hit ? ram_1_24 : _GEN_2082; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2852 = way0_hit ? ram_1_25 : _GEN_2083; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2853 = way0_hit ? ram_1_26 : _GEN_2084; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2854 = way0_hit ? ram_1_27 : _GEN_2085; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2855 = way0_hit ? ram_1_28 : _GEN_2086; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2856 = way0_hit ? ram_1_29 : _GEN_2087; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2857 = way0_hit ? ram_1_30 : _GEN_2088; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2858 = way0_hit ? ram_1_31 : _GEN_2089; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2859 = way0_hit ? ram_1_32 : _GEN_2090; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2860 = way0_hit ? ram_1_33 : _GEN_2091; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2861 = way0_hit ? ram_1_34 : _GEN_2092; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2862 = way0_hit ? ram_1_35 : _GEN_2093; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2863 = way0_hit ? ram_1_36 : _GEN_2094; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2864 = way0_hit ? ram_1_37 : _GEN_2095; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2865 = way0_hit ? ram_1_38 : _GEN_2096; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2866 = way0_hit ? ram_1_39 : _GEN_2097; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2867 = way0_hit ? ram_1_40 : _GEN_2098; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2868 = way0_hit ? ram_1_41 : _GEN_2099; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2869 = way0_hit ? ram_1_42 : _GEN_2100; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2870 = way0_hit ? ram_1_43 : _GEN_2101; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2871 = way0_hit ? ram_1_44 : _GEN_2102; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2872 = way0_hit ? ram_1_45 : _GEN_2103; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2873 = way0_hit ? ram_1_46 : _GEN_2104; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2874 = way0_hit ? ram_1_47 : _GEN_2105; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2875 = way0_hit ? ram_1_48 : _GEN_2106; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2876 = way0_hit ? ram_1_49 : _GEN_2107; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2877 = way0_hit ? ram_1_50 : _GEN_2108; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2878 = way0_hit ? ram_1_51 : _GEN_2109; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2879 = way0_hit ? ram_1_52 : _GEN_2110; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2880 = way0_hit ? ram_1_53 : _GEN_2111; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2881 = way0_hit ? ram_1_54 : _GEN_2112; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2882 = way0_hit ? ram_1_55 : _GEN_2113; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2883 = way0_hit ? ram_1_56 : _GEN_2114; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2884 = way0_hit ? ram_1_57 : _GEN_2115; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2885 = way0_hit ? ram_1_58 : _GEN_2116; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2886 = way0_hit ? ram_1_59 : _GEN_2117; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2887 = way0_hit ? ram_1_60 : _GEN_2118; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2888 = way0_hit ? ram_1_61 : _GEN_2119; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2889 = way0_hit ? ram_1_62 : _GEN_2120; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2890 = way0_hit ? ram_1_63 : _GEN_2121; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2891 = way0_hit ? ram_1_64 : _GEN_2122; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2892 = way0_hit ? ram_1_65 : _GEN_2123; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2893 = way0_hit ? ram_1_66 : _GEN_2124; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2894 = way0_hit ? ram_1_67 : _GEN_2125; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2895 = way0_hit ? ram_1_68 : _GEN_2126; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2896 = way0_hit ? ram_1_69 : _GEN_2127; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2897 = way0_hit ? ram_1_70 : _GEN_2128; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2898 = way0_hit ? ram_1_71 : _GEN_2129; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2899 = way0_hit ? ram_1_72 : _GEN_2130; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2900 = way0_hit ? ram_1_73 : _GEN_2131; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2901 = way0_hit ? ram_1_74 : _GEN_2132; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2902 = way0_hit ? ram_1_75 : _GEN_2133; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2903 = way0_hit ? ram_1_76 : _GEN_2134; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2904 = way0_hit ? ram_1_77 : _GEN_2135; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2905 = way0_hit ? ram_1_78 : _GEN_2136; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2906 = way0_hit ? ram_1_79 : _GEN_2137; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2907 = way0_hit ? ram_1_80 : _GEN_2138; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2908 = way0_hit ? ram_1_81 : _GEN_2139; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2909 = way0_hit ? ram_1_82 : _GEN_2140; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2910 = way0_hit ? ram_1_83 : _GEN_2141; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2911 = way0_hit ? ram_1_84 : _GEN_2142; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2912 = way0_hit ? ram_1_85 : _GEN_2143; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2913 = way0_hit ? ram_1_86 : _GEN_2144; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2914 = way0_hit ? ram_1_87 : _GEN_2145; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2915 = way0_hit ? ram_1_88 : _GEN_2146; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2916 = way0_hit ? ram_1_89 : _GEN_2147; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2917 = way0_hit ? ram_1_90 : _GEN_2148; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2918 = way0_hit ? ram_1_91 : _GEN_2149; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2919 = way0_hit ? ram_1_92 : _GEN_2150; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2920 = way0_hit ? ram_1_93 : _GEN_2151; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2921 = way0_hit ? ram_1_94 : _GEN_2152; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2922 = way0_hit ? ram_1_95 : _GEN_2153; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2923 = way0_hit ? ram_1_96 : _GEN_2154; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2924 = way0_hit ? ram_1_97 : _GEN_2155; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2925 = way0_hit ? ram_1_98 : _GEN_2156; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2926 = way0_hit ? ram_1_99 : _GEN_2157; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2927 = way0_hit ? ram_1_100 : _GEN_2158; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2928 = way0_hit ? ram_1_101 : _GEN_2159; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2929 = way0_hit ? ram_1_102 : _GEN_2160; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2930 = way0_hit ? ram_1_103 : _GEN_2161; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2931 = way0_hit ? ram_1_104 : _GEN_2162; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2932 = way0_hit ? ram_1_105 : _GEN_2163; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2933 = way0_hit ? ram_1_106 : _GEN_2164; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2934 = way0_hit ? ram_1_107 : _GEN_2165; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2935 = way0_hit ? ram_1_108 : _GEN_2166; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2936 = way0_hit ? ram_1_109 : _GEN_2167; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2937 = way0_hit ? ram_1_110 : _GEN_2168; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2938 = way0_hit ? ram_1_111 : _GEN_2169; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2939 = way0_hit ? ram_1_112 : _GEN_2170; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2940 = way0_hit ? ram_1_113 : _GEN_2171; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2941 = way0_hit ? ram_1_114 : _GEN_2172; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2942 = way0_hit ? ram_1_115 : _GEN_2173; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2943 = way0_hit ? ram_1_116 : _GEN_2174; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2944 = way0_hit ? ram_1_117 : _GEN_2175; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2945 = way0_hit ? ram_1_118 : _GEN_2176; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2946 = way0_hit ? ram_1_119 : _GEN_2177; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2947 = way0_hit ? ram_1_120 : _GEN_2178; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2948 = way0_hit ? ram_1_121 : _GEN_2179; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2949 = way0_hit ? ram_1_122 : _GEN_2180; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2950 = way0_hit ? ram_1_123 : _GEN_2181; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2951 = way0_hit ? ram_1_124 : _GEN_2182; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2952 = way0_hit ? ram_1_125 : _GEN_2183; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2953 = way0_hit ? ram_1_126 : _GEN_2184; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2954 = way0_hit ? ram_1_127 : _GEN_2185; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_2955 = way0_hit ? recent_wdata1_0 : _GEN_2186; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2956 = way0_hit ? recent_wdata1_1 : _GEN_2187; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2957 = way0_hit ? recent_wdata1_2 : _GEN_2188; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2958 = way0_hit ? recent_wdata1_3 : _GEN_2189; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2959 = way0_hit ? recent_wdata1_4 : _GEN_2190; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2960 = way0_hit ? recent_wdata1_5 : _GEN_2191; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2961 = way0_hit ? recent_wdata1_6 : _GEN_2192; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2962 = way0_hit ? recent_wdata1_7 : _GEN_2193; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2963 = way0_hit ? recent_wdata1_8 : _GEN_2194; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2964 = way0_hit ? recent_wdata1_9 : _GEN_2195; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2965 = way0_hit ? recent_wdata1_10 : _GEN_2196; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2966 = way0_hit ? recent_wdata1_11 : _GEN_2197; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2967 = way0_hit ? recent_wdata1_12 : _GEN_2198; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2968 = way0_hit ? recent_wdata1_13 : _GEN_2199; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2969 = way0_hit ? recent_wdata1_14 : _GEN_2200; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2970 = way0_hit ? recent_wdata1_15 : _GEN_2201; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2971 = way0_hit ? recent_wdata1_16 : _GEN_2202; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2972 = way0_hit ? recent_wdata1_17 : _GEN_2203; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2973 = way0_hit ? recent_wdata1_18 : _GEN_2204; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2974 = way0_hit ? recent_wdata1_19 : _GEN_2205; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2975 = way0_hit ? recent_wdata1_20 : _GEN_2206; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2976 = way0_hit ? recent_wdata1_21 : _GEN_2207; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2977 = way0_hit ? recent_wdata1_22 : _GEN_2208; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2978 = way0_hit ? recent_wdata1_23 : _GEN_2209; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2979 = way0_hit ? recent_wdata1_24 : _GEN_2210; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2980 = way0_hit ? recent_wdata1_25 : _GEN_2211; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2981 = way0_hit ? recent_wdata1_26 : _GEN_2212; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2982 = way0_hit ? recent_wdata1_27 : _GEN_2213; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2983 = way0_hit ? recent_wdata1_28 : _GEN_2214; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2984 = way0_hit ? recent_wdata1_29 : _GEN_2215; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2985 = way0_hit ? recent_wdata1_30 : _GEN_2216; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2986 = way0_hit ? recent_wdata1_31 : _GEN_2217; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2987 = way0_hit ? recent_wdata1_32 : _GEN_2218; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2988 = way0_hit ? recent_wdata1_33 : _GEN_2219; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2989 = way0_hit ? recent_wdata1_34 : _GEN_2220; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2990 = way0_hit ? recent_wdata1_35 : _GEN_2221; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2991 = way0_hit ? recent_wdata1_36 : _GEN_2222; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2992 = way0_hit ? recent_wdata1_37 : _GEN_2223; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2993 = way0_hit ? recent_wdata1_38 : _GEN_2224; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2994 = way0_hit ? recent_wdata1_39 : _GEN_2225; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2995 = way0_hit ? recent_wdata1_40 : _GEN_2226; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2996 = way0_hit ? recent_wdata1_41 : _GEN_2227; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2997 = way0_hit ? recent_wdata1_42 : _GEN_2228; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2998 = way0_hit ? recent_wdata1_43 : _GEN_2229; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_2999 = way0_hit ? recent_wdata1_44 : _GEN_2230; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3000 = way0_hit ? recent_wdata1_45 : _GEN_2231; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3001 = way0_hit ? recent_wdata1_46 : _GEN_2232; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3002 = way0_hit ? recent_wdata1_47 : _GEN_2233; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3003 = way0_hit ? recent_wdata1_48 : _GEN_2234; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3004 = way0_hit ? recent_wdata1_49 : _GEN_2235; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3005 = way0_hit ? recent_wdata1_50 : _GEN_2236; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3006 = way0_hit ? recent_wdata1_51 : _GEN_2237; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3007 = way0_hit ? recent_wdata1_52 : _GEN_2238; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3008 = way0_hit ? recent_wdata1_53 : _GEN_2239; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3009 = way0_hit ? recent_wdata1_54 : _GEN_2240; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3010 = way0_hit ? recent_wdata1_55 : _GEN_2241; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3011 = way0_hit ? recent_wdata1_56 : _GEN_2242; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3012 = way0_hit ? recent_wdata1_57 : _GEN_2243; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3013 = way0_hit ? recent_wdata1_58 : _GEN_2244; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3014 = way0_hit ? recent_wdata1_59 : _GEN_2245; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3015 = way0_hit ? recent_wdata1_60 : _GEN_2246; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3016 = way0_hit ? recent_wdata1_61 : _GEN_2247; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3017 = way0_hit ? recent_wdata1_62 : _GEN_2248; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3018 = way0_hit ? recent_wdata1_63 : _GEN_2249; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3019 = way0_hit ? recent_wdata1_64 : _GEN_2250; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3020 = way0_hit ? recent_wdata1_65 : _GEN_2251; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3021 = way0_hit ? recent_wdata1_66 : _GEN_2252; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3022 = way0_hit ? recent_wdata1_67 : _GEN_2253; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3023 = way0_hit ? recent_wdata1_68 : _GEN_2254; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3024 = way0_hit ? recent_wdata1_69 : _GEN_2255; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3025 = way0_hit ? recent_wdata1_70 : _GEN_2256; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3026 = way0_hit ? recent_wdata1_71 : _GEN_2257; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3027 = way0_hit ? recent_wdata1_72 : _GEN_2258; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3028 = way0_hit ? recent_wdata1_73 : _GEN_2259; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3029 = way0_hit ? recent_wdata1_74 : _GEN_2260; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3030 = way0_hit ? recent_wdata1_75 : _GEN_2261; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3031 = way0_hit ? recent_wdata1_76 : _GEN_2262; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3032 = way0_hit ? recent_wdata1_77 : _GEN_2263; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3033 = way0_hit ? recent_wdata1_78 : _GEN_2264; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3034 = way0_hit ? recent_wdata1_79 : _GEN_2265; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3035 = way0_hit ? recent_wdata1_80 : _GEN_2266; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3036 = way0_hit ? recent_wdata1_81 : _GEN_2267; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3037 = way0_hit ? recent_wdata1_82 : _GEN_2268; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3038 = way0_hit ? recent_wdata1_83 : _GEN_2269; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3039 = way0_hit ? recent_wdata1_84 : _GEN_2270; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3040 = way0_hit ? recent_wdata1_85 : _GEN_2271; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3041 = way0_hit ? recent_wdata1_86 : _GEN_2272; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3042 = way0_hit ? recent_wdata1_87 : _GEN_2273; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3043 = way0_hit ? recent_wdata1_88 : _GEN_2274; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3044 = way0_hit ? recent_wdata1_89 : _GEN_2275; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3045 = way0_hit ? recent_wdata1_90 : _GEN_2276; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3046 = way0_hit ? recent_wdata1_91 : _GEN_2277; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3047 = way0_hit ? recent_wdata1_92 : _GEN_2278; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3048 = way0_hit ? recent_wdata1_93 : _GEN_2279; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3049 = way0_hit ? recent_wdata1_94 : _GEN_2280; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3050 = way0_hit ? recent_wdata1_95 : _GEN_2281; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3051 = way0_hit ? recent_wdata1_96 : _GEN_2282; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3052 = way0_hit ? recent_wdata1_97 : _GEN_2283; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3053 = way0_hit ? recent_wdata1_98 : _GEN_2284; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3054 = way0_hit ? recent_wdata1_99 : _GEN_2285; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3055 = way0_hit ? recent_wdata1_100 : _GEN_2286; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3056 = way0_hit ? recent_wdata1_101 : _GEN_2287; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3057 = way0_hit ? recent_wdata1_102 : _GEN_2288; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3058 = way0_hit ? recent_wdata1_103 : _GEN_2289; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3059 = way0_hit ? recent_wdata1_104 : _GEN_2290; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3060 = way0_hit ? recent_wdata1_105 : _GEN_2291; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3061 = way0_hit ? recent_wdata1_106 : _GEN_2292; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3062 = way0_hit ? recent_wdata1_107 : _GEN_2293; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3063 = way0_hit ? recent_wdata1_108 : _GEN_2294; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3064 = way0_hit ? recent_wdata1_109 : _GEN_2295; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3065 = way0_hit ? recent_wdata1_110 : _GEN_2296; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3066 = way0_hit ? recent_wdata1_111 : _GEN_2297; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3067 = way0_hit ? recent_wdata1_112 : _GEN_2298; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3068 = way0_hit ? recent_wdata1_113 : _GEN_2299; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3069 = way0_hit ? recent_wdata1_114 : _GEN_2300; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3070 = way0_hit ? recent_wdata1_115 : _GEN_2301; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3071 = way0_hit ? recent_wdata1_116 : _GEN_2302; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3072 = way0_hit ? recent_wdata1_117 : _GEN_2303; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3073 = way0_hit ? recent_wdata1_118 : _GEN_2304; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3074 = way0_hit ? recent_wdata1_119 : _GEN_2305; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3075 = way0_hit ? recent_wdata1_120 : _GEN_2306; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3076 = way0_hit ? recent_wdata1_121 : _GEN_2307; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3077 = way0_hit ? recent_wdata1_122 : _GEN_2308; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3078 = way0_hit ? recent_wdata1_123 : _GEN_2309; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3079 = way0_hit ? recent_wdata1_124 : _GEN_2310; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3080 = way0_hit ? recent_wdata1_125 : _GEN_2311; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3081 = way0_hit ? recent_wdata1_126 : _GEN_2312; // @[d_cache.scala 107:27 21:32]
  wire [63:0] _GEN_3082 = way0_hit ? recent_wdata1_127 : _GEN_2313; // @[d_cache.scala 107:27 21:32]
  wire  _GEN_3083 = way0_hit ? dirty_1_0 : _GEN_2314; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3084 = way0_hit ? dirty_1_1 : _GEN_2315; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3085 = way0_hit ? dirty_1_2 : _GEN_2316; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3086 = way0_hit ? dirty_1_3 : _GEN_2317; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3087 = way0_hit ? dirty_1_4 : _GEN_2318; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3088 = way0_hit ? dirty_1_5 : _GEN_2319; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3089 = way0_hit ? dirty_1_6 : _GEN_2320; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3090 = way0_hit ? dirty_1_7 : _GEN_2321; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3091 = way0_hit ? dirty_1_8 : _GEN_2322; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3092 = way0_hit ? dirty_1_9 : _GEN_2323; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3093 = way0_hit ? dirty_1_10 : _GEN_2324; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3094 = way0_hit ? dirty_1_11 : _GEN_2325; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3095 = way0_hit ? dirty_1_12 : _GEN_2326; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3096 = way0_hit ? dirty_1_13 : _GEN_2327; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3097 = way0_hit ? dirty_1_14 : _GEN_2328; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3098 = way0_hit ? dirty_1_15 : _GEN_2329; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3099 = way0_hit ? dirty_1_16 : _GEN_2330; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3100 = way0_hit ? dirty_1_17 : _GEN_2331; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3101 = way0_hit ? dirty_1_18 : _GEN_2332; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3102 = way0_hit ? dirty_1_19 : _GEN_2333; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3103 = way0_hit ? dirty_1_20 : _GEN_2334; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3104 = way0_hit ? dirty_1_21 : _GEN_2335; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3105 = way0_hit ? dirty_1_22 : _GEN_2336; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3106 = way0_hit ? dirty_1_23 : _GEN_2337; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3107 = way0_hit ? dirty_1_24 : _GEN_2338; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3108 = way0_hit ? dirty_1_25 : _GEN_2339; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3109 = way0_hit ? dirty_1_26 : _GEN_2340; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3110 = way0_hit ? dirty_1_27 : _GEN_2341; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3111 = way0_hit ? dirty_1_28 : _GEN_2342; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3112 = way0_hit ? dirty_1_29 : _GEN_2343; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3113 = way0_hit ? dirty_1_30 : _GEN_2344; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3114 = way0_hit ? dirty_1_31 : _GEN_2345; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3115 = way0_hit ? dirty_1_32 : _GEN_2346; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3116 = way0_hit ? dirty_1_33 : _GEN_2347; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3117 = way0_hit ? dirty_1_34 : _GEN_2348; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3118 = way0_hit ? dirty_1_35 : _GEN_2349; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3119 = way0_hit ? dirty_1_36 : _GEN_2350; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3120 = way0_hit ? dirty_1_37 : _GEN_2351; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3121 = way0_hit ? dirty_1_38 : _GEN_2352; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3122 = way0_hit ? dirty_1_39 : _GEN_2353; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3123 = way0_hit ? dirty_1_40 : _GEN_2354; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3124 = way0_hit ? dirty_1_41 : _GEN_2355; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3125 = way0_hit ? dirty_1_42 : _GEN_2356; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3126 = way0_hit ? dirty_1_43 : _GEN_2357; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3127 = way0_hit ? dirty_1_44 : _GEN_2358; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3128 = way0_hit ? dirty_1_45 : _GEN_2359; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3129 = way0_hit ? dirty_1_46 : _GEN_2360; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3130 = way0_hit ? dirty_1_47 : _GEN_2361; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3131 = way0_hit ? dirty_1_48 : _GEN_2362; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3132 = way0_hit ? dirty_1_49 : _GEN_2363; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3133 = way0_hit ? dirty_1_50 : _GEN_2364; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3134 = way0_hit ? dirty_1_51 : _GEN_2365; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3135 = way0_hit ? dirty_1_52 : _GEN_2366; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3136 = way0_hit ? dirty_1_53 : _GEN_2367; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3137 = way0_hit ? dirty_1_54 : _GEN_2368; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3138 = way0_hit ? dirty_1_55 : _GEN_2369; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3139 = way0_hit ? dirty_1_56 : _GEN_2370; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3140 = way0_hit ? dirty_1_57 : _GEN_2371; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3141 = way0_hit ? dirty_1_58 : _GEN_2372; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3142 = way0_hit ? dirty_1_59 : _GEN_2373; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3143 = way0_hit ? dirty_1_60 : _GEN_2374; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3144 = way0_hit ? dirty_1_61 : _GEN_2375; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3145 = way0_hit ? dirty_1_62 : _GEN_2376; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3146 = way0_hit ? dirty_1_63 : _GEN_2377; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3147 = way0_hit ? dirty_1_64 : _GEN_2378; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3148 = way0_hit ? dirty_1_65 : _GEN_2379; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3149 = way0_hit ? dirty_1_66 : _GEN_2380; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3150 = way0_hit ? dirty_1_67 : _GEN_2381; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3151 = way0_hit ? dirty_1_68 : _GEN_2382; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3152 = way0_hit ? dirty_1_69 : _GEN_2383; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3153 = way0_hit ? dirty_1_70 : _GEN_2384; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3154 = way0_hit ? dirty_1_71 : _GEN_2385; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3155 = way0_hit ? dirty_1_72 : _GEN_2386; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3156 = way0_hit ? dirty_1_73 : _GEN_2387; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3157 = way0_hit ? dirty_1_74 : _GEN_2388; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3158 = way0_hit ? dirty_1_75 : _GEN_2389; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3159 = way0_hit ? dirty_1_76 : _GEN_2390; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3160 = way0_hit ? dirty_1_77 : _GEN_2391; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3161 = way0_hit ? dirty_1_78 : _GEN_2392; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3162 = way0_hit ? dirty_1_79 : _GEN_2393; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3163 = way0_hit ? dirty_1_80 : _GEN_2394; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3164 = way0_hit ? dirty_1_81 : _GEN_2395; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3165 = way0_hit ? dirty_1_82 : _GEN_2396; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3166 = way0_hit ? dirty_1_83 : _GEN_2397; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3167 = way0_hit ? dirty_1_84 : _GEN_2398; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3168 = way0_hit ? dirty_1_85 : _GEN_2399; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3169 = way0_hit ? dirty_1_86 : _GEN_2400; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3170 = way0_hit ? dirty_1_87 : _GEN_2401; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3171 = way0_hit ? dirty_1_88 : _GEN_2402; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3172 = way0_hit ? dirty_1_89 : _GEN_2403; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3173 = way0_hit ? dirty_1_90 : _GEN_2404; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3174 = way0_hit ? dirty_1_91 : _GEN_2405; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3175 = way0_hit ? dirty_1_92 : _GEN_2406; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3176 = way0_hit ? dirty_1_93 : _GEN_2407; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3177 = way0_hit ? dirty_1_94 : _GEN_2408; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3178 = way0_hit ? dirty_1_95 : _GEN_2409; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3179 = way0_hit ? dirty_1_96 : _GEN_2410; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3180 = way0_hit ? dirty_1_97 : _GEN_2411; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3181 = way0_hit ? dirty_1_98 : _GEN_2412; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3182 = way0_hit ? dirty_1_99 : _GEN_2413; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3183 = way0_hit ? dirty_1_100 : _GEN_2414; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3184 = way0_hit ? dirty_1_101 : _GEN_2415; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3185 = way0_hit ? dirty_1_102 : _GEN_2416; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3186 = way0_hit ? dirty_1_103 : _GEN_2417; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3187 = way0_hit ? dirty_1_104 : _GEN_2418; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3188 = way0_hit ? dirty_1_105 : _GEN_2419; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3189 = way0_hit ? dirty_1_106 : _GEN_2420; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3190 = way0_hit ? dirty_1_107 : _GEN_2421; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3191 = way0_hit ? dirty_1_108 : _GEN_2422; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3192 = way0_hit ? dirty_1_109 : _GEN_2423; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3193 = way0_hit ? dirty_1_110 : _GEN_2424; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3194 = way0_hit ? dirty_1_111 : _GEN_2425; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3195 = way0_hit ? dirty_1_112 : _GEN_2426; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3196 = way0_hit ? dirty_1_113 : _GEN_2427; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3197 = way0_hit ? dirty_1_114 : _GEN_2428; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3198 = way0_hit ? dirty_1_115 : _GEN_2429; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3199 = way0_hit ? dirty_1_116 : _GEN_2430; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3200 = way0_hit ? dirty_1_117 : _GEN_2431; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3201 = way0_hit ? dirty_1_118 : _GEN_2432; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3202 = way0_hit ? dirty_1_119 : _GEN_2433; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3203 = way0_hit ? dirty_1_120 : _GEN_2434; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3204 = way0_hit ? dirty_1_121 : _GEN_2435; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3205 = way0_hit ? dirty_1_122 : _GEN_2436; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3206 = way0_hit ? dirty_1_123 : _GEN_2437; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3207 = way0_hit ? dirty_1_124 : _GEN_2438; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3208 = way0_hit ? dirty_1_125 : _GEN_2439; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3209 = way0_hit ? dirty_1_126 : _GEN_2440; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_3210 = way0_hit ? dirty_1_127 : _GEN_2441; // @[d_cache.scala 107:27 27:26]
  wire [2:0] _GEN_3211 = io_from_axi_rvalid ? 3'h5 : state; // @[d_cache.scala 126:37 127:23 76:24]
  wire [63:0] _GEN_3212 = io_from_axi_rvalid ? io_from_axi_rdata : receive_data; // @[d_cache.scala 129:37 130:30 36:31]
  wire [2:0] _GEN_3213 = io_from_axi_bvalid ? 3'h0 : state; // @[d_cache.scala 134:37 135:23 76:24]
  wire [63:0] _GEN_3214 = 7'h0 == index[6:0] ? receive_data : ram_0_0; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3215 = 7'h1 == index[6:0] ? receive_data : ram_0_1; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3216 = 7'h2 == index[6:0] ? receive_data : ram_0_2; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3217 = 7'h3 == index[6:0] ? receive_data : ram_0_3; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3218 = 7'h4 == index[6:0] ? receive_data : ram_0_4; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3219 = 7'h5 == index[6:0] ? receive_data : ram_0_5; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3220 = 7'h6 == index[6:0] ? receive_data : ram_0_6; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3221 = 7'h7 == index[6:0] ? receive_data : ram_0_7; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3222 = 7'h8 == index[6:0] ? receive_data : ram_0_8; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3223 = 7'h9 == index[6:0] ? receive_data : ram_0_9; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3224 = 7'ha == index[6:0] ? receive_data : ram_0_10; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3225 = 7'hb == index[6:0] ? receive_data : ram_0_11; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3226 = 7'hc == index[6:0] ? receive_data : ram_0_12; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3227 = 7'hd == index[6:0] ? receive_data : ram_0_13; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3228 = 7'he == index[6:0] ? receive_data : ram_0_14; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3229 = 7'hf == index[6:0] ? receive_data : ram_0_15; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3230 = 7'h10 == index[6:0] ? receive_data : ram_0_16; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3231 = 7'h11 == index[6:0] ? receive_data : ram_0_17; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3232 = 7'h12 == index[6:0] ? receive_data : ram_0_18; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3233 = 7'h13 == index[6:0] ? receive_data : ram_0_19; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3234 = 7'h14 == index[6:0] ? receive_data : ram_0_20; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3235 = 7'h15 == index[6:0] ? receive_data : ram_0_21; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3236 = 7'h16 == index[6:0] ? receive_data : ram_0_22; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3237 = 7'h17 == index[6:0] ? receive_data : ram_0_23; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3238 = 7'h18 == index[6:0] ? receive_data : ram_0_24; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3239 = 7'h19 == index[6:0] ? receive_data : ram_0_25; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3240 = 7'h1a == index[6:0] ? receive_data : ram_0_26; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3241 = 7'h1b == index[6:0] ? receive_data : ram_0_27; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3242 = 7'h1c == index[6:0] ? receive_data : ram_0_28; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3243 = 7'h1d == index[6:0] ? receive_data : ram_0_29; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3244 = 7'h1e == index[6:0] ? receive_data : ram_0_30; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3245 = 7'h1f == index[6:0] ? receive_data : ram_0_31; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3246 = 7'h20 == index[6:0] ? receive_data : ram_0_32; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3247 = 7'h21 == index[6:0] ? receive_data : ram_0_33; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3248 = 7'h22 == index[6:0] ? receive_data : ram_0_34; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3249 = 7'h23 == index[6:0] ? receive_data : ram_0_35; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3250 = 7'h24 == index[6:0] ? receive_data : ram_0_36; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3251 = 7'h25 == index[6:0] ? receive_data : ram_0_37; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3252 = 7'h26 == index[6:0] ? receive_data : ram_0_38; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3253 = 7'h27 == index[6:0] ? receive_data : ram_0_39; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3254 = 7'h28 == index[6:0] ? receive_data : ram_0_40; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3255 = 7'h29 == index[6:0] ? receive_data : ram_0_41; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3256 = 7'h2a == index[6:0] ? receive_data : ram_0_42; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3257 = 7'h2b == index[6:0] ? receive_data : ram_0_43; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3258 = 7'h2c == index[6:0] ? receive_data : ram_0_44; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3259 = 7'h2d == index[6:0] ? receive_data : ram_0_45; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3260 = 7'h2e == index[6:0] ? receive_data : ram_0_46; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3261 = 7'h2f == index[6:0] ? receive_data : ram_0_47; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3262 = 7'h30 == index[6:0] ? receive_data : ram_0_48; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3263 = 7'h31 == index[6:0] ? receive_data : ram_0_49; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3264 = 7'h32 == index[6:0] ? receive_data : ram_0_50; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3265 = 7'h33 == index[6:0] ? receive_data : ram_0_51; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3266 = 7'h34 == index[6:0] ? receive_data : ram_0_52; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3267 = 7'h35 == index[6:0] ? receive_data : ram_0_53; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3268 = 7'h36 == index[6:0] ? receive_data : ram_0_54; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3269 = 7'h37 == index[6:0] ? receive_data : ram_0_55; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3270 = 7'h38 == index[6:0] ? receive_data : ram_0_56; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3271 = 7'h39 == index[6:0] ? receive_data : ram_0_57; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3272 = 7'h3a == index[6:0] ? receive_data : ram_0_58; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3273 = 7'h3b == index[6:0] ? receive_data : ram_0_59; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3274 = 7'h3c == index[6:0] ? receive_data : ram_0_60; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3275 = 7'h3d == index[6:0] ? receive_data : ram_0_61; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3276 = 7'h3e == index[6:0] ? receive_data : ram_0_62; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3277 = 7'h3f == index[6:0] ? receive_data : ram_0_63; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3278 = 7'h40 == index[6:0] ? receive_data : ram_0_64; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3279 = 7'h41 == index[6:0] ? receive_data : ram_0_65; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3280 = 7'h42 == index[6:0] ? receive_data : ram_0_66; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3281 = 7'h43 == index[6:0] ? receive_data : ram_0_67; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3282 = 7'h44 == index[6:0] ? receive_data : ram_0_68; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3283 = 7'h45 == index[6:0] ? receive_data : ram_0_69; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3284 = 7'h46 == index[6:0] ? receive_data : ram_0_70; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3285 = 7'h47 == index[6:0] ? receive_data : ram_0_71; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3286 = 7'h48 == index[6:0] ? receive_data : ram_0_72; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3287 = 7'h49 == index[6:0] ? receive_data : ram_0_73; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3288 = 7'h4a == index[6:0] ? receive_data : ram_0_74; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3289 = 7'h4b == index[6:0] ? receive_data : ram_0_75; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3290 = 7'h4c == index[6:0] ? receive_data : ram_0_76; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3291 = 7'h4d == index[6:0] ? receive_data : ram_0_77; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3292 = 7'h4e == index[6:0] ? receive_data : ram_0_78; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3293 = 7'h4f == index[6:0] ? receive_data : ram_0_79; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3294 = 7'h50 == index[6:0] ? receive_data : ram_0_80; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3295 = 7'h51 == index[6:0] ? receive_data : ram_0_81; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3296 = 7'h52 == index[6:0] ? receive_data : ram_0_82; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3297 = 7'h53 == index[6:0] ? receive_data : ram_0_83; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3298 = 7'h54 == index[6:0] ? receive_data : ram_0_84; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3299 = 7'h55 == index[6:0] ? receive_data : ram_0_85; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3300 = 7'h56 == index[6:0] ? receive_data : ram_0_86; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3301 = 7'h57 == index[6:0] ? receive_data : ram_0_87; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3302 = 7'h58 == index[6:0] ? receive_data : ram_0_88; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3303 = 7'h59 == index[6:0] ? receive_data : ram_0_89; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3304 = 7'h5a == index[6:0] ? receive_data : ram_0_90; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3305 = 7'h5b == index[6:0] ? receive_data : ram_0_91; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3306 = 7'h5c == index[6:0] ? receive_data : ram_0_92; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3307 = 7'h5d == index[6:0] ? receive_data : ram_0_93; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3308 = 7'h5e == index[6:0] ? receive_data : ram_0_94; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3309 = 7'h5f == index[6:0] ? receive_data : ram_0_95; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3310 = 7'h60 == index[6:0] ? receive_data : ram_0_96; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3311 = 7'h61 == index[6:0] ? receive_data : ram_0_97; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3312 = 7'h62 == index[6:0] ? receive_data : ram_0_98; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3313 = 7'h63 == index[6:0] ? receive_data : ram_0_99; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3314 = 7'h64 == index[6:0] ? receive_data : ram_0_100; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3315 = 7'h65 == index[6:0] ? receive_data : ram_0_101; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3316 = 7'h66 == index[6:0] ? receive_data : ram_0_102; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3317 = 7'h67 == index[6:0] ? receive_data : ram_0_103; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3318 = 7'h68 == index[6:0] ? receive_data : ram_0_104; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3319 = 7'h69 == index[6:0] ? receive_data : ram_0_105; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3320 = 7'h6a == index[6:0] ? receive_data : ram_0_106; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3321 = 7'h6b == index[6:0] ? receive_data : ram_0_107; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3322 = 7'h6c == index[6:0] ? receive_data : ram_0_108; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3323 = 7'h6d == index[6:0] ? receive_data : ram_0_109; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3324 = 7'h6e == index[6:0] ? receive_data : ram_0_110; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3325 = 7'h6f == index[6:0] ? receive_data : ram_0_111; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3326 = 7'h70 == index[6:0] ? receive_data : ram_0_112; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3327 = 7'h71 == index[6:0] ? receive_data : ram_0_113; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3328 = 7'h72 == index[6:0] ? receive_data : ram_0_114; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3329 = 7'h73 == index[6:0] ? receive_data : ram_0_115; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3330 = 7'h74 == index[6:0] ? receive_data : ram_0_116; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3331 = 7'h75 == index[6:0] ? receive_data : ram_0_117; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3332 = 7'h76 == index[6:0] ? receive_data : ram_0_118; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3333 = 7'h77 == index[6:0] ? receive_data : ram_0_119; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3334 = 7'h78 == index[6:0] ? receive_data : ram_0_120; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3335 = 7'h79 == index[6:0] ? receive_data : ram_0_121; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3336 = 7'h7a == index[6:0] ? receive_data : ram_0_122; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3337 = 7'h7b == index[6:0] ? receive_data : ram_0_123; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3338 = 7'h7c == index[6:0] ? receive_data : ram_0_124; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3339 = 7'h7d == index[6:0] ? receive_data : ram_0_125; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3340 = 7'h7e == index[6:0] ? receive_data : ram_0_126; // @[d_cache.scala 141:{30,30} 18:24]
  wire [63:0] _GEN_3341 = 7'h7f == index[6:0] ? receive_data : ram_0_127; // @[d_cache.scala 141:{30,30} 18:24]
  wire [31:0] _GEN_3342 = 7'h0 == index[6:0] ? _GEN_18465 : tag_0_0; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3343 = 7'h1 == index[6:0] ? _GEN_18465 : tag_0_1; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3344 = 7'h2 == index[6:0] ? _GEN_18465 : tag_0_2; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3345 = 7'h3 == index[6:0] ? _GEN_18465 : tag_0_3; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3346 = 7'h4 == index[6:0] ? _GEN_18465 : tag_0_4; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3347 = 7'h5 == index[6:0] ? _GEN_18465 : tag_0_5; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3348 = 7'h6 == index[6:0] ? _GEN_18465 : tag_0_6; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3349 = 7'h7 == index[6:0] ? _GEN_18465 : tag_0_7; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3350 = 7'h8 == index[6:0] ? _GEN_18465 : tag_0_8; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3351 = 7'h9 == index[6:0] ? _GEN_18465 : tag_0_9; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3352 = 7'ha == index[6:0] ? _GEN_18465 : tag_0_10; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3353 = 7'hb == index[6:0] ? _GEN_18465 : tag_0_11; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3354 = 7'hc == index[6:0] ? _GEN_18465 : tag_0_12; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3355 = 7'hd == index[6:0] ? _GEN_18465 : tag_0_13; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3356 = 7'he == index[6:0] ? _GEN_18465 : tag_0_14; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3357 = 7'hf == index[6:0] ? _GEN_18465 : tag_0_15; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3358 = 7'h10 == index[6:0] ? _GEN_18465 : tag_0_16; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3359 = 7'h11 == index[6:0] ? _GEN_18465 : tag_0_17; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3360 = 7'h12 == index[6:0] ? _GEN_18465 : tag_0_18; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3361 = 7'h13 == index[6:0] ? _GEN_18465 : tag_0_19; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3362 = 7'h14 == index[6:0] ? _GEN_18465 : tag_0_20; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3363 = 7'h15 == index[6:0] ? _GEN_18465 : tag_0_21; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3364 = 7'h16 == index[6:0] ? _GEN_18465 : tag_0_22; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3365 = 7'h17 == index[6:0] ? _GEN_18465 : tag_0_23; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3366 = 7'h18 == index[6:0] ? _GEN_18465 : tag_0_24; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3367 = 7'h19 == index[6:0] ? _GEN_18465 : tag_0_25; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3368 = 7'h1a == index[6:0] ? _GEN_18465 : tag_0_26; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3369 = 7'h1b == index[6:0] ? _GEN_18465 : tag_0_27; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3370 = 7'h1c == index[6:0] ? _GEN_18465 : tag_0_28; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3371 = 7'h1d == index[6:0] ? _GEN_18465 : tag_0_29; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3372 = 7'h1e == index[6:0] ? _GEN_18465 : tag_0_30; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3373 = 7'h1f == index[6:0] ? _GEN_18465 : tag_0_31; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3374 = 7'h20 == index[6:0] ? _GEN_18465 : tag_0_32; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3375 = 7'h21 == index[6:0] ? _GEN_18465 : tag_0_33; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3376 = 7'h22 == index[6:0] ? _GEN_18465 : tag_0_34; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3377 = 7'h23 == index[6:0] ? _GEN_18465 : tag_0_35; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3378 = 7'h24 == index[6:0] ? _GEN_18465 : tag_0_36; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3379 = 7'h25 == index[6:0] ? _GEN_18465 : tag_0_37; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3380 = 7'h26 == index[6:0] ? _GEN_18465 : tag_0_38; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3381 = 7'h27 == index[6:0] ? _GEN_18465 : tag_0_39; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3382 = 7'h28 == index[6:0] ? _GEN_18465 : tag_0_40; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3383 = 7'h29 == index[6:0] ? _GEN_18465 : tag_0_41; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3384 = 7'h2a == index[6:0] ? _GEN_18465 : tag_0_42; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3385 = 7'h2b == index[6:0] ? _GEN_18465 : tag_0_43; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3386 = 7'h2c == index[6:0] ? _GEN_18465 : tag_0_44; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3387 = 7'h2d == index[6:0] ? _GEN_18465 : tag_0_45; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3388 = 7'h2e == index[6:0] ? _GEN_18465 : tag_0_46; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3389 = 7'h2f == index[6:0] ? _GEN_18465 : tag_0_47; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3390 = 7'h30 == index[6:0] ? _GEN_18465 : tag_0_48; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3391 = 7'h31 == index[6:0] ? _GEN_18465 : tag_0_49; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3392 = 7'h32 == index[6:0] ? _GEN_18465 : tag_0_50; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3393 = 7'h33 == index[6:0] ? _GEN_18465 : tag_0_51; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3394 = 7'h34 == index[6:0] ? _GEN_18465 : tag_0_52; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3395 = 7'h35 == index[6:0] ? _GEN_18465 : tag_0_53; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3396 = 7'h36 == index[6:0] ? _GEN_18465 : tag_0_54; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3397 = 7'h37 == index[6:0] ? _GEN_18465 : tag_0_55; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3398 = 7'h38 == index[6:0] ? _GEN_18465 : tag_0_56; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3399 = 7'h39 == index[6:0] ? _GEN_18465 : tag_0_57; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3400 = 7'h3a == index[6:0] ? _GEN_18465 : tag_0_58; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3401 = 7'h3b == index[6:0] ? _GEN_18465 : tag_0_59; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3402 = 7'h3c == index[6:0] ? _GEN_18465 : tag_0_60; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3403 = 7'h3d == index[6:0] ? _GEN_18465 : tag_0_61; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3404 = 7'h3e == index[6:0] ? _GEN_18465 : tag_0_62; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3405 = 7'h3f == index[6:0] ? _GEN_18465 : tag_0_63; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3406 = 7'h40 == index[6:0] ? _GEN_18465 : tag_0_64; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3407 = 7'h41 == index[6:0] ? _GEN_18465 : tag_0_65; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3408 = 7'h42 == index[6:0] ? _GEN_18465 : tag_0_66; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3409 = 7'h43 == index[6:0] ? _GEN_18465 : tag_0_67; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3410 = 7'h44 == index[6:0] ? _GEN_18465 : tag_0_68; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3411 = 7'h45 == index[6:0] ? _GEN_18465 : tag_0_69; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3412 = 7'h46 == index[6:0] ? _GEN_18465 : tag_0_70; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3413 = 7'h47 == index[6:0] ? _GEN_18465 : tag_0_71; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3414 = 7'h48 == index[6:0] ? _GEN_18465 : tag_0_72; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3415 = 7'h49 == index[6:0] ? _GEN_18465 : tag_0_73; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3416 = 7'h4a == index[6:0] ? _GEN_18465 : tag_0_74; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3417 = 7'h4b == index[6:0] ? _GEN_18465 : tag_0_75; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3418 = 7'h4c == index[6:0] ? _GEN_18465 : tag_0_76; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3419 = 7'h4d == index[6:0] ? _GEN_18465 : tag_0_77; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3420 = 7'h4e == index[6:0] ? _GEN_18465 : tag_0_78; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3421 = 7'h4f == index[6:0] ? _GEN_18465 : tag_0_79; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3422 = 7'h50 == index[6:0] ? _GEN_18465 : tag_0_80; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3423 = 7'h51 == index[6:0] ? _GEN_18465 : tag_0_81; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3424 = 7'h52 == index[6:0] ? _GEN_18465 : tag_0_82; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3425 = 7'h53 == index[6:0] ? _GEN_18465 : tag_0_83; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3426 = 7'h54 == index[6:0] ? _GEN_18465 : tag_0_84; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3427 = 7'h55 == index[6:0] ? _GEN_18465 : tag_0_85; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3428 = 7'h56 == index[6:0] ? _GEN_18465 : tag_0_86; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3429 = 7'h57 == index[6:0] ? _GEN_18465 : tag_0_87; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3430 = 7'h58 == index[6:0] ? _GEN_18465 : tag_0_88; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3431 = 7'h59 == index[6:0] ? _GEN_18465 : tag_0_89; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3432 = 7'h5a == index[6:0] ? _GEN_18465 : tag_0_90; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3433 = 7'h5b == index[6:0] ? _GEN_18465 : tag_0_91; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3434 = 7'h5c == index[6:0] ? _GEN_18465 : tag_0_92; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3435 = 7'h5d == index[6:0] ? _GEN_18465 : tag_0_93; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3436 = 7'h5e == index[6:0] ? _GEN_18465 : tag_0_94; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3437 = 7'h5f == index[6:0] ? _GEN_18465 : tag_0_95; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3438 = 7'h60 == index[6:0] ? _GEN_18465 : tag_0_96; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3439 = 7'h61 == index[6:0] ? _GEN_18465 : tag_0_97; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3440 = 7'h62 == index[6:0] ? _GEN_18465 : tag_0_98; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3441 = 7'h63 == index[6:0] ? _GEN_18465 : tag_0_99; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3442 = 7'h64 == index[6:0] ? _GEN_18465 : tag_0_100; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3443 = 7'h65 == index[6:0] ? _GEN_18465 : tag_0_101; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3444 = 7'h66 == index[6:0] ? _GEN_18465 : tag_0_102; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3445 = 7'h67 == index[6:0] ? _GEN_18465 : tag_0_103; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3446 = 7'h68 == index[6:0] ? _GEN_18465 : tag_0_104; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3447 = 7'h69 == index[6:0] ? _GEN_18465 : tag_0_105; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3448 = 7'h6a == index[6:0] ? _GEN_18465 : tag_0_106; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3449 = 7'h6b == index[6:0] ? _GEN_18465 : tag_0_107; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3450 = 7'h6c == index[6:0] ? _GEN_18465 : tag_0_108; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3451 = 7'h6d == index[6:0] ? _GEN_18465 : tag_0_109; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3452 = 7'h6e == index[6:0] ? _GEN_18465 : tag_0_110; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3453 = 7'h6f == index[6:0] ? _GEN_18465 : tag_0_111; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3454 = 7'h70 == index[6:0] ? _GEN_18465 : tag_0_112; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3455 = 7'h71 == index[6:0] ? _GEN_18465 : tag_0_113; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3456 = 7'h72 == index[6:0] ? _GEN_18465 : tag_0_114; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3457 = 7'h73 == index[6:0] ? _GEN_18465 : tag_0_115; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3458 = 7'h74 == index[6:0] ? _GEN_18465 : tag_0_116; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3459 = 7'h75 == index[6:0] ? _GEN_18465 : tag_0_117; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3460 = 7'h76 == index[6:0] ? _GEN_18465 : tag_0_118; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3461 = 7'h77 == index[6:0] ? _GEN_18465 : tag_0_119; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3462 = 7'h78 == index[6:0] ? _GEN_18465 : tag_0_120; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3463 = 7'h79 == index[6:0] ? _GEN_18465 : tag_0_121; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3464 = 7'h7a == index[6:0] ? _GEN_18465 : tag_0_122; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3465 = 7'h7b == index[6:0] ? _GEN_18465 : tag_0_123; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3466 = 7'h7c == index[6:0] ? _GEN_18465 : tag_0_124; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3467 = 7'h7d == index[6:0] ? _GEN_18465 : tag_0_125; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3468 = 7'h7e == index[6:0] ? _GEN_18465 : tag_0_126; // @[d_cache.scala 142:{30,30} 22:24]
  wire [31:0] _GEN_3469 = 7'h7f == index[6:0] ? _GEN_18465 : tag_0_127; // @[d_cache.scala 142:{30,30} 22:24]
  wire  _GEN_3470 = _GEN_18470 | valid_0_0; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3471 = _GEN_18471 | valid_0_1; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3472 = _GEN_18472 | valid_0_2; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3473 = _GEN_18473 | valid_0_3; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3474 = _GEN_18474 | valid_0_4; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3475 = _GEN_18475 | valid_0_5; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3476 = _GEN_18476 | valid_0_6; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3477 = _GEN_18477 | valid_0_7; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3478 = _GEN_18478 | valid_0_8; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3479 = _GEN_18479 | valid_0_9; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3480 = _GEN_18480 | valid_0_10; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3481 = _GEN_18481 | valid_0_11; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3482 = _GEN_18482 | valid_0_12; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3483 = _GEN_18483 | valid_0_13; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3484 = _GEN_18484 | valid_0_14; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3485 = _GEN_18485 | valid_0_15; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3486 = _GEN_18486 | valid_0_16; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3487 = _GEN_18487 | valid_0_17; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3488 = _GEN_18488 | valid_0_18; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3489 = _GEN_18489 | valid_0_19; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3490 = _GEN_18490 | valid_0_20; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3491 = _GEN_18491 | valid_0_21; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3492 = _GEN_18492 | valid_0_22; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3493 = _GEN_18493 | valid_0_23; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3494 = _GEN_18494 | valid_0_24; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3495 = _GEN_18495 | valid_0_25; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3496 = _GEN_18496 | valid_0_26; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3497 = _GEN_18497 | valid_0_27; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3498 = _GEN_18498 | valid_0_28; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3499 = _GEN_18499 | valid_0_29; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3500 = _GEN_18500 | valid_0_30; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3501 = _GEN_18501 | valid_0_31; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3502 = _GEN_18502 | valid_0_32; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3503 = _GEN_18503 | valid_0_33; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3504 = _GEN_18504 | valid_0_34; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3505 = _GEN_18505 | valid_0_35; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3506 = _GEN_18506 | valid_0_36; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3507 = _GEN_18507 | valid_0_37; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3508 = _GEN_18508 | valid_0_38; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3509 = _GEN_18509 | valid_0_39; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3510 = _GEN_18510 | valid_0_40; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3511 = _GEN_18511 | valid_0_41; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3512 = _GEN_18512 | valid_0_42; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3513 = _GEN_18513 | valid_0_43; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3514 = _GEN_18514 | valid_0_44; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3515 = _GEN_18515 | valid_0_45; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3516 = _GEN_18516 | valid_0_46; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3517 = _GEN_18517 | valid_0_47; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3518 = _GEN_18518 | valid_0_48; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3519 = _GEN_18519 | valid_0_49; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3520 = _GEN_18520 | valid_0_50; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3521 = _GEN_18521 | valid_0_51; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3522 = _GEN_18522 | valid_0_52; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3523 = _GEN_18523 | valid_0_53; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3524 = _GEN_18524 | valid_0_54; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3525 = _GEN_18525 | valid_0_55; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3526 = _GEN_18526 | valid_0_56; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3527 = _GEN_18527 | valid_0_57; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3528 = _GEN_18528 | valid_0_58; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3529 = _GEN_18529 | valid_0_59; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3530 = _GEN_18530 | valid_0_60; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3531 = _GEN_18531 | valid_0_61; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3532 = _GEN_18532 | valid_0_62; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3533 = _GEN_18533 | valid_0_63; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3534 = _GEN_18534 | valid_0_64; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3535 = _GEN_18535 | valid_0_65; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3536 = _GEN_18536 | valid_0_66; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3537 = _GEN_18537 | valid_0_67; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3538 = _GEN_18538 | valid_0_68; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3539 = _GEN_18539 | valid_0_69; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3540 = _GEN_18540 | valid_0_70; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3541 = _GEN_18541 | valid_0_71; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3542 = _GEN_18542 | valid_0_72; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3543 = _GEN_18543 | valid_0_73; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3544 = _GEN_18544 | valid_0_74; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3545 = _GEN_18545 | valid_0_75; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3546 = _GEN_18546 | valid_0_76; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3547 = _GEN_18547 | valid_0_77; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3548 = _GEN_18548 | valid_0_78; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3549 = _GEN_18549 | valid_0_79; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3550 = _GEN_18550 | valid_0_80; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3551 = _GEN_18551 | valid_0_81; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3552 = _GEN_18552 | valid_0_82; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3553 = _GEN_18553 | valid_0_83; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3554 = _GEN_18554 | valid_0_84; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3555 = _GEN_18555 | valid_0_85; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3556 = _GEN_18556 | valid_0_86; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3557 = _GEN_18557 | valid_0_87; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3558 = _GEN_18558 | valid_0_88; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3559 = _GEN_18559 | valid_0_89; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3560 = _GEN_18560 | valid_0_90; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3561 = _GEN_18561 | valid_0_91; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3562 = _GEN_18562 | valid_0_92; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3563 = _GEN_18563 | valid_0_93; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3564 = _GEN_18564 | valid_0_94; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3565 = _GEN_18565 | valid_0_95; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3566 = _GEN_18566 | valid_0_96; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3567 = _GEN_18567 | valid_0_97; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3568 = _GEN_18568 | valid_0_98; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3569 = _GEN_18569 | valid_0_99; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3570 = _GEN_18570 | valid_0_100; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3571 = _GEN_18571 | valid_0_101; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3572 = _GEN_18572 | valid_0_102; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3573 = _GEN_18573 | valid_0_103; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3574 = _GEN_18574 | valid_0_104; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3575 = _GEN_18575 | valid_0_105; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3576 = _GEN_18576 | valid_0_106; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3577 = _GEN_18577 | valid_0_107; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3578 = _GEN_18578 | valid_0_108; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3579 = _GEN_18579 | valid_0_109; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3580 = _GEN_18580 | valid_0_110; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3581 = _GEN_18581 | valid_0_111; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3582 = _GEN_18582 | valid_0_112; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3583 = _GEN_18583 | valid_0_113; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3584 = _GEN_18584 | valid_0_114; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3585 = _GEN_18585 | valid_0_115; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3586 = _GEN_18586 | valid_0_116; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3587 = _GEN_18587 | valid_0_117; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3588 = _GEN_18588 | valid_0_118; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3589 = _GEN_18589 | valid_0_119; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3590 = _GEN_18590 | valid_0_120; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3591 = _GEN_18591 | valid_0_121; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3592 = _GEN_18592 | valid_0_122; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3593 = _GEN_18593 | valid_0_123; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3594 = _GEN_18594 | valid_0_124; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3595 = _GEN_18595 | valid_0_125; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3596 = _GEN_18596 | valid_0_126; // @[d_cache.scala 143:{32,32} 24:26]
  wire  _GEN_3597 = _GEN_18597 | valid_0_127; // @[d_cache.scala 143:{32,32} 24:26]
  wire [63:0] _GEN_3598 = 7'h0 == index[6:0] ? receive_data : ram_1_0; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3599 = 7'h1 == index[6:0] ? receive_data : ram_1_1; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3600 = 7'h2 == index[6:0] ? receive_data : ram_1_2; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3601 = 7'h3 == index[6:0] ? receive_data : ram_1_3; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3602 = 7'h4 == index[6:0] ? receive_data : ram_1_4; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3603 = 7'h5 == index[6:0] ? receive_data : ram_1_5; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3604 = 7'h6 == index[6:0] ? receive_data : ram_1_6; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3605 = 7'h7 == index[6:0] ? receive_data : ram_1_7; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3606 = 7'h8 == index[6:0] ? receive_data : ram_1_8; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3607 = 7'h9 == index[6:0] ? receive_data : ram_1_9; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3608 = 7'ha == index[6:0] ? receive_data : ram_1_10; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3609 = 7'hb == index[6:0] ? receive_data : ram_1_11; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3610 = 7'hc == index[6:0] ? receive_data : ram_1_12; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3611 = 7'hd == index[6:0] ? receive_data : ram_1_13; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3612 = 7'he == index[6:0] ? receive_data : ram_1_14; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3613 = 7'hf == index[6:0] ? receive_data : ram_1_15; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3614 = 7'h10 == index[6:0] ? receive_data : ram_1_16; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3615 = 7'h11 == index[6:0] ? receive_data : ram_1_17; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3616 = 7'h12 == index[6:0] ? receive_data : ram_1_18; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3617 = 7'h13 == index[6:0] ? receive_data : ram_1_19; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3618 = 7'h14 == index[6:0] ? receive_data : ram_1_20; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3619 = 7'h15 == index[6:0] ? receive_data : ram_1_21; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3620 = 7'h16 == index[6:0] ? receive_data : ram_1_22; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3621 = 7'h17 == index[6:0] ? receive_data : ram_1_23; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3622 = 7'h18 == index[6:0] ? receive_data : ram_1_24; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3623 = 7'h19 == index[6:0] ? receive_data : ram_1_25; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3624 = 7'h1a == index[6:0] ? receive_data : ram_1_26; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3625 = 7'h1b == index[6:0] ? receive_data : ram_1_27; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3626 = 7'h1c == index[6:0] ? receive_data : ram_1_28; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3627 = 7'h1d == index[6:0] ? receive_data : ram_1_29; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3628 = 7'h1e == index[6:0] ? receive_data : ram_1_30; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3629 = 7'h1f == index[6:0] ? receive_data : ram_1_31; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3630 = 7'h20 == index[6:0] ? receive_data : ram_1_32; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3631 = 7'h21 == index[6:0] ? receive_data : ram_1_33; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3632 = 7'h22 == index[6:0] ? receive_data : ram_1_34; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3633 = 7'h23 == index[6:0] ? receive_data : ram_1_35; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3634 = 7'h24 == index[6:0] ? receive_data : ram_1_36; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3635 = 7'h25 == index[6:0] ? receive_data : ram_1_37; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3636 = 7'h26 == index[6:0] ? receive_data : ram_1_38; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3637 = 7'h27 == index[6:0] ? receive_data : ram_1_39; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3638 = 7'h28 == index[6:0] ? receive_data : ram_1_40; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3639 = 7'h29 == index[6:0] ? receive_data : ram_1_41; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3640 = 7'h2a == index[6:0] ? receive_data : ram_1_42; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3641 = 7'h2b == index[6:0] ? receive_data : ram_1_43; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3642 = 7'h2c == index[6:0] ? receive_data : ram_1_44; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3643 = 7'h2d == index[6:0] ? receive_data : ram_1_45; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3644 = 7'h2e == index[6:0] ? receive_data : ram_1_46; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3645 = 7'h2f == index[6:0] ? receive_data : ram_1_47; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3646 = 7'h30 == index[6:0] ? receive_data : ram_1_48; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3647 = 7'h31 == index[6:0] ? receive_data : ram_1_49; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3648 = 7'h32 == index[6:0] ? receive_data : ram_1_50; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3649 = 7'h33 == index[6:0] ? receive_data : ram_1_51; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3650 = 7'h34 == index[6:0] ? receive_data : ram_1_52; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3651 = 7'h35 == index[6:0] ? receive_data : ram_1_53; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3652 = 7'h36 == index[6:0] ? receive_data : ram_1_54; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3653 = 7'h37 == index[6:0] ? receive_data : ram_1_55; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3654 = 7'h38 == index[6:0] ? receive_data : ram_1_56; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3655 = 7'h39 == index[6:0] ? receive_data : ram_1_57; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3656 = 7'h3a == index[6:0] ? receive_data : ram_1_58; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3657 = 7'h3b == index[6:0] ? receive_data : ram_1_59; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3658 = 7'h3c == index[6:0] ? receive_data : ram_1_60; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3659 = 7'h3d == index[6:0] ? receive_data : ram_1_61; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3660 = 7'h3e == index[6:0] ? receive_data : ram_1_62; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3661 = 7'h3f == index[6:0] ? receive_data : ram_1_63; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3662 = 7'h40 == index[6:0] ? receive_data : ram_1_64; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3663 = 7'h41 == index[6:0] ? receive_data : ram_1_65; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3664 = 7'h42 == index[6:0] ? receive_data : ram_1_66; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3665 = 7'h43 == index[6:0] ? receive_data : ram_1_67; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3666 = 7'h44 == index[6:0] ? receive_data : ram_1_68; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3667 = 7'h45 == index[6:0] ? receive_data : ram_1_69; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3668 = 7'h46 == index[6:0] ? receive_data : ram_1_70; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3669 = 7'h47 == index[6:0] ? receive_data : ram_1_71; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3670 = 7'h48 == index[6:0] ? receive_data : ram_1_72; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3671 = 7'h49 == index[6:0] ? receive_data : ram_1_73; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3672 = 7'h4a == index[6:0] ? receive_data : ram_1_74; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3673 = 7'h4b == index[6:0] ? receive_data : ram_1_75; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3674 = 7'h4c == index[6:0] ? receive_data : ram_1_76; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3675 = 7'h4d == index[6:0] ? receive_data : ram_1_77; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3676 = 7'h4e == index[6:0] ? receive_data : ram_1_78; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3677 = 7'h4f == index[6:0] ? receive_data : ram_1_79; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3678 = 7'h50 == index[6:0] ? receive_data : ram_1_80; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3679 = 7'h51 == index[6:0] ? receive_data : ram_1_81; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3680 = 7'h52 == index[6:0] ? receive_data : ram_1_82; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3681 = 7'h53 == index[6:0] ? receive_data : ram_1_83; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3682 = 7'h54 == index[6:0] ? receive_data : ram_1_84; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3683 = 7'h55 == index[6:0] ? receive_data : ram_1_85; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3684 = 7'h56 == index[6:0] ? receive_data : ram_1_86; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3685 = 7'h57 == index[6:0] ? receive_data : ram_1_87; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3686 = 7'h58 == index[6:0] ? receive_data : ram_1_88; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3687 = 7'h59 == index[6:0] ? receive_data : ram_1_89; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3688 = 7'h5a == index[6:0] ? receive_data : ram_1_90; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3689 = 7'h5b == index[6:0] ? receive_data : ram_1_91; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3690 = 7'h5c == index[6:0] ? receive_data : ram_1_92; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3691 = 7'h5d == index[6:0] ? receive_data : ram_1_93; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3692 = 7'h5e == index[6:0] ? receive_data : ram_1_94; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3693 = 7'h5f == index[6:0] ? receive_data : ram_1_95; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3694 = 7'h60 == index[6:0] ? receive_data : ram_1_96; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3695 = 7'h61 == index[6:0] ? receive_data : ram_1_97; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3696 = 7'h62 == index[6:0] ? receive_data : ram_1_98; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3697 = 7'h63 == index[6:0] ? receive_data : ram_1_99; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3698 = 7'h64 == index[6:0] ? receive_data : ram_1_100; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3699 = 7'h65 == index[6:0] ? receive_data : ram_1_101; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3700 = 7'h66 == index[6:0] ? receive_data : ram_1_102; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3701 = 7'h67 == index[6:0] ? receive_data : ram_1_103; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3702 = 7'h68 == index[6:0] ? receive_data : ram_1_104; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3703 = 7'h69 == index[6:0] ? receive_data : ram_1_105; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3704 = 7'h6a == index[6:0] ? receive_data : ram_1_106; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3705 = 7'h6b == index[6:0] ? receive_data : ram_1_107; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3706 = 7'h6c == index[6:0] ? receive_data : ram_1_108; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3707 = 7'h6d == index[6:0] ? receive_data : ram_1_109; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3708 = 7'h6e == index[6:0] ? receive_data : ram_1_110; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3709 = 7'h6f == index[6:0] ? receive_data : ram_1_111; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3710 = 7'h70 == index[6:0] ? receive_data : ram_1_112; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3711 = 7'h71 == index[6:0] ? receive_data : ram_1_113; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3712 = 7'h72 == index[6:0] ? receive_data : ram_1_114; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3713 = 7'h73 == index[6:0] ? receive_data : ram_1_115; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3714 = 7'h74 == index[6:0] ? receive_data : ram_1_116; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3715 = 7'h75 == index[6:0] ? receive_data : ram_1_117; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3716 = 7'h76 == index[6:0] ? receive_data : ram_1_118; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3717 = 7'h77 == index[6:0] ? receive_data : ram_1_119; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3718 = 7'h78 == index[6:0] ? receive_data : ram_1_120; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3719 = 7'h79 == index[6:0] ? receive_data : ram_1_121; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3720 = 7'h7a == index[6:0] ? receive_data : ram_1_122; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3721 = 7'h7b == index[6:0] ? receive_data : ram_1_123; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3722 = 7'h7c == index[6:0] ? receive_data : ram_1_124; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3723 = 7'h7d == index[6:0] ? receive_data : ram_1_125; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3724 = 7'h7e == index[6:0] ? receive_data : ram_1_126; // @[d_cache.scala 147:{30,30} 19:24]
  wire [63:0] _GEN_3725 = 7'h7f == index[6:0] ? receive_data : ram_1_127; // @[d_cache.scala 147:{30,30} 19:24]
  wire [31:0] _GEN_3726 = 7'h0 == index[6:0] ? _GEN_18465 : tag_1_0; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3727 = 7'h1 == index[6:0] ? _GEN_18465 : tag_1_1; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3728 = 7'h2 == index[6:0] ? _GEN_18465 : tag_1_2; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3729 = 7'h3 == index[6:0] ? _GEN_18465 : tag_1_3; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3730 = 7'h4 == index[6:0] ? _GEN_18465 : tag_1_4; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3731 = 7'h5 == index[6:0] ? _GEN_18465 : tag_1_5; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3732 = 7'h6 == index[6:0] ? _GEN_18465 : tag_1_6; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3733 = 7'h7 == index[6:0] ? _GEN_18465 : tag_1_7; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3734 = 7'h8 == index[6:0] ? _GEN_18465 : tag_1_8; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3735 = 7'h9 == index[6:0] ? _GEN_18465 : tag_1_9; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3736 = 7'ha == index[6:0] ? _GEN_18465 : tag_1_10; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3737 = 7'hb == index[6:0] ? _GEN_18465 : tag_1_11; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3738 = 7'hc == index[6:0] ? _GEN_18465 : tag_1_12; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3739 = 7'hd == index[6:0] ? _GEN_18465 : tag_1_13; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3740 = 7'he == index[6:0] ? _GEN_18465 : tag_1_14; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3741 = 7'hf == index[6:0] ? _GEN_18465 : tag_1_15; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3742 = 7'h10 == index[6:0] ? _GEN_18465 : tag_1_16; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3743 = 7'h11 == index[6:0] ? _GEN_18465 : tag_1_17; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3744 = 7'h12 == index[6:0] ? _GEN_18465 : tag_1_18; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3745 = 7'h13 == index[6:0] ? _GEN_18465 : tag_1_19; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3746 = 7'h14 == index[6:0] ? _GEN_18465 : tag_1_20; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3747 = 7'h15 == index[6:0] ? _GEN_18465 : tag_1_21; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3748 = 7'h16 == index[6:0] ? _GEN_18465 : tag_1_22; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3749 = 7'h17 == index[6:0] ? _GEN_18465 : tag_1_23; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3750 = 7'h18 == index[6:0] ? _GEN_18465 : tag_1_24; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3751 = 7'h19 == index[6:0] ? _GEN_18465 : tag_1_25; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3752 = 7'h1a == index[6:0] ? _GEN_18465 : tag_1_26; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3753 = 7'h1b == index[6:0] ? _GEN_18465 : tag_1_27; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3754 = 7'h1c == index[6:0] ? _GEN_18465 : tag_1_28; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3755 = 7'h1d == index[6:0] ? _GEN_18465 : tag_1_29; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3756 = 7'h1e == index[6:0] ? _GEN_18465 : tag_1_30; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3757 = 7'h1f == index[6:0] ? _GEN_18465 : tag_1_31; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3758 = 7'h20 == index[6:0] ? _GEN_18465 : tag_1_32; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3759 = 7'h21 == index[6:0] ? _GEN_18465 : tag_1_33; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3760 = 7'h22 == index[6:0] ? _GEN_18465 : tag_1_34; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3761 = 7'h23 == index[6:0] ? _GEN_18465 : tag_1_35; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3762 = 7'h24 == index[6:0] ? _GEN_18465 : tag_1_36; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3763 = 7'h25 == index[6:0] ? _GEN_18465 : tag_1_37; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3764 = 7'h26 == index[6:0] ? _GEN_18465 : tag_1_38; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3765 = 7'h27 == index[6:0] ? _GEN_18465 : tag_1_39; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3766 = 7'h28 == index[6:0] ? _GEN_18465 : tag_1_40; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3767 = 7'h29 == index[6:0] ? _GEN_18465 : tag_1_41; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3768 = 7'h2a == index[6:0] ? _GEN_18465 : tag_1_42; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3769 = 7'h2b == index[6:0] ? _GEN_18465 : tag_1_43; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3770 = 7'h2c == index[6:0] ? _GEN_18465 : tag_1_44; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3771 = 7'h2d == index[6:0] ? _GEN_18465 : tag_1_45; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3772 = 7'h2e == index[6:0] ? _GEN_18465 : tag_1_46; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3773 = 7'h2f == index[6:0] ? _GEN_18465 : tag_1_47; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3774 = 7'h30 == index[6:0] ? _GEN_18465 : tag_1_48; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3775 = 7'h31 == index[6:0] ? _GEN_18465 : tag_1_49; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3776 = 7'h32 == index[6:0] ? _GEN_18465 : tag_1_50; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3777 = 7'h33 == index[6:0] ? _GEN_18465 : tag_1_51; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3778 = 7'h34 == index[6:0] ? _GEN_18465 : tag_1_52; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3779 = 7'h35 == index[6:0] ? _GEN_18465 : tag_1_53; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3780 = 7'h36 == index[6:0] ? _GEN_18465 : tag_1_54; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3781 = 7'h37 == index[6:0] ? _GEN_18465 : tag_1_55; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3782 = 7'h38 == index[6:0] ? _GEN_18465 : tag_1_56; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3783 = 7'h39 == index[6:0] ? _GEN_18465 : tag_1_57; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3784 = 7'h3a == index[6:0] ? _GEN_18465 : tag_1_58; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3785 = 7'h3b == index[6:0] ? _GEN_18465 : tag_1_59; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3786 = 7'h3c == index[6:0] ? _GEN_18465 : tag_1_60; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3787 = 7'h3d == index[6:0] ? _GEN_18465 : tag_1_61; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3788 = 7'h3e == index[6:0] ? _GEN_18465 : tag_1_62; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3789 = 7'h3f == index[6:0] ? _GEN_18465 : tag_1_63; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3790 = 7'h40 == index[6:0] ? _GEN_18465 : tag_1_64; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3791 = 7'h41 == index[6:0] ? _GEN_18465 : tag_1_65; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3792 = 7'h42 == index[6:0] ? _GEN_18465 : tag_1_66; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3793 = 7'h43 == index[6:0] ? _GEN_18465 : tag_1_67; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3794 = 7'h44 == index[6:0] ? _GEN_18465 : tag_1_68; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3795 = 7'h45 == index[6:0] ? _GEN_18465 : tag_1_69; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3796 = 7'h46 == index[6:0] ? _GEN_18465 : tag_1_70; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3797 = 7'h47 == index[6:0] ? _GEN_18465 : tag_1_71; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3798 = 7'h48 == index[6:0] ? _GEN_18465 : tag_1_72; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3799 = 7'h49 == index[6:0] ? _GEN_18465 : tag_1_73; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3800 = 7'h4a == index[6:0] ? _GEN_18465 : tag_1_74; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3801 = 7'h4b == index[6:0] ? _GEN_18465 : tag_1_75; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3802 = 7'h4c == index[6:0] ? _GEN_18465 : tag_1_76; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3803 = 7'h4d == index[6:0] ? _GEN_18465 : tag_1_77; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3804 = 7'h4e == index[6:0] ? _GEN_18465 : tag_1_78; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3805 = 7'h4f == index[6:0] ? _GEN_18465 : tag_1_79; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3806 = 7'h50 == index[6:0] ? _GEN_18465 : tag_1_80; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3807 = 7'h51 == index[6:0] ? _GEN_18465 : tag_1_81; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3808 = 7'h52 == index[6:0] ? _GEN_18465 : tag_1_82; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3809 = 7'h53 == index[6:0] ? _GEN_18465 : tag_1_83; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3810 = 7'h54 == index[6:0] ? _GEN_18465 : tag_1_84; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3811 = 7'h55 == index[6:0] ? _GEN_18465 : tag_1_85; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3812 = 7'h56 == index[6:0] ? _GEN_18465 : tag_1_86; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3813 = 7'h57 == index[6:0] ? _GEN_18465 : tag_1_87; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3814 = 7'h58 == index[6:0] ? _GEN_18465 : tag_1_88; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3815 = 7'h59 == index[6:0] ? _GEN_18465 : tag_1_89; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3816 = 7'h5a == index[6:0] ? _GEN_18465 : tag_1_90; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3817 = 7'h5b == index[6:0] ? _GEN_18465 : tag_1_91; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3818 = 7'h5c == index[6:0] ? _GEN_18465 : tag_1_92; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3819 = 7'h5d == index[6:0] ? _GEN_18465 : tag_1_93; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3820 = 7'h5e == index[6:0] ? _GEN_18465 : tag_1_94; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3821 = 7'h5f == index[6:0] ? _GEN_18465 : tag_1_95; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3822 = 7'h60 == index[6:0] ? _GEN_18465 : tag_1_96; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3823 = 7'h61 == index[6:0] ? _GEN_18465 : tag_1_97; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3824 = 7'h62 == index[6:0] ? _GEN_18465 : tag_1_98; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3825 = 7'h63 == index[6:0] ? _GEN_18465 : tag_1_99; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3826 = 7'h64 == index[6:0] ? _GEN_18465 : tag_1_100; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3827 = 7'h65 == index[6:0] ? _GEN_18465 : tag_1_101; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3828 = 7'h66 == index[6:0] ? _GEN_18465 : tag_1_102; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3829 = 7'h67 == index[6:0] ? _GEN_18465 : tag_1_103; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3830 = 7'h68 == index[6:0] ? _GEN_18465 : tag_1_104; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3831 = 7'h69 == index[6:0] ? _GEN_18465 : tag_1_105; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3832 = 7'h6a == index[6:0] ? _GEN_18465 : tag_1_106; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3833 = 7'h6b == index[6:0] ? _GEN_18465 : tag_1_107; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3834 = 7'h6c == index[6:0] ? _GEN_18465 : tag_1_108; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3835 = 7'h6d == index[6:0] ? _GEN_18465 : tag_1_109; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3836 = 7'h6e == index[6:0] ? _GEN_18465 : tag_1_110; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3837 = 7'h6f == index[6:0] ? _GEN_18465 : tag_1_111; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3838 = 7'h70 == index[6:0] ? _GEN_18465 : tag_1_112; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3839 = 7'h71 == index[6:0] ? _GEN_18465 : tag_1_113; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3840 = 7'h72 == index[6:0] ? _GEN_18465 : tag_1_114; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3841 = 7'h73 == index[6:0] ? _GEN_18465 : tag_1_115; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3842 = 7'h74 == index[6:0] ? _GEN_18465 : tag_1_116; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3843 = 7'h75 == index[6:0] ? _GEN_18465 : tag_1_117; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3844 = 7'h76 == index[6:0] ? _GEN_18465 : tag_1_118; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3845 = 7'h77 == index[6:0] ? _GEN_18465 : tag_1_119; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3846 = 7'h78 == index[6:0] ? _GEN_18465 : tag_1_120; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3847 = 7'h79 == index[6:0] ? _GEN_18465 : tag_1_121; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3848 = 7'h7a == index[6:0] ? _GEN_18465 : tag_1_122; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3849 = 7'h7b == index[6:0] ? _GEN_18465 : tag_1_123; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3850 = 7'h7c == index[6:0] ? _GEN_18465 : tag_1_124; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3851 = 7'h7d == index[6:0] ? _GEN_18465 : tag_1_125; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3852 = 7'h7e == index[6:0] ? _GEN_18465 : tag_1_126; // @[d_cache.scala 148:{30,30} 23:24]
  wire [31:0] _GEN_3853 = 7'h7f == index[6:0] ? _GEN_18465 : tag_1_127; // @[d_cache.scala 148:{30,30} 23:24]
  wire  _GEN_3854 = _GEN_18470 | valid_1_0; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3855 = _GEN_18471 | valid_1_1; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3856 = _GEN_18472 | valid_1_2; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3857 = _GEN_18473 | valid_1_3; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3858 = _GEN_18474 | valid_1_4; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3859 = _GEN_18475 | valid_1_5; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3860 = _GEN_18476 | valid_1_6; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3861 = _GEN_18477 | valid_1_7; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3862 = _GEN_18478 | valid_1_8; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3863 = _GEN_18479 | valid_1_9; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3864 = _GEN_18480 | valid_1_10; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3865 = _GEN_18481 | valid_1_11; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3866 = _GEN_18482 | valid_1_12; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3867 = _GEN_18483 | valid_1_13; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3868 = _GEN_18484 | valid_1_14; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3869 = _GEN_18485 | valid_1_15; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3870 = _GEN_18486 | valid_1_16; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3871 = _GEN_18487 | valid_1_17; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3872 = _GEN_18488 | valid_1_18; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3873 = _GEN_18489 | valid_1_19; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3874 = _GEN_18490 | valid_1_20; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3875 = _GEN_18491 | valid_1_21; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3876 = _GEN_18492 | valid_1_22; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3877 = _GEN_18493 | valid_1_23; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3878 = _GEN_18494 | valid_1_24; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3879 = _GEN_18495 | valid_1_25; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3880 = _GEN_18496 | valid_1_26; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3881 = _GEN_18497 | valid_1_27; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3882 = _GEN_18498 | valid_1_28; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3883 = _GEN_18499 | valid_1_29; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3884 = _GEN_18500 | valid_1_30; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3885 = _GEN_18501 | valid_1_31; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3886 = _GEN_18502 | valid_1_32; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3887 = _GEN_18503 | valid_1_33; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3888 = _GEN_18504 | valid_1_34; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3889 = _GEN_18505 | valid_1_35; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3890 = _GEN_18506 | valid_1_36; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3891 = _GEN_18507 | valid_1_37; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3892 = _GEN_18508 | valid_1_38; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3893 = _GEN_18509 | valid_1_39; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3894 = _GEN_18510 | valid_1_40; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3895 = _GEN_18511 | valid_1_41; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3896 = _GEN_18512 | valid_1_42; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3897 = _GEN_18513 | valid_1_43; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3898 = _GEN_18514 | valid_1_44; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3899 = _GEN_18515 | valid_1_45; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3900 = _GEN_18516 | valid_1_46; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3901 = _GEN_18517 | valid_1_47; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3902 = _GEN_18518 | valid_1_48; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3903 = _GEN_18519 | valid_1_49; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3904 = _GEN_18520 | valid_1_50; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3905 = _GEN_18521 | valid_1_51; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3906 = _GEN_18522 | valid_1_52; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3907 = _GEN_18523 | valid_1_53; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3908 = _GEN_18524 | valid_1_54; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3909 = _GEN_18525 | valid_1_55; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3910 = _GEN_18526 | valid_1_56; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3911 = _GEN_18527 | valid_1_57; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3912 = _GEN_18528 | valid_1_58; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3913 = _GEN_18529 | valid_1_59; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3914 = _GEN_18530 | valid_1_60; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3915 = _GEN_18531 | valid_1_61; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3916 = _GEN_18532 | valid_1_62; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3917 = _GEN_18533 | valid_1_63; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3918 = _GEN_18534 | valid_1_64; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3919 = _GEN_18535 | valid_1_65; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3920 = _GEN_18536 | valid_1_66; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3921 = _GEN_18537 | valid_1_67; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3922 = _GEN_18538 | valid_1_68; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3923 = _GEN_18539 | valid_1_69; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3924 = _GEN_18540 | valid_1_70; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3925 = _GEN_18541 | valid_1_71; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3926 = _GEN_18542 | valid_1_72; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3927 = _GEN_18543 | valid_1_73; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3928 = _GEN_18544 | valid_1_74; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3929 = _GEN_18545 | valid_1_75; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3930 = _GEN_18546 | valid_1_76; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3931 = _GEN_18547 | valid_1_77; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3932 = _GEN_18548 | valid_1_78; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3933 = _GEN_18549 | valid_1_79; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3934 = _GEN_18550 | valid_1_80; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3935 = _GEN_18551 | valid_1_81; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3936 = _GEN_18552 | valid_1_82; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3937 = _GEN_18553 | valid_1_83; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3938 = _GEN_18554 | valid_1_84; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3939 = _GEN_18555 | valid_1_85; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3940 = _GEN_18556 | valid_1_86; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3941 = _GEN_18557 | valid_1_87; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3942 = _GEN_18558 | valid_1_88; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3943 = _GEN_18559 | valid_1_89; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3944 = _GEN_18560 | valid_1_90; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3945 = _GEN_18561 | valid_1_91; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3946 = _GEN_18562 | valid_1_92; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3947 = _GEN_18563 | valid_1_93; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3948 = _GEN_18564 | valid_1_94; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3949 = _GEN_18565 | valid_1_95; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3950 = _GEN_18566 | valid_1_96; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3951 = _GEN_18567 | valid_1_97; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3952 = _GEN_18568 | valid_1_98; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3953 = _GEN_18569 | valid_1_99; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3954 = _GEN_18570 | valid_1_100; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3955 = _GEN_18571 | valid_1_101; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3956 = _GEN_18572 | valid_1_102; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3957 = _GEN_18573 | valid_1_103; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3958 = _GEN_18574 | valid_1_104; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3959 = _GEN_18575 | valid_1_105; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3960 = _GEN_18576 | valid_1_106; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3961 = _GEN_18577 | valid_1_107; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3962 = _GEN_18578 | valid_1_108; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3963 = _GEN_18579 | valid_1_109; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3964 = _GEN_18580 | valid_1_110; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3965 = _GEN_18581 | valid_1_111; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3966 = _GEN_18582 | valid_1_112; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3967 = _GEN_18583 | valid_1_113; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3968 = _GEN_18584 | valid_1_114; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3969 = _GEN_18585 | valid_1_115; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3970 = _GEN_18586 | valid_1_116; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3971 = _GEN_18587 | valid_1_117; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3972 = _GEN_18588 | valid_1_118; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3973 = _GEN_18589 | valid_1_119; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3974 = _GEN_18590 | valid_1_120; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3975 = _GEN_18591 | valid_1_121; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3976 = _GEN_18592 | valid_1_122; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3977 = _GEN_18593 | valid_1_123; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3978 = _GEN_18594 | valid_1_124; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3979 = _GEN_18595 | valid_1_125; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3980 = _GEN_18596 | valid_1_126; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _GEN_3981 = _GEN_18597 | valid_1_127; // @[d_cache.scala 149:{32,32} 25:26]
  wire  _T_46 = ~quene; // @[d_cache.scala 152:27]
  wire [41:0] _write_back_addr_T_1 = {_GEN_127, 10'h0}; // @[d_cache.scala 156:58]
  wire [34:0] _write_back_addr_T_2 = {index, 3'h0}; // @[d_cache.scala 156:74]
  wire [41:0] _GEN_18985 = {{7'd0}, _write_back_addr_T_2}; // @[d_cache.scala 156:65]
  wire [41:0] _write_back_addr_T_3 = _write_back_addr_T_1 | _GEN_18985; // @[d_cache.scala 156:65]
  wire  _GEN_4622 = 7'h0 == index[6:0] ? 1'h0 : dirty_0_0; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4623 = 7'h1 == index[6:0] ? 1'h0 : dirty_0_1; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4624 = 7'h2 == index[6:0] ? 1'h0 : dirty_0_2; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4625 = 7'h3 == index[6:0] ? 1'h0 : dirty_0_3; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4626 = 7'h4 == index[6:0] ? 1'h0 : dirty_0_4; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4627 = 7'h5 == index[6:0] ? 1'h0 : dirty_0_5; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4628 = 7'h6 == index[6:0] ? 1'h0 : dirty_0_6; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4629 = 7'h7 == index[6:0] ? 1'h0 : dirty_0_7; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4630 = 7'h8 == index[6:0] ? 1'h0 : dirty_0_8; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4631 = 7'h9 == index[6:0] ? 1'h0 : dirty_0_9; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4632 = 7'ha == index[6:0] ? 1'h0 : dirty_0_10; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4633 = 7'hb == index[6:0] ? 1'h0 : dirty_0_11; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4634 = 7'hc == index[6:0] ? 1'h0 : dirty_0_12; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4635 = 7'hd == index[6:0] ? 1'h0 : dirty_0_13; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4636 = 7'he == index[6:0] ? 1'h0 : dirty_0_14; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4637 = 7'hf == index[6:0] ? 1'h0 : dirty_0_15; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4638 = 7'h10 == index[6:0] ? 1'h0 : dirty_0_16; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4639 = 7'h11 == index[6:0] ? 1'h0 : dirty_0_17; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4640 = 7'h12 == index[6:0] ? 1'h0 : dirty_0_18; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4641 = 7'h13 == index[6:0] ? 1'h0 : dirty_0_19; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4642 = 7'h14 == index[6:0] ? 1'h0 : dirty_0_20; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4643 = 7'h15 == index[6:0] ? 1'h0 : dirty_0_21; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4644 = 7'h16 == index[6:0] ? 1'h0 : dirty_0_22; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4645 = 7'h17 == index[6:0] ? 1'h0 : dirty_0_23; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4646 = 7'h18 == index[6:0] ? 1'h0 : dirty_0_24; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4647 = 7'h19 == index[6:0] ? 1'h0 : dirty_0_25; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4648 = 7'h1a == index[6:0] ? 1'h0 : dirty_0_26; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4649 = 7'h1b == index[6:0] ? 1'h0 : dirty_0_27; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4650 = 7'h1c == index[6:0] ? 1'h0 : dirty_0_28; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4651 = 7'h1d == index[6:0] ? 1'h0 : dirty_0_29; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4652 = 7'h1e == index[6:0] ? 1'h0 : dirty_0_30; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4653 = 7'h1f == index[6:0] ? 1'h0 : dirty_0_31; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4654 = 7'h20 == index[6:0] ? 1'h0 : dirty_0_32; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4655 = 7'h21 == index[6:0] ? 1'h0 : dirty_0_33; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4656 = 7'h22 == index[6:0] ? 1'h0 : dirty_0_34; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4657 = 7'h23 == index[6:0] ? 1'h0 : dirty_0_35; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4658 = 7'h24 == index[6:0] ? 1'h0 : dirty_0_36; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4659 = 7'h25 == index[6:0] ? 1'h0 : dirty_0_37; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4660 = 7'h26 == index[6:0] ? 1'h0 : dirty_0_38; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4661 = 7'h27 == index[6:0] ? 1'h0 : dirty_0_39; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4662 = 7'h28 == index[6:0] ? 1'h0 : dirty_0_40; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4663 = 7'h29 == index[6:0] ? 1'h0 : dirty_0_41; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4664 = 7'h2a == index[6:0] ? 1'h0 : dirty_0_42; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4665 = 7'h2b == index[6:0] ? 1'h0 : dirty_0_43; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4666 = 7'h2c == index[6:0] ? 1'h0 : dirty_0_44; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4667 = 7'h2d == index[6:0] ? 1'h0 : dirty_0_45; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4668 = 7'h2e == index[6:0] ? 1'h0 : dirty_0_46; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4669 = 7'h2f == index[6:0] ? 1'h0 : dirty_0_47; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4670 = 7'h30 == index[6:0] ? 1'h0 : dirty_0_48; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4671 = 7'h31 == index[6:0] ? 1'h0 : dirty_0_49; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4672 = 7'h32 == index[6:0] ? 1'h0 : dirty_0_50; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4673 = 7'h33 == index[6:0] ? 1'h0 : dirty_0_51; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4674 = 7'h34 == index[6:0] ? 1'h0 : dirty_0_52; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4675 = 7'h35 == index[6:0] ? 1'h0 : dirty_0_53; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4676 = 7'h36 == index[6:0] ? 1'h0 : dirty_0_54; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4677 = 7'h37 == index[6:0] ? 1'h0 : dirty_0_55; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4678 = 7'h38 == index[6:0] ? 1'h0 : dirty_0_56; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4679 = 7'h39 == index[6:0] ? 1'h0 : dirty_0_57; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4680 = 7'h3a == index[6:0] ? 1'h0 : dirty_0_58; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4681 = 7'h3b == index[6:0] ? 1'h0 : dirty_0_59; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4682 = 7'h3c == index[6:0] ? 1'h0 : dirty_0_60; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4683 = 7'h3d == index[6:0] ? 1'h0 : dirty_0_61; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4684 = 7'h3e == index[6:0] ? 1'h0 : dirty_0_62; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4685 = 7'h3f == index[6:0] ? 1'h0 : dirty_0_63; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4686 = 7'h40 == index[6:0] ? 1'h0 : dirty_0_64; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4687 = 7'h41 == index[6:0] ? 1'h0 : dirty_0_65; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4688 = 7'h42 == index[6:0] ? 1'h0 : dirty_0_66; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4689 = 7'h43 == index[6:0] ? 1'h0 : dirty_0_67; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4690 = 7'h44 == index[6:0] ? 1'h0 : dirty_0_68; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4691 = 7'h45 == index[6:0] ? 1'h0 : dirty_0_69; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4692 = 7'h46 == index[6:0] ? 1'h0 : dirty_0_70; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4693 = 7'h47 == index[6:0] ? 1'h0 : dirty_0_71; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4694 = 7'h48 == index[6:0] ? 1'h0 : dirty_0_72; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4695 = 7'h49 == index[6:0] ? 1'h0 : dirty_0_73; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4696 = 7'h4a == index[6:0] ? 1'h0 : dirty_0_74; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4697 = 7'h4b == index[6:0] ? 1'h0 : dirty_0_75; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4698 = 7'h4c == index[6:0] ? 1'h0 : dirty_0_76; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4699 = 7'h4d == index[6:0] ? 1'h0 : dirty_0_77; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4700 = 7'h4e == index[6:0] ? 1'h0 : dirty_0_78; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4701 = 7'h4f == index[6:0] ? 1'h0 : dirty_0_79; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4702 = 7'h50 == index[6:0] ? 1'h0 : dirty_0_80; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4703 = 7'h51 == index[6:0] ? 1'h0 : dirty_0_81; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4704 = 7'h52 == index[6:0] ? 1'h0 : dirty_0_82; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4705 = 7'h53 == index[6:0] ? 1'h0 : dirty_0_83; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4706 = 7'h54 == index[6:0] ? 1'h0 : dirty_0_84; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4707 = 7'h55 == index[6:0] ? 1'h0 : dirty_0_85; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4708 = 7'h56 == index[6:0] ? 1'h0 : dirty_0_86; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4709 = 7'h57 == index[6:0] ? 1'h0 : dirty_0_87; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4710 = 7'h58 == index[6:0] ? 1'h0 : dirty_0_88; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4711 = 7'h59 == index[6:0] ? 1'h0 : dirty_0_89; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4712 = 7'h5a == index[6:0] ? 1'h0 : dirty_0_90; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4713 = 7'h5b == index[6:0] ? 1'h0 : dirty_0_91; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4714 = 7'h5c == index[6:0] ? 1'h0 : dirty_0_92; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4715 = 7'h5d == index[6:0] ? 1'h0 : dirty_0_93; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4716 = 7'h5e == index[6:0] ? 1'h0 : dirty_0_94; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4717 = 7'h5f == index[6:0] ? 1'h0 : dirty_0_95; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4718 = 7'h60 == index[6:0] ? 1'h0 : dirty_0_96; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4719 = 7'h61 == index[6:0] ? 1'h0 : dirty_0_97; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4720 = 7'h62 == index[6:0] ? 1'h0 : dirty_0_98; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4721 = 7'h63 == index[6:0] ? 1'h0 : dirty_0_99; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4722 = 7'h64 == index[6:0] ? 1'h0 : dirty_0_100; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4723 = 7'h65 == index[6:0] ? 1'h0 : dirty_0_101; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4724 = 7'h66 == index[6:0] ? 1'h0 : dirty_0_102; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4725 = 7'h67 == index[6:0] ? 1'h0 : dirty_0_103; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4726 = 7'h68 == index[6:0] ? 1'h0 : dirty_0_104; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4727 = 7'h69 == index[6:0] ? 1'h0 : dirty_0_105; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4728 = 7'h6a == index[6:0] ? 1'h0 : dirty_0_106; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4729 = 7'h6b == index[6:0] ? 1'h0 : dirty_0_107; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4730 = 7'h6c == index[6:0] ? 1'h0 : dirty_0_108; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4731 = 7'h6d == index[6:0] ? 1'h0 : dirty_0_109; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4732 = 7'h6e == index[6:0] ? 1'h0 : dirty_0_110; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4733 = 7'h6f == index[6:0] ? 1'h0 : dirty_0_111; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4734 = 7'h70 == index[6:0] ? 1'h0 : dirty_0_112; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4735 = 7'h71 == index[6:0] ? 1'h0 : dirty_0_113; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4736 = 7'h72 == index[6:0] ? 1'h0 : dirty_0_114; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4737 = 7'h73 == index[6:0] ? 1'h0 : dirty_0_115; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4738 = 7'h74 == index[6:0] ? 1'h0 : dirty_0_116; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4739 = 7'h75 == index[6:0] ? 1'h0 : dirty_0_117; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4740 = 7'h76 == index[6:0] ? 1'h0 : dirty_0_118; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4741 = 7'h77 == index[6:0] ? 1'h0 : dirty_0_119; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4742 = 7'h78 == index[6:0] ? 1'h0 : dirty_0_120; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4743 = 7'h79 == index[6:0] ? 1'h0 : dirty_0_121; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4744 = 7'h7a == index[6:0] ? 1'h0 : dirty_0_122; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4745 = 7'h7b == index[6:0] ? 1'h0 : dirty_0_123; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4746 = 7'h7c == index[6:0] ? 1'h0 : dirty_0_124; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4747 = 7'h7d == index[6:0] ? 1'h0 : dirty_0_125; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4748 = 7'h7e == index[6:0] ? 1'h0 : dirty_0_126; // @[d_cache.scala 159:{40,40} 26:26]
  wire  _GEN_4749 = 7'h7f == index[6:0] ? 1'h0 : dirty_0_127; // @[d_cache.scala 159:{40,40} 26:26]
  wire [63:0] _GEN_5262 = _GEN_901 ? _GEN_1160 : write_back_data; // @[d_cache.scala 154:47 155:41 31:34]
  wire [41:0] _GEN_5263 = _GEN_901 ? _write_back_addr_T_3 : {{10'd0}, write_back_addr}; // @[d_cache.scala 154:47 156:41 32:34]
  wire [63:0] _GEN_5264 = _GEN_901 ? _GEN_3214 : _GEN_3214; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5265 = _GEN_901 ? _GEN_3215 : _GEN_3215; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5266 = _GEN_901 ? _GEN_3216 : _GEN_3216; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5267 = _GEN_901 ? _GEN_3217 : _GEN_3217; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5268 = _GEN_901 ? _GEN_3218 : _GEN_3218; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5269 = _GEN_901 ? _GEN_3219 : _GEN_3219; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5270 = _GEN_901 ? _GEN_3220 : _GEN_3220; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5271 = _GEN_901 ? _GEN_3221 : _GEN_3221; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5272 = _GEN_901 ? _GEN_3222 : _GEN_3222; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5273 = _GEN_901 ? _GEN_3223 : _GEN_3223; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5274 = _GEN_901 ? _GEN_3224 : _GEN_3224; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5275 = _GEN_901 ? _GEN_3225 : _GEN_3225; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5276 = _GEN_901 ? _GEN_3226 : _GEN_3226; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5277 = _GEN_901 ? _GEN_3227 : _GEN_3227; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5278 = _GEN_901 ? _GEN_3228 : _GEN_3228; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5279 = _GEN_901 ? _GEN_3229 : _GEN_3229; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5280 = _GEN_901 ? _GEN_3230 : _GEN_3230; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5281 = _GEN_901 ? _GEN_3231 : _GEN_3231; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5282 = _GEN_901 ? _GEN_3232 : _GEN_3232; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5283 = _GEN_901 ? _GEN_3233 : _GEN_3233; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5284 = _GEN_901 ? _GEN_3234 : _GEN_3234; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5285 = _GEN_901 ? _GEN_3235 : _GEN_3235; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5286 = _GEN_901 ? _GEN_3236 : _GEN_3236; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5287 = _GEN_901 ? _GEN_3237 : _GEN_3237; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5288 = _GEN_901 ? _GEN_3238 : _GEN_3238; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5289 = _GEN_901 ? _GEN_3239 : _GEN_3239; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5290 = _GEN_901 ? _GEN_3240 : _GEN_3240; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5291 = _GEN_901 ? _GEN_3241 : _GEN_3241; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5292 = _GEN_901 ? _GEN_3242 : _GEN_3242; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5293 = _GEN_901 ? _GEN_3243 : _GEN_3243; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5294 = _GEN_901 ? _GEN_3244 : _GEN_3244; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5295 = _GEN_901 ? _GEN_3245 : _GEN_3245; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5296 = _GEN_901 ? _GEN_3246 : _GEN_3246; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5297 = _GEN_901 ? _GEN_3247 : _GEN_3247; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5298 = _GEN_901 ? _GEN_3248 : _GEN_3248; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5299 = _GEN_901 ? _GEN_3249 : _GEN_3249; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5300 = _GEN_901 ? _GEN_3250 : _GEN_3250; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5301 = _GEN_901 ? _GEN_3251 : _GEN_3251; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5302 = _GEN_901 ? _GEN_3252 : _GEN_3252; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5303 = _GEN_901 ? _GEN_3253 : _GEN_3253; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5304 = _GEN_901 ? _GEN_3254 : _GEN_3254; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5305 = _GEN_901 ? _GEN_3255 : _GEN_3255; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5306 = _GEN_901 ? _GEN_3256 : _GEN_3256; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5307 = _GEN_901 ? _GEN_3257 : _GEN_3257; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5308 = _GEN_901 ? _GEN_3258 : _GEN_3258; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5309 = _GEN_901 ? _GEN_3259 : _GEN_3259; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5310 = _GEN_901 ? _GEN_3260 : _GEN_3260; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5311 = _GEN_901 ? _GEN_3261 : _GEN_3261; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5312 = _GEN_901 ? _GEN_3262 : _GEN_3262; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5313 = _GEN_901 ? _GEN_3263 : _GEN_3263; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5314 = _GEN_901 ? _GEN_3264 : _GEN_3264; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5315 = _GEN_901 ? _GEN_3265 : _GEN_3265; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5316 = _GEN_901 ? _GEN_3266 : _GEN_3266; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5317 = _GEN_901 ? _GEN_3267 : _GEN_3267; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5318 = _GEN_901 ? _GEN_3268 : _GEN_3268; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5319 = _GEN_901 ? _GEN_3269 : _GEN_3269; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5320 = _GEN_901 ? _GEN_3270 : _GEN_3270; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5321 = _GEN_901 ? _GEN_3271 : _GEN_3271; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5322 = _GEN_901 ? _GEN_3272 : _GEN_3272; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5323 = _GEN_901 ? _GEN_3273 : _GEN_3273; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5324 = _GEN_901 ? _GEN_3274 : _GEN_3274; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5325 = _GEN_901 ? _GEN_3275 : _GEN_3275; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5326 = _GEN_901 ? _GEN_3276 : _GEN_3276; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5327 = _GEN_901 ? _GEN_3277 : _GEN_3277; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5328 = _GEN_901 ? _GEN_3278 : _GEN_3278; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5329 = _GEN_901 ? _GEN_3279 : _GEN_3279; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5330 = _GEN_901 ? _GEN_3280 : _GEN_3280; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5331 = _GEN_901 ? _GEN_3281 : _GEN_3281; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5332 = _GEN_901 ? _GEN_3282 : _GEN_3282; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5333 = _GEN_901 ? _GEN_3283 : _GEN_3283; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5334 = _GEN_901 ? _GEN_3284 : _GEN_3284; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5335 = _GEN_901 ? _GEN_3285 : _GEN_3285; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5336 = _GEN_901 ? _GEN_3286 : _GEN_3286; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5337 = _GEN_901 ? _GEN_3287 : _GEN_3287; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5338 = _GEN_901 ? _GEN_3288 : _GEN_3288; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5339 = _GEN_901 ? _GEN_3289 : _GEN_3289; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5340 = _GEN_901 ? _GEN_3290 : _GEN_3290; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5341 = _GEN_901 ? _GEN_3291 : _GEN_3291; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5342 = _GEN_901 ? _GEN_3292 : _GEN_3292; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5343 = _GEN_901 ? _GEN_3293 : _GEN_3293; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5344 = _GEN_901 ? _GEN_3294 : _GEN_3294; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5345 = _GEN_901 ? _GEN_3295 : _GEN_3295; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5346 = _GEN_901 ? _GEN_3296 : _GEN_3296; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5347 = _GEN_901 ? _GEN_3297 : _GEN_3297; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5348 = _GEN_901 ? _GEN_3298 : _GEN_3298; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5349 = _GEN_901 ? _GEN_3299 : _GEN_3299; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5350 = _GEN_901 ? _GEN_3300 : _GEN_3300; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5351 = _GEN_901 ? _GEN_3301 : _GEN_3301; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5352 = _GEN_901 ? _GEN_3302 : _GEN_3302; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5353 = _GEN_901 ? _GEN_3303 : _GEN_3303; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5354 = _GEN_901 ? _GEN_3304 : _GEN_3304; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5355 = _GEN_901 ? _GEN_3305 : _GEN_3305; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5356 = _GEN_901 ? _GEN_3306 : _GEN_3306; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5357 = _GEN_901 ? _GEN_3307 : _GEN_3307; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5358 = _GEN_901 ? _GEN_3308 : _GEN_3308; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5359 = _GEN_901 ? _GEN_3309 : _GEN_3309; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5360 = _GEN_901 ? _GEN_3310 : _GEN_3310; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5361 = _GEN_901 ? _GEN_3311 : _GEN_3311; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5362 = _GEN_901 ? _GEN_3312 : _GEN_3312; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5363 = _GEN_901 ? _GEN_3313 : _GEN_3313; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5364 = _GEN_901 ? _GEN_3314 : _GEN_3314; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5365 = _GEN_901 ? _GEN_3315 : _GEN_3315; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5366 = _GEN_901 ? _GEN_3316 : _GEN_3316; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5367 = _GEN_901 ? _GEN_3317 : _GEN_3317; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5368 = _GEN_901 ? _GEN_3318 : _GEN_3318; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5369 = _GEN_901 ? _GEN_3319 : _GEN_3319; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5370 = _GEN_901 ? _GEN_3320 : _GEN_3320; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5371 = _GEN_901 ? _GEN_3321 : _GEN_3321; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5372 = _GEN_901 ? _GEN_3322 : _GEN_3322; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5373 = _GEN_901 ? _GEN_3323 : _GEN_3323; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5374 = _GEN_901 ? _GEN_3324 : _GEN_3324; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5375 = _GEN_901 ? _GEN_3325 : _GEN_3325; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5376 = _GEN_901 ? _GEN_3326 : _GEN_3326; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5377 = _GEN_901 ? _GEN_3327 : _GEN_3327; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5378 = _GEN_901 ? _GEN_3328 : _GEN_3328; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5379 = _GEN_901 ? _GEN_3329 : _GEN_3329; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5380 = _GEN_901 ? _GEN_3330 : _GEN_3330; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5381 = _GEN_901 ? _GEN_3331 : _GEN_3331; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5382 = _GEN_901 ? _GEN_3332 : _GEN_3332; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5383 = _GEN_901 ? _GEN_3333 : _GEN_3333; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5384 = _GEN_901 ? _GEN_3334 : _GEN_3334; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5385 = _GEN_901 ? _GEN_3335 : _GEN_3335; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5386 = _GEN_901 ? _GEN_3336 : _GEN_3336; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5387 = _GEN_901 ? _GEN_3337 : _GEN_3337; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5388 = _GEN_901 ? _GEN_3338 : _GEN_3338; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5389 = _GEN_901 ? _GEN_3339 : _GEN_3339; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5390 = _GEN_901 ? _GEN_3340 : _GEN_3340; // @[d_cache.scala 154:47]
  wire [63:0] _GEN_5391 = _GEN_901 ? _GEN_3341 : _GEN_3341; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5392 = _GEN_901 ? _GEN_3342 : _GEN_3342; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5393 = _GEN_901 ? _GEN_3343 : _GEN_3343; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5394 = _GEN_901 ? _GEN_3344 : _GEN_3344; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5395 = _GEN_901 ? _GEN_3345 : _GEN_3345; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5396 = _GEN_901 ? _GEN_3346 : _GEN_3346; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5397 = _GEN_901 ? _GEN_3347 : _GEN_3347; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5398 = _GEN_901 ? _GEN_3348 : _GEN_3348; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5399 = _GEN_901 ? _GEN_3349 : _GEN_3349; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5400 = _GEN_901 ? _GEN_3350 : _GEN_3350; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5401 = _GEN_901 ? _GEN_3351 : _GEN_3351; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5402 = _GEN_901 ? _GEN_3352 : _GEN_3352; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5403 = _GEN_901 ? _GEN_3353 : _GEN_3353; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5404 = _GEN_901 ? _GEN_3354 : _GEN_3354; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5405 = _GEN_901 ? _GEN_3355 : _GEN_3355; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5406 = _GEN_901 ? _GEN_3356 : _GEN_3356; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5407 = _GEN_901 ? _GEN_3357 : _GEN_3357; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5408 = _GEN_901 ? _GEN_3358 : _GEN_3358; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5409 = _GEN_901 ? _GEN_3359 : _GEN_3359; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5410 = _GEN_901 ? _GEN_3360 : _GEN_3360; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5411 = _GEN_901 ? _GEN_3361 : _GEN_3361; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5412 = _GEN_901 ? _GEN_3362 : _GEN_3362; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5413 = _GEN_901 ? _GEN_3363 : _GEN_3363; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5414 = _GEN_901 ? _GEN_3364 : _GEN_3364; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5415 = _GEN_901 ? _GEN_3365 : _GEN_3365; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5416 = _GEN_901 ? _GEN_3366 : _GEN_3366; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5417 = _GEN_901 ? _GEN_3367 : _GEN_3367; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5418 = _GEN_901 ? _GEN_3368 : _GEN_3368; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5419 = _GEN_901 ? _GEN_3369 : _GEN_3369; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5420 = _GEN_901 ? _GEN_3370 : _GEN_3370; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5421 = _GEN_901 ? _GEN_3371 : _GEN_3371; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5422 = _GEN_901 ? _GEN_3372 : _GEN_3372; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5423 = _GEN_901 ? _GEN_3373 : _GEN_3373; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5424 = _GEN_901 ? _GEN_3374 : _GEN_3374; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5425 = _GEN_901 ? _GEN_3375 : _GEN_3375; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5426 = _GEN_901 ? _GEN_3376 : _GEN_3376; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5427 = _GEN_901 ? _GEN_3377 : _GEN_3377; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5428 = _GEN_901 ? _GEN_3378 : _GEN_3378; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5429 = _GEN_901 ? _GEN_3379 : _GEN_3379; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5430 = _GEN_901 ? _GEN_3380 : _GEN_3380; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5431 = _GEN_901 ? _GEN_3381 : _GEN_3381; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5432 = _GEN_901 ? _GEN_3382 : _GEN_3382; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5433 = _GEN_901 ? _GEN_3383 : _GEN_3383; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5434 = _GEN_901 ? _GEN_3384 : _GEN_3384; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5435 = _GEN_901 ? _GEN_3385 : _GEN_3385; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5436 = _GEN_901 ? _GEN_3386 : _GEN_3386; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5437 = _GEN_901 ? _GEN_3387 : _GEN_3387; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5438 = _GEN_901 ? _GEN_3388 : _GEN_3388; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5439 = _GEN_901 ? _GEN_3389 : _GEN_3389; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5440 = _GEN_901 ? _GEN_3390 : _GEN_3390; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5441 = _GEN_901 ? _GEN_3391 : _GEN_3391; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5442 = _GEN_901 ? _GEN_3392 : _GEN_3392; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5443 = _GEN_901 ? _GEN_3393 : _GEN_3393; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5444 = _GEN_901 ? _GEN_3394 : _GEN_3394; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5445 = _GEN_901 ? _GEN_3395 : _GEN_3395; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5446 = _GEN_901 ? _GEN_3396 : _GEN_3396; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5447 = _GEN_901 ? _GEN_3397 : _GEN_3397; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5448 = _GEN_901 ? _GEN_3398 : _GEN_3398; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5449 = _GEN_901 ? _GEN_3399 : _GEN_3399; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5450 = _GEN_901 ? _GEN_3400 : _GEN_3400; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5451 = _GEN_901 ? _GEN_3401 : _GEN_3401; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5452 = _GEN_901 ? _GEN_3402 : _GEN_3402; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5453 = _GEN_901 ? _GEN_3403 : _GEN_3403; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5454 = _GEN_901 ? _GEN_3404 : _GEN_3404; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5455 = _GEN_901 ? _GEN_3405 : _GEN_3405; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5456 = _GEN_901 ? _GEN_3406 : _GEN_3406; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5457 = _GEN_901 ? _GEN_3407 : _GEN_3407; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5458 = _GEN_901 ? _GEN_3408 : _GEN_3408; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5459 = _GEN_901 ? _GEN_3409 : _GEN_3409; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5460 = _GEN_901 ? _GEN_3410 : _GEN_3410; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5461 = _GEN_901 ? _GEN_3411 : _GEN_3411; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5462 = _GEN_901 ? _GEN_3412 : _GEN_3412; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5463 = _GEN_901 ? _GEN_3413 : _GEN_3413; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5464 = _GEN_901 ? _GEN_3414 : _GEN_3414; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5465 = _GEN_901 ? _GEN_3415 : _GEN_3415; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5466 = _GEN_901 ? _GEN_3416 : _GEN_3416; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5467 = _GEN_901 ? _GEN_3417 : _GEN_3417; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5468 = _GEN_901 ? _GEN_3418 : _GEN_3418; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5469 = _GEN_901 ? _GEN_3419 : _GEN_3419; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5470 = _GEN_901 ? _GEN_3420 : _GEN_3420; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5471 = _GEN_901 ? _GEN_3421 : _GEN_3421; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5472 = _GEN_901 ? _GEN_3422 : _GEN_3422; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5473 = _GEN_901 ? _GEN_3423 : _GEN_3423; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5474 = _GEN_901 ? _GEN_3424 : _GEN_3424; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5475 = _GEN_901 ? _GEN_3425 : _GEN_3425; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5476 = _GEN_901 ? _GEN_3426 : _GEN_3426; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5477 = _GEN_901 ? _GEN_3427 : _GEN_3427; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5478 = _GEN_901 ? _GEN_3428 : _GEN_3428; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5479 = _GEN_901 ? _GEN_3429 : _GEN_3429; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5480 = _GEN_901 ? _GEN_3430 : _GEN_3430; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5481 = _GEN_901 ? _GEN_3431 : _GEN_3431; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5482 = _GEN_901 ? _GEN_3432 : _GEN_3432; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5483 = _GEN_901 ? _GEN_3433 : _GEN_3433; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5484 = _GEN_901 ? _GEN_3434 : _GEN_3434; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5485 = _GEN_901 ? _GEN_3435 : _GEN_3435; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5486 = _GEN_901 ? _GEN_3436 : _GEN_3436; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5487 = _GEN_901 ? _GEN_3437 : _GEN_3437; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5488 = _GEN_901 ? _GEN_3438 : _GEN_3438; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5489 = _GEN_901 ? _GEN_3439 : _GEN_3439; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5490 = _GEN_901 ? _GEN_3440 : _GEN_3440; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5491 = _GEN_901 ? _GEN_3441 : _GEN_3441; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5492 = _GEN_901 ? _GEN_3442 : _GEN_3442; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5493 = _GEN_901 ? _GEN_3443 : _GEN_3443; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5494 = _GEN_901 ? _GEN_3444 : _GEN_3444; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5495 = _GEN_901 ? _GEN_3445 : _GEN_3445; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5496 = _GEN_901 ? _GEN_3446 : _GEN_3446; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5497 = _GEN_901 ? _GEN_3447 : _GEN_3447; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5498 = _GEN_901 ? _GEN_3448 : _GEN_3448; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5499 = _GEN_901 ? _GEN_3449 : _GEN_3449; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5500 = _GEN_901 ? _GEN_3450 : _GEN_3450; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5501 = _GEN_901 ? _GEN_3451 : _GEN_3451; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5502 = _GEN_901 ? _GEN_3452 : _GEN_3452; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5503 = _GEN_901 ? _GEN_3453 : _GEN_3453; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5504 = _GEN_901 ? _GEN_3454 : _GEN_3454; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5505 = _GEN_901 ? _GEN_3455 : _GEN_3455; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5506 = _GEN_901 ? _GEN_3456 : _GEN_3456; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5507 = _GEN_901 ? _GEN_3457 : _GEN_3457; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5508 = _GEN_901 ? _GEN_3458 : _GEN_3458; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5509 = _GEN_901 ? _GEN_3459 : _GEN_3459; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5510 = _GEN_901 ? _GEN_3460 : _GEN_3460; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5511 = _GEN_901 ? _GEN_3461 : _GEN_3461; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5512 = _GEN_901 ? _GEN_3462 : _GEN_3462; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5513 = _GEN_901 ? _GEN_3463 : _GEN_3463; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5514 = _GEN_901 ? _GEN_3464 : _GEN_3464; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5515 = _GEN_901 ? _GEN_3465 : _GEN_3465; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5516 = _GEN_901 ? _GEN_3466 : _GEN_3466; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5517 = _GEN_901 ? _GEN_3467 : _GEN_3467; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5518 = _GEN_901 ? _GEN_3468 : _GEN_3468; // @[d_cache.scala 154:47]
  wire [31:0] _GEN_5519 = _GEN_901 ? _GEN_3469 : _GEN_3469; // @[d_cache.scala 154:47]
  wire  _GEN_5520 = _GEN_901 ? _GEN_4622 : dirty_0_0; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5521 = _GEN_901 ? _GEN_4623 : dirty_0_1; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5522 = _GEN_901 ? _GEN_4624 : dirty_0_2; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5523 = _GEN_901 ? _GEN_4625 : dirty_0_3; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5524 = _GEN_901 ? _GEN_4626 : dirty_0_4; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5525 = _GEN_901 ? _GEN_4627 : dirty_0_5; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5526 = _GEN_901 ? _GEN_4628 : dirty_0_6; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5527 = _GEN_901 ? _GEN_4629 : dirty_0_7; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5528 = _GEN_901 ? _GEN_4630 : dirty_0_8; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5529 = _GEN_901 ? _GEN_4631 : dirty_0_9; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5530 = _GEN_901 ? _GEN_4632 : dirty_0_10; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5531 = _GEN_901 ? _GEN_4633 : dirty_0_11; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5532 = _GEN_901 ? _GEN_4634 : dirty_0_12; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5533 = _GEN_901 ? _GEN_4635 : dirty_0_13; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5534 = _GEN_901 ? _GEN_4636 : dirty_0_14; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5535 = _GEN_901 ? _GEN_4637 : dirty_0_15; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5536 = _GEN_901 ? _GEN_4638 : dirty_0_16; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5537 = _GEN_901 ? _GEN_4639 : dirty_0_17; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5538 = _GEN_901 ? _GEN_4640 : dirty_0_18; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5539 = _GEN_901 ? _GEN_4641 : dirty_0_19; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5540 = _GEN_901 ? _GEN_4642 : dirty_0_20; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5541 = _GEN_901 ? _GEN_4643 : dirty_0_21; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5542 = _GEN_901 ? _GEN_4644 : dirty_0_22; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5543 = _GEN_901 ? _GEN_4645 : dirty_0_23; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5544 = _GEN_901 ? _GEN_4646 : dirty_0_24; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5545 = _GEN_901 ? _GEN_4647 : dirty_0_25; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5546 = _GEN_901 ? _GEN_4648 : dirty_0_26; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5547 = _GEN_901 ? _GEN_4649 : dirty_0_27; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5548 = _GEN_901 ? _GEN_4650 : dirty_0_28; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5549 = _GEN_901 ? _GEN_4651 : dirty_0_29; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5550 = _GEN_901 ? _GEN_4652 : dirty_0_30; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5551 = _GEN_901 ? _GEN_4653 : dirty_0_31; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5552 = _GEN_901 ? _GEN_4654 : dirty_0_32; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5553 = _GEN_901 ? _GEN_4655 : dirty_0_33; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5554 = _GEN_901 ? _GEN_4656 : dirty_0_34; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5555 = _GEN_901 ? _GEN_4657 : dirty_0_35; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5556 = _GEN_901 ? _GEN_4658 : dirty_0_36; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5557 = _GEN_901 ? _GEN_4659 : dirty_0_37; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5558 = _GEN_901 ? _GEN_4660 : dirty_0_38; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5559 = _GEN_901 ? _GEN_4661 : dirty_0_39; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5560 = _GEN_901 ? _GEN_4662 : dirty_0_40; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5561 = _GEN_901 ? _GEN_4663 : dirty_0_41; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5562 = _GEN_901 ? _GEN_4664 : dirty_0_42; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5563 = _GEN_901 ? _GEN_4665 : dirty_0_43; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5564 = _GEN_901 ? _GEN_4666 : dirty_0_44; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5565 = _GEN_901 ? _GEN_4667 : dirty_0_45; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5566 = _GEN_901 ? _GEN_4668 : dirty_0_46; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5567 = _GEN_901 ? _GEN_4669 : dirty_0_47; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5568 = _GEN_901 ? _GEN_4670 : dirty_0_48; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5569 = _GEN_901 ? _GEN_4671 : dirty_0_49; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5570 = _GEN_901 ? _GEN_4672 : dirty_0_50; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5571 = _GEN_901 ? _GEN_4673 : dirty_0_51; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5572 = _GEN_901 ? _GEN_4674 : dirty_0_52; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5573 = _GEN_901 ? _GEN_4675 : dirty_0_53; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5574 = _GEN_901 ? _GEN_4676 : dirty_0_54; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5575 = _GEN_901 ? _GEN_4677 : dirty_0_55; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5576 = _GEN_901 ? _GEN_4678 : dirty_0_56; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5577 = _GEN_901 ? _GEN_4679 : dirty_0_57; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5578 = _GEN_901 ? _GEN_4680 : dirty_0_58; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5579 = _GEN_901 ? _GEN_4681 : dirty_0_59; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5580 = _GEN_901 ? _GEN_4682 : dirty_0_60; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5581 = _GEN_901 ? _GEN_4683 : dirty_0_61; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5582 = _GEN_901 ? _GEN_4684 : dirty_0_62; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5583 = _GEN_901 ? _GEN_4685 : dirty_0_63; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5584 = _GEN_901 ? _GEN_4686 : dirty_0_64; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5585 = _GEN_901 ? _GEN_4687 : dirty_0_65; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5586 = _GEN_901 ? _GEN_4688 : dirty_0_66; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5587 = _GEN_901 ? _GEN_4689 : dirty_0_67; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5588 = _GEN_901 ? _GEN_4690 : dirty_0_68; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5589 = _GEN_901 ? _GEN_4691 : dirty_0_69; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5590 = _GEN_901 ? _GEN_4692 : dirty_0_70; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5591 = _GEN_901 ? _GEN_4693 : dirty_0_71; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5592 = _GEN_901 ? _GEN_4694 : dirty_0_72; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5593 = _GEN_901 ? _GEN_4695 : dirty_0_73; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5594 = _GEN_901 ? _GEN_4696 : dirty_0_74; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5595 = _GEN_901 ? _GEN_4697 : dirty_0_75; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5596 = _GEN_901 ? _GEN_4698 : dirty_0_76; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5597 = _GEN_901 ? _GEN_4699 : dirty_0_77; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5598 = _GEN_901 ? _GEN_4700 : dirty_0_78; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5599 = _GEN_901 ? _GEN_4701 : dirty_0_79; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5600 = _GEN_901 ? _GEN_4702 : dirty_0_80; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5601 = _GEN_901 ? _GEN_4703 : dirty_0_81; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5602 = _GEN_901 ? _GEN_4704 : dirty_0_82; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5603 = _GEN_901 ? _GEN_4705 : dirty_0_83; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5604 = _GEN_901 ? _GEN_4706 : dirty_0_84; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5605 = _GEN_901 ? _GEN_4707 : dirty_0_85; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5606 = _GEN_901 ? _GEN_4708 : dirty_0_86; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5607 = _GEN_901 ? _GEN_4709 : dirty_0_87; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5608 = _GEN_901 ? _GEN_4710 : dirty_0_88; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5609 = _GEN_901 ? _GEN_4711 : dirty_0_89; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5610 = _GEN_901 ? _GEN_4712 : dirty_0_90; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5611 = _GEN_901 ? _GEN_4713 : dirty_0_91; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5612 = _GEN_901 ? _GEN_4714 : dirty_0_92; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5613 = _GEN_901 ? _GEN_4715 : dirty_0_93; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5614 = _GEN_901 ? _GEN_4716 : dirty_0_94; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5615 = _GEN_901 ? _GEN_4717 : dirty_0_95; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5616 = _GEN_901 ? _GEN_4718 : dirty_0_96; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5617 = _GEN_901 ? _GEN_4719 : dirty_0_97; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5618 = _GEN_901 ? _GEN_4720 : dirty_0_98; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5619 = _GEN_901 ? _GEN_4721 : dirty_0_99; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5620 = _GEN_901 ? _GEN_4722 : dirty_0_100; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5621 = _GEN_901 ? _GEN_4723 : dirty_0_101; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5622 = _GEN_901 ? _GEN_4724 : dirty_0_102; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5623 = _GEN_901 ? _GEN_4725 : dirty_0_103; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5624 = _GEN_901 ? _GEN_4726 : dirty_0_104; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5625 = _GEN_901 ? _GEN_4727 : dirty_0_105; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5626 = _GEN_901 ? _GEN_4728 : dirty_0_106; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5627 = _GEN_901 ? _GEN_4729 : dirty_0_107; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5628 = _GEN_901 ? _GEN_4730 : dirty_0_108; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5629 = _GEN_901 ? _GEN_4731 : dirty_0_109; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5630 = _GEN_901 ? _GEN_4732 : dirty_0_110; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5631 = _GEN_901 ? _GEN_4733 : dirty_0_111; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5632 = _GEN_901 ? _GEN_4734 : dirty_0_112; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5633 = _GEN_901 ? _GEN_4735 : dirty_0_113; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5634 = _GEN_901 ? _GEN_4736 : dirty_0_114; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5635 = _GEN_901 ? _GEN_4737 : dirty_0_115; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5636 = _GEN_901 ? _GEN_4738 : dirty_0_116; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5637 = _GEN_901 ? _GEN_4739 : dirty_0_117; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5638 = _GEN_901 ? _GEN_4740 : dirty_0_118; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5639 = _GEN_901 ? _GEN_4741 : dirty_0_119; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5640 = _GEN_901 ? _GEN_4742 : dirty_0_120; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5641 = _GEN_901 ? _GEN_4743 : dirty_0_121; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5642 = _GEN_901 ? _GEN_4744 : dirty_0_122; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5643 = _GEN_901 ? _GEN_4745 : dirty_0_123; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5644 = _GEN_901 ? _GEN_4746 : dirty_0_124; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5645 = _GEN_901 ? _GEN_4747 : dirty_0_125; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5646 = _GEN_901 ? _GEN_4748 : dirty_0_126; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5647 = _GEN_901 ? _GEN_4749 : dirty_0_127; // @[d_cache.scala 154:47 26:26]
  wire  _GEN_5648 = _GEN_901 ? _GEN_3470 : _GEN_3470; // @[d_cache.scala 154:47]
  wire  _GEN_5649 = _GEN_901 ? _GEN_3471 : _GEN_3471; // @[d_cache.scala 154:47]
  wire  _GEN_5650 = _GEN_901 ? _GEN_3472 : _GEN_3472; // @[d_cache.scala 154:47]
  wire  _GEN_5651 = _GEN_901 ? _GEN_3473 : _GEN_3473; // @[d_cache.scala 154:47]
  wire  _GEN_5652 = _GEN_901 ? _GEN_3474 : _GEN_3474; // @[d_cache.scala 154:47]
  wire  _GEN_5653 = _GEN_901 ? _GEN_3475 : _GEN_3475; // @[d_cache.scala 154:47]
  wire  _GEN_5654 = _GEN_901 ? _GEN_3476 : _GEN_3476; // @[d_cache.scala 154:47]
  wire  _GEN_5655 = _GEN_901 ? _GEN_3477 : _GEN_3477; // @[d_cache.scala 154:47]
  wire  _GEN_5656 = _GEN_901 ? _GEN_3478 : _GEN_3478; // @[d_cache.scala 154:47]
  wire  _GEN_5657 = _GEN_901 ? _GEN_3479 : _GEN_3479; // @[d_cache.scala 154:47]
  wire  _GEN_5658 = _GEN_901 ? _GEN_3480 : _GEN_3480; // @[d_cache.scala 154:47]
  wire  _GEN_5659 = _GEN_901 ? _GEN_3481 : _GEN_3481; // @[d_cache.scala 154:47]
  wire  _GEN_5660 = _GEN_901 ? _GEN_3482 : _GEN_3482; // @[d_cache.scala 154:47]
  wire  _GEN_5661 = _GEN_901 ? _GEN_3483 : _GEN_3483; // @[d_cache.scala 154:47]
  wire  _GEN_5662 = _GEN_901 ? _GEN_3484 : _GEN_3484; // @[d_cache.scala 154:47]
  wire  _GEN_5663 = _GEN_901 ? _GEN_3485 : _GEN_3485; // @[d_cache.scala 154:47]
  wire  _GEN_5664 = _GEN_901 ? _GEN_3486 : _GEN_3486; // @[d_cache.scala 154:47]
  wire  _GEN_5665 = _GEN_901 ? _GEN_3487 : _GEN_3487; // @[d_cache.scala 154:47]
  wire  _GEN_5666 = _GEN_901 ? _GEN_3488 : _GEN_3488; // @[d_cache.scala 154:47]
  wire  _GEN_5667 = _GEN_901 ? _GEN_3489 : _GEN_3489; // @[d_cache.scala 154:47]
  wire  _GEN_5668 = _GEN_901 ? _GEN_3490 : _GEN_3490; // @[d_cache.scala 154:47]
  wire  _GEN_5669 = _GEN_901 ? _GEN_3491 : _GEN_3491; // @[d_cache.scala 154:47]
  wire  _GEN_5670 = _GEN_901 ? _GEN_3492 : _GEN_3492; // @[d_cache.scala 154:47]
  wire  _GEN_5671 = _GEN_901 ? _GEN_3493 : _GEN_3493; // @[d_cache.scala 154:47]
  wire  _GEN_5672 = _GEN_901 ? _GEN_3494 : _GEN_3494; // @[d_cache.scala 154:47]
  wire  _GEN_5673 = _GEN_901 ? _GEN_3495 : _GEN_3495; // @[d_cache.scala 154:47]
  wire  _GEN_5674 = _GEN_901 ? _GEN_3496 : _GEN_3496; // @[d_cache.scala 154:47]
  wire  _GEN_5675 = _GEN_901 ? _GEN_3497 : _GEN_3497; // @[d_cache.scala 154:47]
  wire  _GEN_5676 = _GEN_901 ? _GEN_3498 : _GEN_3498; // @[d_cache.scala 154:47]
  wire  _GEN_5677 = _GEN_901 ? _GEN_3499 : _GEN_3499; // @[d_cache.scala 154:47]
  wire  _GEN_5678 = _GEN_901 ? _GEN_3500 : _GEN_3500; // @[d_cache.scala 154:47]
  wire  _GEN_5679 = _GEN_901 ? _GEN_3501 : _GEN_3501; // @[d_cache.scala 154:47]
  wire  _GEN_5680 = _GEN_901 ? _GEN_3502 : _GEN_3502; // @[d_cache.scala 154:47]
  wire  _GEN_5681 = _GEN_901 ? _GEN_3503 : _GEN_3503; // @[d_cache.scala 154:47]
  wire  _GEN_5682 = _GEN_901 ? _GEN_3504 : _GEN_3504; // @[d_cache.scala 154:47]
  wire  _GEN_5683 = _GEN_901 ? _GEN_3505 : _GEN_3505; // @[d_cache.scala 154:47]
  wire  _GEN_5684 = _GEN_901 ? _GEN_3506 : _GEN_3506; // @[d_cache.scala 154:47]
  wire  _GEN_5685 = _GEN_901 ? _GEN_3507 : _GEN_3507; // @[d_cache.scala 154:47]
  wire  _GEN_5686 = _GEN_901 ? _GEN_3508 : _GEN_3508; // @[d_cache.scala 154:47]
  wire  _GEN_5687 = _GEN_901 ? _GEN_3509 : _GEN_3509; // @[d_cache.scala 154:47]
  wire  _GEN_5688 = _GEN_901 ? _GEN_3510 : _GEN_3510; // @[d_cache.scala 154:47]
  wire  _GEN_5689 = _GEN_901 ? _GEN_3511 : _GEN_3511; // @[d_cache.scala 154:47]
  wire  _GEN_5690 = _GEN_901 ? _GEN_3512 : _GEN_3512; // @[d_cache.scala 154:47]
  wire  _GEN_5691 = _GEN_901 ? _GEN_3513 : _GEN_3513; // @[d_cache.scala 154:47]
  wire  _GEN_5692 = _GEN_901 ? _GEN_3514 : _GEN_3514; // @[d_cache.scala 154:47]
  wire  _GEN_5693 = _GEN_901 ? _GEN_3515 : _GEN_3515; // @[d_cache.scala 154:47]
  wire  _GEN_5694 = _GEN_901 ? _GEN_3516 : _GEN_3516; // @[d_cache.scala 154:47]
  wire  _GEN_5695 = _GEN_901 ? _GEN_3517 : _GEN_3517; // @[d_cache.scala 154:47]
  wire  _GEN_5696 = _GEN_901 ? _GEN_3518 : _GEN_3518; // @[d_cache.scala 154:47]
  wire  _GEN_5697 = _GEN_901 ? _GEN_3519 : _GEN_3519; // @[d_cache.scala 154:47]
  wire  _GEN_5698 = _GEN_901 ? _GEN_3520 : _GEN_3520; // @[d_cache.scala 154:47]
  wire  _GEN_5699 = _GEN_901 ? _GEN_3521 : _GEN_3521; // @[d_cache.scala 154:47]
  wire  _GEN_5700 = _GEN_901 ? _GEN_3522 : _GEN_3522; // @[d_cache.scala 154:47]
  wire  _GEN_5701 = _GEN_901 ? _GEN_3523 : _GEN_3523; // @[d_cache.scala 154:47]
  wire  _GEN_5702 = _GEN_901 ? _GEN_3524 : _GEN_3524; // @[d_cache.scala 154:47]
  wire  _GEN_5703 = _GEN_901 ? _GEN_3525 : _GEN_3525; // @[d_cache.scala 154:47]
  wire  _GEN_5704 = _GEN_901 ? _GEN_3526 : _GEN_3526; // @[d_cache.scala 154:47]
  wire  _GEN_5705 = _GEN_901 ? _GEN_3527 : _GEN_3527; // @[d_cache.scala 154:47]
  wire  _GEN_5706 = _GEN_901 ? _GEN_3528 : _GEN_3528; // @[d_cache.scala 154:47]
  wire  _GEN_5707 = _GEN_901 ? _GEN_3529 : _GEN_3529; // @[d_cache.scala 154:47]
  wire  _GEN_5708 = _GEN_901 ? _GEN_3530 : _GEN_3530; // @[d_cache.scala 154:47]
  wire  _GEN_5709 = _GEN_901 ? _GEN_3531 : _GEN_3531; // @[d_cache.scala 154:47]
  wire  _GEN_5710 = _GEN_901 ? _GEN_3532 : _GEN_3532; // @[d_cache.scala 154:47]
  wire  _GEN_5711 = _GEN_901 ? _GEN_3533 : _GEN_3533; // @[d_cache.scala 154:47]
  wire  _GEN_5712 = _GEN_901 ? _GEN_3534 : _GEN_3534; // @[d_cache.scala 154:47]
  wire  _GEN_5713 = _GEN_901 ? _GEN_3535 : _GEN_3535; // @[d_cache.scala 154:47]
  wire  _GEN_5714 = _GEN_901 ? _GEN_3536 : _GEN_3536; // @[d_cache.scala 154:47]
  wire  _GEN_5715 = _GEN_901 ? _GEN_3537 : _GEN_3537; // @[d_cache.scala 154:47]
  wire  _GEN_5716 = _GEN_901 ? _GEN_3538 : _GEN_3538; // @[d_cache.scala 154:47]
  wire  _GEN_5717 = _GEN_901 ? _GEN_3539 : _GEN_3539; // @[d_cache.scala 154:47]
  wire  _GEN_5718 = _GEN_901 ? _GEN_3540 : _GEN_3540; // @[d_cache.scala 154:47]
  wire  _GEN_5719 = _GEN_901 ? _GEN_3541 : _GEN_3541; // @[d_cache.scala 154:47]
  wire  _GEN_5720 = _GEN_901 ? _GEN_3542 : _GEN_3542; // @[d_cache.scala 154:47]
  wire  _GEN_5721 = _GEN_901 ? _GEN_3543 : _GEN_3543; // @[d_cache.scala 154:47]
  wire  _GEN_5722 = _GEN_901 ? _GEN_3544 : _GEN_3544; // @[d_cache.scala 154:47]
  wire  _GEN_5723 = _GEN_901 ? _GEN_3545 : _GEN_3545; // @[d_cache.scala 154:47]
  wire  _GEN_5724 = _GEN_901 ? _GEN_3546 : _GEN_3546; // @[d_cache.scala 154:47]
  wire  _GEN_5725 = _GEN_901 ? _GEN_3547 : _GEN_3547; // @[d_cache.scala 154:47]
  wire  _GEN_5726 = _GEN_901 ? _GEN_3548 : _GEN_3548; // @[d_cache.scala 154:47]
  wire  _GEN_5727 = _GEN_901 ? _GEN_3549 : _GEN_3549; // @[d_cache.scala 154:47]
  wire  _GEN_5728 = _GEN_901 ? _GEN_3550 : _GEN_3550; // @[d_cache.scala 154:47]
  wire  _GEN_5729 = _GEN_901 ? _GEN_3551 : _GEN_3551; // @[d_cache.scala 154:47]
  wire  _GEN_5730 = _GEN_901 ? _GEN_3552 : _GEN_3552; // @[d_cache.scala 154:47]
  wire  _GEN_5731 = _GEN_901 ? _GEN_3553 : _GEN_3553; // @[d_cache.scala 154:47]
  wire  _GEN_5732 = _GEN_901 ? _GEN_3554 : _GEN_3554; // @[d_cache.scala 154:47]
  wire  _GEN_5733 = _GEN_901 ? _GEN_3555 : _GEN_3555; // @[d_cache.scala 154:47]
  wire  _GEN_5734 = _GEN_901 ? _GEN_3556 : _GEN_3556; // @[d_cache.scala 154:47]
  wire  _GEN_5735 = _GEN_901 ? _GEN_3557 : _GEN_3557; // @[d_cache.scala 154:47]
  wire  _GEN_5736 = _GEN_901 ? _GEN_3558 : _GEN_3558; // @[d_cache.scala 154:47]
  wire  _GEN_5737 = _GEN_901 ? _GEN_3559 : _GEN_3559; // @[d_cache.scala 154:47]
  wire  _GEN_5738 = _GEN_901 ? _GEN_3560 : _GEN_3560; // @[d_cache.scala 154:47]
  wire  _GEN_5739 = _GEN_901 ? _GEN_3561 : _GEN_3561; // @[d_cache.scala 154:47]
  wire  _GEN_5740 = _GEN_901 ? _GEN_3562 : _GEN_3562; // @[d_cache.scala 154:47]
  wire  _GEN_5741 = _GEN_901 ? _GEN_3563 : _GEN_3563; // @[d_cache.scala 154:47]
  wire  _GEN_5742 = _GEN_901 ? _GEN_3564 : _GEN_3564; // @[d_cache.scala 154:47]
  wire  _GEN_5743 = _GEN_901 ? _GEN_3565 : _GEN_3565; // @[d_cache.scala 154:47]
  wire  _GEN_5744 = _GEN_901 ? _GEN_3566 : _GEN_3566; // @[d_cache.scala 154:47]
  wire  _GEN_5745 = _GEN_901 ? _GEN_3567 : _GEN_3567; // @[d_cache.scala 154:47]
  wire  _GEN_5746 = _GEN_901 ? _GEN_3568 : _GEN_3568; // @[d_cache.scala 154:47]
  wire  _GEN_5747 = _GEN_901 ? _GEN_3569 : _GEN_3569; // @[d_cache.scala 154:47]
  wire  _GEN_5748 = _GEN_901 ? _GEN_3570 : _GEN_3570; // @[d_cache.scala 154:47]
  wire  _GEN_5749 = _GEN_901 ? _GEN_3571 : _GEN_3571; // @[d_cache.scala 154:47]
  wire  _GEN_5750 = _GEN_901 ? _GEN_3572 : _GEN_3572; // @[d_cache.scala 154:47]
  wire  _GEN_5751 = _GEN_901 ? _GEN_3573 : _GEN_3573; // @[d_cache.scala 154:47]
  wire  _GEN_5752 = _GEN_901 ? _GEN_3574 : _GEN_3574; // @[d_cache.scala 154:47]
  wire  _GEN_5753 = _GEN_901 ? _GEN_3575 : _GEN_3575; // @[d_cache.scala 154:47]
  wire  _GEN_5754 = _GEN_901 ? _GEN_3576 : _GEN_3576; // @[d_cache.scala 154:47]
  wire  _GEN_5755 = _GEN_901 ? _GEN_3577 : _GEN_3577; // @[d_cache.scala 154:47]
  wire  _GEN_5756 = _GEN_901 ? _GEN_3578 : _GEN_3578; // @[d_cache.scala 154:47]
  wire  _GEN_5757 = _GEN_901 ? _GEN_3579 : _GEN_3579; // @[d_cache.scala 154:47]
  wire  _GEN_5758 = _GEN_901 ? _GEN_3580 : _GEN_3580; // @[d_cache.scala 154:47]
  wire  _GEN_5759 = _GEN_901 ? _GEN_3581 : _GEN_3581; // @[d_cache.scala 154:47]
  wire  _GEN_5760 = _GEN_901 ? _GEN_3582 : _GEN_3582; // @[d_cache.scala 154:47]
  wire  _GEN_5761 = _GEN_901 ? _GEN_3583 : _GEN_3583; // @[d_cache.scala 154:47]
  wire  _GEN_5762 = _GEN_901 ? _GEN_3584 : _GEN_3584; // @[d_cache.scala 154:47]
  wire  _GEN_5763 = _GEN_901 ? _GEN_3585 : _GEN_3585; // @[d_cache.scala 154:47]
  wire  _GEN_5764 = _GEN_901 ? _GEN_3586 : _GEN_3586; // @[d_cache.scala 154:47]
  wire  _GEN_5765 = _GEN_901 ? _GEN_3587 : _GEN_3587; // @[d_cache.scala 154:47]
  wire  _GEN_5766 = _GEN_901 ? _GEN_3588 : _GEN_3588; // @[d_cache.scala 154:47]
  wire  _GEN_5767 = _GEN_901 ? _GEN_3589 : _GEN_3589; // @[d_cache.scala 154:47]
  wire  _GEN_5768 = _GEN_901 ? _GEN_3590 : _GEN_3590; // @[d_cache.scala 154:47]
  wire  _GEN_5769 = _GEN_901 ? _GEN_3591 : _GEN_3591; // @[d_cache.scala 154:47]
  wire  _GEN_5770 = _GEN_901 ? _GEN_3592 : _GEN_3592; // @[d_cache.scala 154:47]
  wire  _GEN_5771 = _GEN_901 ? _GEN_3593 : _GEN_3593; // @[d_cache.scala 154:47]
  wire  _GEN_5772 = _GEN_901 ? _GEN_3594 : _GEN_3594; // @[d_cache.scala 154:47]
  wire  _GEN_5773 = _GEN_901 ? _GEN_3595 : _GEN_3595; // @[d_cache.scala 154:47]
  wire  _GEN_5774 = _GEN_901 ? _GEN_3596 : _GEN_3596; // @[d_cache.scala 154:47]
  wire  _GEN_5775 = _GEN_901 ? _GEN_3597 : _GEN_3597; // @[d_cache.scala 154:47]
  wire [2:0] _GEN_5776 = _GEN_901 ? 3'h6 : 3'h7; // @[d_cache.scala 154:47 161:31 164:31]
  wire [41:0] _write_back_addr_T_5 = {_GEN_384, 10'h0}; // @[d_cache.scala 173:58]
  wire [41:0] _write_back_addr_T_7 = _write_back_addr_T_5 | _GEN_18985; // @[d_cache.scala 173:65]
  wire  _GEN_6418 = 7'h0 == index[6:0] ? 1'h0 : dirty_1_0; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6419 = 7'h1 == index[6:0] ? 1'h0 : dirty_1_1; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6420 = 7'h2 == index[6:0] ? 1'h0 : dirty_1_2; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6421 = 7'h3 == index[6:0] ? 1'h0 : dirty_1_3; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6422 = 7'h4 == index[6:0] ? 1'h0 : dirty_1_4; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6423 = 7'h5 == index[6:0] ? 1'h0 : dirty_1_5; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6424 = 7'h6 == index[6:0] ? 1'h0 : dirty_1_6; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6425 = 7'h7 == index[6:0] ? 1'h0 : dirty_1_7; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6426 = 7'h8 == index[6:0] ? 1'h0 : dirty_1_8; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6427 = 7'h9 == index[6:0] ? 1'h0 : dirty_1_9; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6428 = 7'ha == index[6:0] ? 1'h0 : dirty_1_10; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6429 = 7'hb == index[6:0] ? 1'h0 : dirty_1_11; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6430 = 7'hc == index[6:0] ? 1'h0 : dirty_1_12; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6431 = 7'hd == index[6:0] ? 1'h0 : dirty_1_13; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6432 = 7'he == index[6:0] ? 1'h0 : dirty_1_14; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6433 = 7'hf == index[6:0] ? 1'h0 : dirty_1_15; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6434 = 7'h10 == index[6:0] ? 1'h0 : dirty_1_16; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6435 = 7'h11 == index[6:0] ? 1'h0 : dirty_1_17; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6436 = 7'h12 == index[6:0] ? 1'h0 : dirty_1_18; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6437 = 7'h13 == index[6:0] ? 1'h0 : dirty_1_19; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6438 = 7'h14 == index[6:0] ? 1'h0 : dirty_1_20; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6439 = 7'h15 == index[6:0] ? 1'h0 : dirty_1_21; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6440 = 7'h16 == index[6:0] ? 1'h0 : dirty_1_22; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6441 = 7'h17 == index[6:0] ? 1'h0 : dirty_1_23; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6442 = 7'h18 == index[6:0] ? 1'h0 : dirty_1_24; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6443 = 7'h19 == index[6:0] ? 1'h0 : dirty_1_25; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6444 = 7'h1a == index[6:0] ? 1'h0 : dirty_1_26; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6445 = 7'h1b == index[6:0] ? 1'h0 : dirty_1_27; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6446 = 7'h1c == index[6:0] ? 1'h0 : dirty_1_28; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6447 = 7'h1d == index[6:0] ? 1'h0 : dirty_1_29; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6448 = 7'h1e == index[6:0] ? 1'h0 : dirty_1_30; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6449 = 7'h1f == index[6:0] ? 1'h0 : dirty_1_31; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6450 = 7'h20 == index[6:0] ? 1'h0 : dirty_1_32; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6451 = 7'h21 == index[6:0] ? 1'h0 : dirty_1_33; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6452 = 7'h22 == index[6:0] ? 1'h0 : dirty_1_34; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6453 = 7'h23 == index[6:0] ? 1'h0 : dirty_1_35; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6454 = 7'h24 == index[6:0] ? 1'h0 : dirty_1_36; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6455 = 7'h25 == index[6:0] ? 1'h0 : dirty_1_37; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6456 = 7'h26 == index[6:0] ? 1'h0 : dirty_1_38; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6457 = 7'h27 == index[6:0] ? 1'h0 : dirty_1_39; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6458 = 7'h28 == index[6:0] ? 1'h0 : dirty_1_40; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6459 = 7'h29 == index[6:0] ? 1'h0 : dirty_1_41; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6460 = 7'h2a == index[6:0] ? 1'h0 : dirty_1_42; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6461 = 7'h2b == index[6:0] ? 1'h0 : dirty_1_43; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6462 = 7'h2c == index[6:0] ? 1'h0 : dirty_1_44; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6463 = 7'h2d == index[6:0] ? 1'h0 : dirty_1_45; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6464 = 7'h2e == index[6:0] ? 1'h0 : dirty_1_46; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6465 = 7'h2f == index[6:0] ? 1'h0 : dirty_1_47; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6466 = 7'h30 == index[6:0] ? 1'h0 : dirty_1_48; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6467 = 7'h31 == index[6:0] ? 1'h0 : dirty_1_49; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6468 = 7'h32 == index[6:0] ? 1'h0 : dirty_1_50; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6469 = 7'h33 == index[6:0] ? 1'h0 : dirty_1_51; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6470 = 7'h34 == index[6:0] ? 1'h0 : dirty_1_52; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6471 = 7'h35 == index[6:0] ? 1'h0 : dirty_1_53; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6472 = 7'h36 == index[6:0] ? 1'h0 : dirty_1_54; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6473 = 7'h37 == index[6:0] ? 1'h0 : dirty_1_55; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6474 = 7'h38 == index[6:0] ? 1'h0 : dirty_1_56; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6475 = 7'h39 == index[6:0] ? 1'h0 : dirty_1_57; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6476 = 7'h3a == index[6:0] ? 1'h0 : dirty_1_58; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6477 = 7'h3b == index[6:0] ? 1'h0 : dirty_1_59; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6478 = 7'h3c == index[6:0] ? 1'h0 : dirty_1_60; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6479 = 7'h3d == index[6:0] ? 1'h0 : dirty_1_61; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6480 = 7'h3e == index[6:0] ? 1'h0 : dirty_1_62; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6481 = 7'h3f == index[6:0] ? 1'h0 : dirty_1_63; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6482 = 7'h40 == index[6:0] ? 1'h0 : dirty_1_64; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6483 = 7'h41 == index[6:0] ? 1'h0 : dirty_1_65; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6484 = 7'h42 == index[6:0] ? 1'h0 : dirty_1_66; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6485 = 7'h43 == index[6:0] ? 1'h0 : dirty_1_67; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6486 = 7'h44 == index[6:0] ? 1'h0 : dirty_1_68; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6487 = 7'h45 == index[6:0] ? 1'h0 : dirty_1_69; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6488 = 7'h46 == index[6:0] ? 1'h0 : dirty_1_70; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6489 = 7'h47 == index[6:0] ? 1'h0 : dirty_1_71; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6490 = 7'h48 == index[6:0] ? 1'h0 : dirty_1_72; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6491 = 7'h49 == index[6:0] ? 1'h0 : dirty_1_73; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6492 = 7'h4a == index[6:0] ? 1'h0 : dirty_1_74; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6493 = 7'h4b == index[6:0] ? 1'h0 : dirty_1_75; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6494 = 7'h4c == index[6:0] ? 1'h0 : dirty_1_76; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6495 = 7'h4d == index[6:0] ? 1'h0 : dirty_1_77; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6496 = 7'h4e == index[6:0] ? 1'h0 : dirty_1_78; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6497 = 7'h4f == index[6:0] ? 1'h0 : dirty_1_79; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6498 = 7'h50 == index[6:0] ? 1'h0 : dirty_1_80; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6499 = 7'h51 == index[6:0] ? 1'h0 : dirty_1_81; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6500 = 7'h52 == index[6:0] ? 1'h0 : dirty_1_82; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6501 = 7'h53 == index[6:0] ? 1'h0 : dirty_1_83; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6502 = 7'h54 == index[6:0] ? 1'h0 : dirty_1_84; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6503 = 7'h55 == index[6:0] ? 1'h0 : dirty_1_85; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6504 = 7'h56 == index[6:0] ? 1'h0 : dirty_1_86; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6505 = 7'h57 == index[6:0] ? 1'h0 : dirty_1_87; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6506 = 7'h58 == index[6:0] ? 1'h0 : dirty_1_88; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6507 = 7'h59 == index[6:0] ? 1'h0 : dirty_1_89; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6508 = 7'h5a == index[6:0] ? 1'h0 : dirty_1_90; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6509 = 7'h5b == index[6:0] ? 1'h0 : dirty_1_91; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6510 = 7'h5c == index[6:0] ? 1'h0 : dirty_1_92; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6511 = 7'h5d == index[6:0] ? 1'h0 : dirty_1_93; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6512 = 7'h5e == index[6:0] ? 1'h0 : dirty_1_94; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6513 = 7'h5f == index[6:0] ? 1'h0 : dirty_1_95; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6514 = 7'h60 == index[6:0] ? 1'h0 : dirty_1_96; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6515 = 7'h61 == index[6:0] ? 1'h0 : dirty_1_97; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6516 = 7'h62 == index[6:0] ? 1'h0 : dirty_1_98; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6517 = 7'h63 == index[6:0] ? 1'h0 : dirty_1_99; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6518 = 7'h64 == index[6:0] ? 1'h0 : dirty_1_100; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6519 = 7'h65 == index[6:0] ? 1'h0 : dirty_1_101; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6520 = 7'h66 == index[6:0] ? 1'h0 : dirty_1_102; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6521 = 7'h67 == index[6:0] ? 1'h0 : dirty_1_103; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6522 = 7'h68 == index[6:0] ? 1'h0 : dirty_1_104; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6523 = 7'h69 == index[6:0] ? 1'h0 : dirty_1_105; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6524 = 7'h6a == index[6:0] ? 1'h0 : dirty_1_106; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6525 = 7'h6b == index[6:0] ? 1'h0 : dirty_1_107; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6526 = 7'h6c == index[6:0] ? 1'h0 : dirty_1_108; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6527 = 7'h6d == index[6:0] ? 1'h0 : dirty_1_109; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6528 = 7'h6e == index[6:0] ? 1'h0 : dirty_1_110; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6529 = 7'h6f == index[6:0] ? 1'h0 : dirty_1_111; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6530 = 7'h70 == index[6:0] ? 1'h0 : dirty_1_112; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6531 = 7'h71 == index[6:0] ? 1'h0 : dirty_1_113; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6532 = 7'h72 == index[6:0] ? 1'h0 : dirty_1_114; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6533 = 7'h73 == index[6:0] ? 1'h0 : dirty_1_115; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6534 = 7'h74 == index[6:0] ? 1'h0 : dirty_1_116; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6535 = 7'h75 == index[6:0] ? 1'h0 : dirty_1_117; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6536 = 7'h76 == index[6:0] ? 1'h0 : dirty_1_118; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6537 = 7'h77 == index[6:0] ? 1'h0 : dirty_1_119; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6538 = 7'h78 == index[6:0] ? 1'h0 : dirty_1_120; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6539 = 7'h79 == index[6:0] ? 1'h0 : dirty_1_121; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6540 = 7'h7a == index[6:0] ? 1'h0 : dirty_1_122; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6541 = 7'h7b == index[6:0] ? 1'h0 : dirty_1_123; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6542 = 7'h7c == index[6:0] ? 1'h0 : dirty_1_124; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6543 = 7'h7d == index[6:0] ? 1'h0 : dirty_1_125; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6544 = 7'h7e == index[6:0] ? 1'h0 : dirty_1_126; // @[d_cache.scala 176:{40,40} 27:26]
  wire  _GEN_6545 = 7'h7f == index[6:0] ? 1'h0 : dirty_1_127; // @[d_cache.scala 176:{40,40} 27:26]
  wire [63:0] _GEN_7058 = _GEN_1030 ? _GEN_1672 : write_back_data; // @[d_cache.scala 171:47 172:41 31:34]
  wire [41:0] _GEN_7059 = _GEN_1030 ? _write_back_addr_T_7 : {{10'd0}, write_back_addr}; // @[d_cache.scala 171:47 173:41 32:34]
  wire [63:0] _GEN_7060 = _GEN_1030 ? _GEN_3598 : _GEN_3598; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7061 = _GEN_1030 ? _GEN_3599 : _GEN_3599; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7062 = _GEN_1030 ? _GEN_3600 : _GEN_3600; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7063 = _GEN_1030 ? _GEN_3601 : _GEN_3601; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7064 = _GEN_1030 ? _GEN_3602 : _GEN_3602; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7065 = _GEN_1030 ? _GEN_3603 : _GEN_3603; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7066 = _GEN_1030 ? _GEN_3604 : _GEN_3604; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7067 = _GEN_1030 ? _GEN_3605 : _GEN_3605; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7068 = _GEN_1030 ? _GEN_3606 : _GEN_3606; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7069 = _GEN_1030 ? _GEN_3607 : _GEN_3607; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7070 = _GEN_1030 ? _GEN_3608 : _GEN_3608; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7071 = _GEN_1030 ? _GEN_3609 : _GEN_3609; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7072 = _GEN_1030 ? _GEN_3610 : _GEN_3610; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7073 = _GEN_1030 ? _GEN_3611 : _GEN_3611; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7074 = _GEN_1030 ? _GEN_3612 : _GEN_3612; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7075 = _GEN_1030 ? _GEN_3613 : _GEN_3613; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7076 = _GEN_1030 ? _GEN_3614 : _GEN_3614; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7077 = _GEN_1030 ? _GEN_3615 : _GEN_3615; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7078 = _GEN_1030 ? _GEN_3616 : _GEN_3616; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7079 = _GEN_1030 ? _GEN_3617 : _GEN_3617; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7080 = _GEN_1030 ? _GEN_3618 : _GEN_3618; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7081 = _GEN_1030 ? _GEN_3619 : _GEN_3619; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7082 = _GEN_1030 ? _GEN_3620 : _GEN_3620; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7083 = _GEN_1030 ? _GEN_3621 : _GEN_3621; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7084 = _GEN_1030 ? _GEN_3622 : _GEN_3622; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7085 = _GEN_1030 ? _GEN_3623 : _GEN_3623; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7086 = _GEN_1030 ? _GEN_3624 : _GEN_3624; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7087 = _GEN_1030 ? _GEN_3625 : _GEN_3625; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7088 = _GEN_1030 ? _GEN_3626 : _GEN_3626; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7089 = _GEN_1030 ? _GEN_3627 : _GEN_3627; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7090 = _GEN_1030 ? _GEN_3628 : _GEN_3628; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7091 = _GEN_1030 ? _GEN_3629 : _GEN_3629; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7092 = _GEN_1030 ? _GEN_3630 : _GEN_3630; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7093 = _GEN_1030 ? _GEN_3631 : _GEN_3631; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7094 = _GEN_1030 ? _GEN_3632 : _GEN_3632; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7095 = _GEN_1030 ? _GEN_3633 : _GEN_3633; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7096 = _GEN_1030 ? _GEN_3634 : _GEN_3634; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7097 = _GEN_1030 ? _GEN_3635 : _GEN_3635; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7098 = _GEN_1030 ? _GEN_3636 : _GEN_3636; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7099 = _GEN_1030 ? _GEN_3637 : _GEN_3637; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7100 = _GEN_1030 ? _GEN_3638 : _GEN_3638; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7101 = _GEN_1030 ? _GEN_3639 : _GEN_3639; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7102 = _GEN_1030 ? _GEN_3640 : _GEN_3640; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7103 = _GEN_1030 ? _GEN_3641 : _GEN_3641; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7104 = _GEN_1030 ? _GEN_3642 : _GEN_3642; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7105 = _GEN_1030 ? _GEN_3643 : _GEN_3643; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7106 = _GEN_1030 ? _GEN_3644 : _GEN_3644; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7107 = _GEN_1030 ? _GEN_3645 : _GEN_3645; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7108 = _GEN_1030 ? _GEN_3646 : _GEN_3646; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7109 = _GEN_1030 ? _GEN_3647 : _GEN_3647; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7110 = _GEN_1030 ? _GEN_3648 : _GEN_3648; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7111 = _GEN_1030 ? _GEN_3649 : _GEN_3649; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7112 = _GEN_1030 ? _GEN_3650 : _GEN_3650; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7113 = _GEN_1030 ? _GEN_3651 : _GEN_3651; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7114 = _GEN_1030 ? _GEN_3652 : _GEN_3652; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7115 = _GEN_1030 ? _GEN_3653 : _GEN_3653; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7116 = _GEN_1030 ? _GEN_3654 : _GEN_3654; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7117 = _GEN_1030 ? _GEN_3655 : _GEN_3655; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7118 = _GEN_1030 ? _GEN_3656 : _GEN_3656; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7119 = _GEN_1030 ? _GEN_3657 : _GEN_3657; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7120 = _GEN_1030 ? _GEN_3658 : _GEN_3658; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7121 = _GEN_1030 ? _GEN_3659 : _GEN_3659; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7122 = _GEN_1030 ? _GEN_3660 : _GEN_3660; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7123 = _GEN_1030 ? _GEN_3661 : _GEN_3661; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7124 = _GEN_1030 ? _GEN_3662 : _GEN_3662; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7125 = _GEN_1030 ? _GEN_3663 : _GEN_3663; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7126 = _GEN_1030 ? _GEN_3664 : _GEN_3664; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7127 = _GEN_1030 ? _GEN_3665 : _GEN_3665; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7128 = _GEN_1030 ? _GEN_3666 : _GEN_3666; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7129 = _GEN_1030 ? _GEN_3667 : _GEN_3667; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7130 = _GEN_1030 ? _GEN_3668 : _GEN_3668; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7131 = _GEN_1030 ? _GEN_3669 : _GEN_3669; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7132 = _GEN_1030 ? _GEN_3670 : _GEN_3670; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7133 = _GEN_1030 ? _GEN_3671 : _GEN_3671; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7134 = _GEN_1030 ? _GEN_3672 : _GEN_3672; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7135 = _GEN_1030 ? _GEN_3673 : _GEN_3673; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7136 = _GEN_1030 ? _GEN_3674 : _GEN_3674; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7137 = _GEN_1030 ? _GEN_3675 : _GEN_3675; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7138 = _GEN_1030 ? _GEN_3676 : _GEN_3676; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7139 = _GEN_1030 ? _GEN_3677 : _GEN_3677; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7140 = _GEN_1030 ? _GEN_3678 : _GEN_3678; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7141 = _GEN_1030 ? _GEN_3679 : _GEN_3679; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7142 = _GEN_1030 ? _GEN_3680 : _GEN_3680; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7143 = _GEN_1030 ? _GEN_3681 : _GEN_3681; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7144 = _GEN_1030 ? _GEN_3682 : _GEN_3682; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7145 = _GEN_1030 ? _GEN_3683 : _GEN_3683; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7146 = _GEN_1030 ? _GEN_3684 : _GEN_3684; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7147 = _GEN_1030 ? _GEN_3685 : _GEN_3685; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7148 = _GEN_1030 ? _GEN_3686 : _GEN_3686; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7149 = _GEN_1030 ? _GEN_3687 : _GEN_3687; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7150 = _GEN_1030 ? _GEN_3688 : _GEN_3688; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7151 = _GEN_1030 ? _GEN_3689 : _GEN_3689; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7152 = _GEN_1030 ? _GEN_3690 : _GEN_3690; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7153 = _GEN_1030 ? _GEN_3691 : _GEN_3691; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7154 = _GEN_1030 ? _GEN_3692 : _GEN_3692; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7155 = _GEN_1030 ? _GEN_3693 : _GEN_3693; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7156 = _GEN_1030 ? _GEN_3694 : _GEN_3694; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7157 = _GEN_1030 ? _GEN_3695 : _GEN_3695; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7158 = _GEN_1030 ? _GEN_3696 : _GEN_3696; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7159 = _GEN_1030 ? _GEN_3697 : _GEN_3697; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7160 = _GEN_1030 ? _GEN_3698 : _GEN_3698; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7161 = _GEN_1030 ? _GEN_3699 : _GEN_3699; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7162 = _GEN_1030 ? _GEN_3700 : _GEN_3700; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7163 = _GEN_1030 ? _GEN_3701 : _GEN_3701; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7164 = _GEN_1030 ? _GEN_3702 : _GEN_3702; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7165 = _GEN_1030 ? _GEN_3703 : _GEN_3703; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7166 = _GEN_1030 ? _GEN_3704 : _GEN_3704; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7167 = _GEN_1030 ? _GEN_3705 : _GEN_3705; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7168 = _GEN_1030 ? _GEN_3706 : _GEN_3706; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7169 = _GEN_1030 ? _GEN_3707 : _GEN_3707; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7170 = _GEN_1030 ? _GEN_3708 : _GEN_3708; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7171 = _GEN_1030 ? _GEN_3709 : _GEN_3709; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7172 = _GEN_1030 ? _GEN_3710 : _GEN_3710; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7173 = _GEN_1030 ? _GEN_3711 : _GEN_3711; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7174 = _GEN_1030 ? _GEN_3712 : _GEN_3712; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7175 = _GEN_1030 ? _GEN_3713 : _GEN_3713; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7176 = _GEN_1030 ? _GEN_3714 : _GEN_3714; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7177 = _GEN_1030 ? _GEN_3715 : _GEN_3715; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7178 = _GEN_1030 ? _GEN_3716 : _GEN_3716; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7179 = _GEN_1030 ? _GEN_3717 : _GEN_3717; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7180 = _GEN_1030 ? _GEN_3718 : _GEN_3718; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7181 = _GEN_1030 ? _GEN_3719 : _GEN_3719; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7182 = _GEN_1030 ? _GEN_3720 : _GEN_3720; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7183 = _GEN_1030 ? _GEN_3721 : _GEN_3721; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7184 = _GEN_1030 ? _GEN_3722 : _GEN_3722; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7185 = _GEN_1030 ? _GEN_3723 : _GEN_3723; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7186 = _GEN_1030 ? _GEN_3724 : _GEN_3724; // @[d_cache.scala 171:47]
  wire [63:0] _GEN_7187 = _GEN_1030 ? _GEN_3725 : _GEN_3725; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7188 = _GEN_1030 ? _GEN_3726 : _GEN_3726; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7189 = _GEN_1030 ? _GEN_3727 : _GEN_3727; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7190 = _GEN_1030 ? _GEN_3728 : _GEN_3728; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7191 = _GEN_1030 ? _GEN_3729 : _GEN_3729; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7192 = _GEN_1030 ? _GEN_3730 : _GEN_3730; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7193 = _GEN_1030 ? _GEN_3731 : _GEN_3731; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7194 = _GEN_1030 ? _GEN_3732 : _GEN_3732; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7195 = _GEN_1030 ? _GEN_3733 : _GEN_3733; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7196 = _GEN_1030 ? _GEN_3734 : _GEN_3734; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7197 = _GEN_1030 ? _GEN_3735 : _GEN_3735; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7198 = _GEN_1030 ? _GEN_3736 : _GEN_3736; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7199 = _GEN_1030 ? _GEN_3737 : _GEN_3737; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7200 = _GEN_1030 ? _GEN_3738 : _GEN_3738; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7201 = _GEN_1030 ? _GEN_3739 : _GEN_3739; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7202 = _GEN_1030 ? _GEN_3740 : _GEN_3740; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7203 = _GEN_1030 ? _GEN_3741 : _GEN_3741; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7204 = _GEN_1030 ? _GEN_3742 : _GEN_3742; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7205 = _GEN_1030 ? _GEN_3743 : _GEN_3743; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7206 = _GEN_1030 ? _GEN_3744 : _GEN_3744; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7207 = _GEN_1030 ? _GEN_3745 : _GEN_3745; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7208 = _GEN_1030 ? _GEN_3746 : _GEN_3746; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7209 = _GEN_1030 ? _GEN_3747 : _GEN_3747; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7210 = _GEN_1030 ? _GEN_3748 : _GEN_3748; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7211 = _GEN_1030 ? _GEN_3749 : _GEN_3749; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7212 = _GEN_1030 ? _GEN_3750 : _GEN_3750; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7213 = _GEN_1030 ? _GEN_3751 : _GEN_3751; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7214 = _GEN_1030 ? _GEN_3752 : _GEN_3752; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7215 = _GEN_1030 ? _GEN_3753 : _GEN_3753; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7216 = _GEN_1030 ? _GEN_3754 : _GEN_3754; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7217 = _GEN_1030 ? _GEN_3755 : _GEN_3755; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7218 = _GEN_1030 ? _GEN_3756 : _GEN_3756; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7219 = _GEN_1030 ? _GEN_3757 : _GEN_3757; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7220 = _GEN_1030 ? _GEN_3758 : _GEN_3758; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7221 = _GEN_1030 ? _GEN_3759 : _GEN_3759; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7222 = _GEN_1030 ? _GEN_3760 : _GEN_3760; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7223 = _GEN_1030 ? _GEN_3761 : _GEN_3761; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7224 = _GEN_1030 ? _GEN_3762 : _GEN_3762; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7225 = _GEN_1030 ? _GEN_3763 : _GEN_3763; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7226 = _GEN_1030 ? _GEN_3764 : _GEN_3764; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7227 = _GEN_1030 ? _GEN_3765 : _GEN_3765; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7228 = _GEN_1030 ? _GEN_3766 : _GEN_3766; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7229 = _GEN_1030 ? _GEN_3767 : _GEN_3767; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7230 = _GEN_1030 ? _GEN_3768 : _GEN_3768; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7231 = _GEN_1030 ? _GEN_3769 : _GEN_3769; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7232 = _GEN_1030 ? _GEN_3770 : _GEN_3770; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7233 = _GEN_1030 ? _GEN_3771 : _GEN_3771; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7234 = _GEN_1030 ? _GEN_3772 : _GEN_3772; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7235 = _GEN_1030 ? _GEN_3773 : _GEN_3773; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7236 = _GEN_1030 ? _GEN_3774 : _GEN_3774; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7237 = _GEN_1030 ? _GEN_3775 : _GEN_3775; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7238 = _GEN_1030 ? _GEN_3776 : _GEN_3776; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7239 = _GEN_1030 ? _GEN_3777 : _GEN_3777; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7240 = _GEN_1030 ? _GEN_3778 : _GEN_3778; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7241 = _GEN_1030 ? _GEN_3779 : _GEN_3779; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7242 = _GEN_1030 ? _GEN_3780 : _GEN_3780; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7243 = _GEN_1030 ? _GEN_3781 : _GEN_3781; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7244 = _GEN_1030 ? _GEN_3782 : _GEN_3782; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7245 = _GEN_1030 ? _GEN_3783 : _GEN_3783; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7246 = _GEN_1030 ? _GEN_3784 : _GEN_3784; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7247 = _GEN_1030 ? _GEN_3785 : _GEN_3785; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7248 = _GEN_1030 ? _GEN_3786 : _GEN_3786; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7249 = _GEN_1030 ? _GEN_3787 : _GEN_3787; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7250 = _GEN_1030 ? _GEN_3788 : _GEN_3788; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7251 = _GEN_1030 ? _GEN_3789 : _GEN_3789; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7252 = _GEN_1030 ? _GEN_3790 : _GEN_3790; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7253 = _GEN_1030 ? _GEN_3791 : _GEN_3791; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7254 = _GEN_1030 ? _GEN_3792 : _GEN_3792; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7255 = _GEN_1030 ? _GEN_3793 : _GEN_3793; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7256 = _GEN_1030 ? _GEN_3794 : _GEN_3794; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7257 = _GEN_1030 ? _GEN_3795 : _GEN_3795; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7258 = _GEN_1030 ? _GEN_3796 : _GEN_3796; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7259 = _GEN_1030 ? _GEN_3797 : _GEN_3797; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7260 = _GEN_1030 ? _GEN_3798 : _GEN_3798; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7261 = _GEN_1030 ? _GEN_3799 : _GEN_3799; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7262 = _GEN_1030 ? _GEN_3800 : _GEN_3800; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7263 = _GEN_1030 ? _GEN_3801 : _GEN_3801; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7264 = _GEN_1030 ? _GEN_3802 : _GEN_3802; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7265 = _GEN_1030 ? _GEN_3803 : _GEN_3803; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7266 = _GEN_1030 ? _GEN_3804 : _GEN_3804; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7267 = _GEN_1030 ? _GEN_3805 : _GEN_3805; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7268 = _GEN_1030 ? _GEN_3806 : _GEN_3806; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7269 = _GEN_1030 ? _GEN_3807 : _GEN_3807; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7270 = _GEN_1030 ? _GEN_3808 : _GEN_3808; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7271 = _GEN_1030 ? _GEN_3809 : _GEN_3809; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7272 = _GEN_1030 ? _GEN_3810 : _GEN_3810; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7273 = _GEN_1030 ? _GEN_3811 : _GEN_3811; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7274 = _GEN_1030 ? _GEN_3812 : _GEN_3812; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7275 = _GEN_1030 ? _GEN_3813 : _GEN_3813; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7276 = _GEN_1030 ? _GEN_3814 : _GEN_3814; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7277 = _GEN_1030 ? _GEN_3815 : _GEN_3815; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7278 = _GEN_1030 ? _GEN_3816 : _GEN_3816; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7279 = _GEN_1030 ? _GEN_3817 : _GEN_3817; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7280 = _GEN_1030 ? _GEN_3818 : _GEN_3818; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7281 = _GEN_1030 ? _GEN_3819 : _GEN_3819; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7282 = _GEN_1030 ? _GEN_3820 : _GEN_3820; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7283 = _GEN_1030 ? _GEN_3821 : _GEN_3821; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7284 = _GEN_1030 ? _GEN_3822 : _GEN_3822; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7285 = _GEN_1030 ? _GEN_3823 : _GEN_3823; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7286 = _GEN_1030 ? _GEN_3824 : _GEN_3824; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7287 = _GEN_1030 ? _GEN_3825 : _GEN_3825; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7288 = _GEN_1030 ? _GEN_3826 : _GEN_3826; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7289 = _GEN_1030 ? _GEN_3827 : _GEN_3827; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7290 = _GEN_1030 ? _GEN_3828 : _GEN_3828; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7291 = _GEN_1030 ? _GEN_3829 : _GEN_3829; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7292 = _GEN_1030 ? _GEN_3830 : _GEN_3830; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7293 = _GEN_1030 ? _GEN_3831 : _GEN_3831; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7294 = _GEN_1030 ? _GEN_3832 : _GEN_3832; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7295 = _GEN_1030 ? _GEN_3833 : _GEN_3833; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7296 = _GEN_1030 ? _GEN_3834 : _GEN_3834; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7297 = _GEN_1030 ? _GEN_3835 : _GEN_3835; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7298 = _GEN_1030 ? _GEN_3836 : _GEN_3836; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7299 = _GEN_1030 ? _GEN_3837 : _GEN_3837; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7300 = _GEN_1030 ? _GEN_3838 : _GEN_3838; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7301 = _GEN_1030 ? _GEN_3839 : _GEN_3839; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7302 = _GEN_1030 ? _GEN_3840 : _GEN_3840; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7303 = _GEN_1030 ? _GEN_3841 : _GEN_3841; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7304 = _GEN_1030 ? _GEN_3842 : _GEN_3842; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7305 = _GEN_1030 ? _GEN_3843 : _GEN_3843; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7306 = _GEN_1030 ? _GEN_3844 : _GEN_3844; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7307 = _GEN_1030 ? _GEN_3845 : _GEN_3845; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7308 = _GEN_1030 ? _GEN_3846 : _GEN_3846; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7309 = _GEN_1030 ? _GEN_3847 : _GEN_3847; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7310 = _GEN_1030 ? _GEN_3848 : _GEN_3848; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7311 = _GEN_1030 ? _GEN_3849 : _GEN_3849; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7312 = _GEN_1030 ? _GEN_3850 : _GEN_3850; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7313 = _GEN_1030 ? _GEN_3851 : _GEN_3851; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7314 = _GEN_1030 ? _GEN_3852 : _GEN_3852; // @[d_cache.scala 171:47]
  wire [31:0] _GEN_7315 = _GEN_1030 ? _GEN_3853 : _GEN_3853; // @[d_cache.scala 171:47]
  wire  _GEN_7316 = _GEN_1030 ? _GEN_6418 : dirty_1_0; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7317 = _GEN_1030 ? _GEN_6419 : dirty_1_1; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7318 = _GEN_1030 ? _GEN_6420 : dirty_1_2; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7319 = _GEN_1030 ? _GEN_6421 : dirty_1_3; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7320 = _GEN_1030 ? _GEN_6422 : dirty_1_4; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7321 = _GEN_1030 ? _GEN_6423 : dirty_1_5; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7322 = _GEN_1030 ? _GEN_6424 : dirty_1_6; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7323 = _GEN_1030 ? _GEN_6425 : dirty_1_7; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7324 = _GEN_1030 ? _GEN_6426 : dirty_1_8; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7325 = _GEN_1030 ? _GEN_6427 : dirty_1_9; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7326 = _GEN_1030 ? _GEN_6428 : dirty_1_10; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7327 = _GEN_1030 ? _GEN_6429 : dirty_1_11; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7328 = _GEN_1030 ? _GEN_6430 : dirty_1_12; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7329 = _GEN_1030 ? _GEN_6431 : dirty_1_13; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7330 = _GEN_1030 ? _GEN_6432 : dirty_1_14; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7331 = _GEN_1030 ? _GEN_6433 : dirty_1_15; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7332 = _GEN_1030 ? _GEN_6434 : dirty_1_16; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7333 = _GEN_1030 ? _GEN_6435 : dirty_1_17; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7334 = _GEN_1030 ? _GEN_6436 : dirty_1_18; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7335 = _GEN_1030 ? _GEN_6437 : dirty_1_19; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7336 = _GEN_1030 ? _GEN_6438 : dirty_1_20; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7337 = _GEN_1030 ? _GEN_6439 : dirty_1_21; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7338 = _GEN_1030 ? _GEN_6440 : dirty_1_22; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7339 = _GEN_1030 ? _GEN_6441 : dirty_1_23; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7340 = _GEN_1030 ? _GEN_6442 : dirty_1_24; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7341 = _GEN_1030 ? _GEN_6443 : dirty_1_25; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7342 = _GEN_1030 ? _GEN_6444 : dirty_1_26; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7343 = _GEN_1030 ? _GEN_6445 : dirty_1_27; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7344 = _GEN_1030 ? _GEN_6446 : dirty_1_28; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7345 = _GEN_1030 ? _GEN_6447 : dirty_1_29; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7346 = _GEN_1030 ? _GEN_6448 : dirty_1_30; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7347 = _GEN_1030 ? _GEN_6449 : dirty_1_31; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7348 = _GEN_1030 ? _GEN_6450 : dirty_1_32; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7349 = _GEN_1030 ? _GEN_6451 : dirty_1_33; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7350 = _GEN_1030 ? _GEN_6452 : dirty_1_34; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7351 = _GEN_1030 ? _GEN_6453 : dirty_1_35; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7352 = _GEN_1030 ? _GEN_6454 : dirty_1_36; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7353 = _GEN_1030 ? _GEN_6455 : dirty_1_37; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7354 = _GEN_1030 ? _GEN_6456 : dirty_1_38; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7355 = _GEN_1030 ? _GEN_6457 : dirty_1_39; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7356 = _GEN_1030 ? _GEN_6458 : dirty_1_40; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7357 = _GEN_1030 ? _GEN_6459 : dirty_1_41; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7358 = _GEN_1030 ? _GEN_6460 : dirty_1_42; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7359 = _GEN_1030 ? _GEN_6461 : dirty_1_43; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7360 = _GEN_1030 ? _GEN_6462 : dirty_1_44; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7361 = _GEN_1030 ? _GEN_6463 : dirty_1_45; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7362 = _GEN_1030 ? _GEN_6464 : dirty_1_46; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7363 = _GEN_1030 ? _GEN_6465 : dirty_1_47; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7364 = _GEN_1030 ? _GEN_6466 : dirty_1_48; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7365 = _GEN_1030 ? _GEN_6467 : dirty_1_49; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7366 = _GEN_1030 ? _GEN_6468 : dirty_1_50; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7367 = _GEN_1030 ? _GEN_6469 : dirty_1_51; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7368 = _GEN_1030 ? _GEN_6470 : dirty_1_52; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7369 = _GEN_1030 ? _GEN_6471 : dirty_1_53; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7370 = _GEN_1030 ? _GEN_6472 : dirty_1_54; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7371 = _GEN_1030 ? _GEN_6473 : dirty_1_55; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7372 = _GEN_1030 ? _GEN_6474 : dirty_1_56; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7373 = _GEN_1030 ? _GEN_6475 : dirty_1_57; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7374 = _GEN_1030 ? _GEN_6476 : dirty_1_58; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7375 = _GEN_1030 ? _GEN_6477 : dirty_1_59; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7376 = _GEN_1030 ? _GEN_6478 : dirty_1_60; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7377 = _GEN_1030 ? _GEN_6479 : dirty_1_61; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7378 = _GEN_1030 ? _GEN_6480 : dirty_1_62; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7379 = _GEN_1030 ? _GEN_6481 : dirty_1_63; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7380 = _GEN_1030 ? _GEN_6482 : dirty_1_64; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7381 = _GEN_1030 ? _GEN_6483 : dirty_1_65; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7382 = _GEN_1030 ? _GEN_6484 : dirty_1_66; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7383 = _GEN_1030 ? _GEN_6485 : dirty_1_67; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7384 = _GEN_1030 ? _GEN_6486 : dirty_1_68; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7385 = _GEN_1030 ? _GEN_6487 : dirty_1_69; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7386 = _GEN_1030 ? _GEN_6488 : dirty_1_70; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7387 = _GEN_1030 ? _GEN_6489 : dirty_1_71; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7388 = _GEN_1030 ? _GEN_6490 : dirty_1_72; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7389 = _GEN_1030 ? _GEN_6491 : dirty_1_73; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7390 = _GEN_1030 ? _GEN_6492 : dirty_1_74; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7391 = _GEN_1030 ? _GEN_6493 : dirty_1_75; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7392 = _GEN_1030 ? _GEN_6494 : dirty_1_76; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7393 = _GEN_1030 ? _GEN_6495 : dirty_1_77; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7394 = _GEN_1030 ? _GEN_6496 : dirty_1_78; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7395 = _GEN_1030 ? _GEN_6497 : dirty_1_79; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7396 = _GEN_1030 ? _GEN_6498 : dirty_1_80; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7397 = _GEN_1030 ? _GEN_6499 : dirty_1_81; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7398 = _GEN_1030 ? _GEN_6500 : dirty_1_82; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7399 = _GEN_1030 ? _GEN_6501 : dirty_1_83; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7400 = _GEN_1030 ? _GEN_6502 : dirty_1_84; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7401 = _GEN_1030 ? _GEN_6503 : dirty_1_85; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7402 = _GEN_1030 ? _GEN_6504 : dirty_1_86; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7403 = _GEN_1030 ? _GEN_6505 : dirty_1_87; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7404 = _GEN_1030 ? _GEN_6506 : dirty_1_88; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7405 = _GEN_1030 ? _GEN_6507 : dirty_1_89; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7406 = _GEN_1030 ? _GEN_6508 : dirty_1_90; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7407 = _GEN_1030 ? _GEN_6509 : dirty_1_91; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7408 = _GEN_1030 ? _GEN_6510 : dirty_1_92; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7409 = _GEN_1030 ? _GEN_6511 : dirty_1_93; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7410 = _GEN_1030 ? _GEN_6512 : dirty_1_94; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7411 = _GEN_1030 ? _GEN_6513 : dirty_1_95; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7412 = _GEN_1030 ? _GEN_6514 : dirty_1_96; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7413 = _GEN_1030 ? _GEN_6515 : dirty_1_97; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7414 = _GEN_1030 ? _GEN_6516 : dirty_1_98; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7415 = _GEN_1030 ? _GEN_6517 : dirty_1_99; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7416 = _GEN_1030 ? _GEN_6518 : dirty_1_100; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7417 = _GEN_1030 ? _GEN_6519 : dirty_1_101; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7418 = _GEN_1030 ? _GEN_6520 : dirty_1_102; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7419 = _GEN_1030 ? _GEN_6521 : dirty_1_103; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7420 = _GEN_1030 ? _GEN_6522 : dirty_1_104; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7421 = _GEN_1030 ? _GEN_6523 : dirty_1_105; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7422 = _GEN_1030 ? _GEN_6524 : dirty_1_106; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7423 = _GEN_1030 ? _GEN_6525 : dirty_1_107; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7424 = _GEN_1030 ? _GEN_6526 : dirty_1_108; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7425 = _GEN_1030 ? _GEN_6527 : dirty_1_109; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7426 = _GEN_1030 ? _GEN_6528 : dirty_1_110; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7427 = _GEN_1030 ? _GEN_6529 : dirty_1_111; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7428 = _GEN_1030 ? _GEN_6530 : dirty_1_112; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7429 = _GEN_1030 ? _GEN_6531 : dirty_1_113; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7430 = _GEN_1030 ? _GEN_6532 : dirty_1_114; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7431 = _GEN_1030 ? _GEN_6533 : dirty_1_115; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7432 = _GEN_1030 ? _GEN_6534 : dirty_1_116; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7433 = _GEN_1030 ? _GEN_6535 : dirty_1_117; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7434 = _GEN_1030 ? _GEN_6536 : dirty_1_118; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7435 = _GEN_1030 ? _GEN_6537 : dirty_1_119; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7436 = _GEN_1030 ? _GEN_6538 : dirty_1_120; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7437 = _GEN_1030 ? _GEN_6539 : dirty_1_121; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7438 = _GEN_1030 ? _GEN_6540 : dirty_1_122; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7439 = _GEN_1030 ? _GEN_6541 : dirty_1_123; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7440 = _GEN_1030 ? _GEN_6542 : dirty_1_124; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7441 = _GEN_1030 ? _GEN_6543 : dirty_1_125; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7442 = _GEN_1030 ? _GEN_6544 : dirty_1_126; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7443 = _GEN_1030 ? _GEN_6545 : dirty_1_127; // @[d_cache.scala 171:47 27:26]
  wire  _GEN_7444 = _GEN_1030 ? _GEN_3854 : _GEN_3854; // @[d_cache.scala 171:47]
  wire  _GEN_7445 = _GEN_1030 ? _GEN_3855 : _GEN_3855; // @[d_cache.scala 171:47]
  wire  _GEN_7446 = _GEN_1030 ? _GEN_3856 : _GEN_3856; // @[d_cache.scala 171:47]
  wire  _GEN_7447 = _GEN_1030 ? _GEN_3857 : _GEN_3857; // @[d_cache.scala 171:47]
  wire  _GEN_7448 = _GEN_1030 ? _GEN_3858 : _GEN_3858; // @[d_cache.scala 171:47]
  wire  _GEN_7449 = _GEN_1030 ? _GEN_3859 : _GEN_3859; // @[d_cache.scala 171:47]
  wire  _GEN_7450 = _GEN_1030 ? _GEN_3860 : _GEN_3860; // @[d_cache.scala 171:47]
  wire  _GEN_7451 = _GEN_1030 ? _GEN_3861 : _GEN_3861; // @[d_cache.scala 171:47]
  wire  _GEN_7452 = _GEN_1030 ? _GEN_3862 : _GEN_3862; // @[d_cache.scala 171:47]
  wire  _GEN_7453 = _GEN_1030 ? _GEN_3863 : _GEN_3863; // @[d_cache.scala 171:47]
  wire  _GEN_7454 = _GEN_1030 ? _GEN_3864 : _GEN_3864; // @[d_cache.scala 171:47]
  wire  _GEN_7455 = _GEN_1030 ? _GEN_3865 : _GEN_3865; // @[d_cache.scala 171:47]
  wire  _GEN_7456 = _GEN_1030 ? _GEN_3866 : _GEN_3866; // @[d_cache.scala 171:47]
  wire  _GEN_7457 = _GEN_1030 ? _GEN_3867 : _GEN_3867; // @[d_cache.scala 171:47]
  wire  _GEN_7458 = _GEN_1030 ? _GEN_3868 : _GEN_3868; // @[d_cache.scala 171:47]
  wire  _GEN_7459 = _GEN_1030 ? _GEN_3869 : _GEN_3869; // @[d_cache.scala 171:47]
  wire  _GEN_7460 = _GEN_1030 ? _GEN_3870 : _GEN_3870; // @[d_cache.scala 171:47]
  wire  _GEN_7461 = _GEN_1030 ? _GEN_3871 : _GEN_3871; // @[d_cache.scala 171:47]
  wire  _GEN_7462 = _GEN_1030 ? _GEN_3872 : _GEN_3872; // @[d_cache.scala 171:47]
  wire  _GEN_7463 = _GEN_1030 ? _GEN_3873 : _GEN_3873; // @[d_cache.scala 171:47]
  wire  _GEN_7464 = _GEN_1030 ? _GEN_3874 : _GEN_3874; // @[d_cache.scala 171:47]
  wire  _GEN_7465 = _GEN_1030 ? _GEN_3875 : _GEN_3875; // @[d_cache.scala 171:47]
  wire  _GEN_7466 = _GEN_1030 ? _GEN_3876 : _GEN_3876; // @[d_cache.scala 171:47]
  wire  _GEN_7467 = _GEN_1030 ? _GEN_3877 : _GEN_3877; // @[d_cache.scala 171:47]
  wire  _GEN_7468 = _GEN_1030 ? _GEN_3878 : _GEN_3878; // @[d_cache.scala 171:47]
  wire  _GEN_7469 = _GEN_1030 ? _GEN_3879 : _GEN_3879; // @[d_cache.scala 171:47]
  wire  _GEN_7470 = _GEN_1030 ? _GEN_3880 : _GEN_3880; // @[d_cache.scala 171:47]
  wire  _GEN_7471 = _GEN_1030 ? _GEN_3881 : _GEN_3881; // @[d_cache.scala 171:47]
  wire  _GEN_7472 = _GEN_1030 ? _GEN_3882 : _GEN_3882; // @[d_cache.scala 171:47]
  wire  _GEN_7473 = _GEN_1030 ? _GEN_3883 : _GEN_3883; // @[d_cache.scala 171:47]
  wire  _GEN_7474 = _GEN_1030 ? _GEN_3884 : _GEN_3884; // @[d_cache.scala 171:47]
  wire  _GEN_7475 = _GEN_1030 ? _GEN_3885 : _GEN_3885; // @[d_cache.scala 171:47]
  wire  _GEN_7476 = _GEN_1030 ? _GEN_3886 : _GEN_3886; // @[d_cache.scala 171:47]
  wire  _GEN_7477 = _GEN_1030 ? _GEN_3887 : _GEN_3887; // @[d_cache.scala 171:47]
  wire  _GEN_7478 = _GEN_1030 ? _GEN_3888 : _GEN_3888; // @[d_cache.scala 171:47]
  wire  _GEN_7479 = _GEN_1030 ? _GEN_3889 : _GEN_3889; // @[d_cache.scala 171:47]
  wire  _GEN_7480 = _GEN_1030 ? _GEN_3890 : _GEN_3890; // @[d_cache.scala 171:47]
  wire  _GEN_7481 = _GEN_1030 ? _GEN_3891 : _GEN_3891; // @[d_cache.scala 171:47]
  wire  _GEN_7482 = _GEN_1030 ? _GEN_3892 : _GEN_3892; // @[d_cache.scala 171:47]
  wire  _GEN_7483 = _GEN_1030 ? _GEN_3893 : _GEN_3893; // @[d_cache.scala 171:47]
  wire  _GEN_7484 = _GEN_1030 ? _GEN_3894 : _GEN_3894; // @[d_cache.scala 171:47]
  wire  _GEN_7485 = _GEN_1030 ? _GEN_3895 : _GEN_3895; // @[d_cache.scala 171:47]
  wire  _GEN_7486 = _GEN_1030 ? _GEN_3896 : _GEN_3896; // @[d_cache.scala 171:47]
  wire  _GEN_7487 = _GEN_1030 ? _GEN_3897 : _GEN_3897; // @[d_cache.scala 171:47]
  wire  _GEN_7488 = _GEN_1030 ? _GEN_3898 : _GEN_3898; // @[d_cache.scala 171:47]
  wire  _GEN_7489 = _GEN_1030 ? _GEN_3899 : _GEN_3899; // @[d_cache.scala 171:47]
  wire  _GEN_7490 = _GEN_1030 ? _GEN_3900 : _GEN_3900; // @[d_cache.scala 171:47]
  wire  _GEN_7491 = _GEN_1030 ? _GEN_3901 : _GEN_3901; // @[d_cache.scala 171:47]
  wire  _GEN_7492 = _GEN_1030 ? _GEN_3902 : _GEN_3902; // @[d_cache.scala 171:47]
  wire  _GEN_7493 = _GEN_1030 ? _GEN_3903 : _GEN_3903; // @[d_cache.scala 171:47]
  wire  _GEN_7494 = _GEN_1030 ? _GEN_3904 : _GEN_3904; // @[d_cache.scala 171:47]
  wire  _GEN_7495 = _GEN_1030 ? _GEN_3905 : _GEN_3905; // @[d_cache.scala 171:47]
  wire  _GEN_7496 = _GEN_1030 ? _GEN_3906 : _GEN_3906; // @[d_cache.scala 171:47]
  wire  _GEN_7497 = _GEN_1030 ? _GEN_3907 : _GEN_3907; // @[d_cache.scala 171:47]
  wire  _GEN_7498 = _GEN_1030 ? _GEN_3908 : _GEN_3908; // @[d_cache.scala 171:47]
  wire  _GEN_7499 = _GEN_1030 ? _GEN_3909 : _GEN_3909; // @[d_cache.scala 171:47]
  wire  _GEN_7500 = _GEN_1030 ? _GEN_3910 : _GEN_3910; // @[d_cache.scala 171:47]
  wire  _GEN_7501 = _GEN_1030 ? _GEN_3911 : _GEN_3911; // @[d_cache.scala 171:47]
  wire  _GEN_7502 = _GEN_1030 ? _GEN_3912 : _GEN_3912; // @[d_cache.scala 171:47]
  wire  _GEN_7503 = _GEN_1030 ? _GEN_3913 : _GEN_3913; // @[d_cache.scala 171:47]
  wire  _GEN_7504 = _GEN_1030 ? _GEN_3914 : _GEN_3914; // @[d_cache.scala 171:47]
  wire  _GEN_7505 = _GEN_1030 ? _GEN_3915 : _GEN_3915; // @[d_cache.scala 171:47]
  wire  _GEN_7506 = _GEN_1030 ? _GEN_3916 : _GEN_3916; // @[d_cache.scala 171:47]
  wire  _GEN_7507 = _GEN_1030 ? _GEN_3917 : _GEN_3917; // @[d_cache.scala 171:47]
  wire  _GEN_7508 = _GEN_1030 ? _GEN_3918 : _GEN_3918; // @[d_cache.scala 171:47]
  wire  _GEN_7509 = _GEN_1030 ? _GEN_3919 : _GEN_3919; // @[d_cache.scala 171:47]
  wire  _GEN_7510 = _GEN_1030 ? _GEN_3920 : _GEN_3920; // @[d_cache.scala 171:47]
  wire  _GEN_7511 = _GEN_1030 ? _GEN_3921 : _GEN_3921; // @[d_cache.scala 171:47]
  wire  _GEN_7512 = _GEN_1030 ? _GEN_3922 : _GEN_3922; // @[d_cache.scala 171:47]
  wire  _GEN_7513 = _GEN_1030 ? _GEN_3923 : _GEN_3923; // @[d_cache.scala 171:47]
  wire  _GEN_7514 = _GEN_1030 ? _GEN_3924 : _GEN_3924; // @[d_cache.scala 171:47]
  wire  _GEN_7515 = _GEN_1030 ? _GEN_3925 : _GEN_3925; // @[d_cache.scala 171:47]
  wire  _GEN_7516 = _GEN_1030 ? _GEN_3926 : _GEN_3926; // @[d_cache.scala 171:47]
  wire  _GEN_7517 = _GEN_1030 ? _GEN_3927 : _GEN_3927; // @[d_cache.scala 171:47]
  wire  _GEN_7518 = _GEN_1030 ? _GEN_3928 : _GEN_3928; // @[d_cache.scala 171:47]
  wire  _GEN_7519 = _GEN_1030 ? _GEN_3929 : _GEN_3929; // @[d_cache.scala 171:47]
  wire  _GEN_7520 = _GEN_1030 ? _GEN_3930 : _GEN_3930; // @[d_cache.scala 171:47]
  wire  _GEN_7521 = _GEN_1030 ? _GEN_3931 : _GEN_3931; // @[d_cache.scala 171:47]
  wire  _GEN_7522 = _GEN_1030 ? _GEN_3932 : _GEN_3932; // @[d_cache.scala 171:47]
  wire  _GEN_7523 = _GEN_1030 ? _GEN_3933 : _GEN_3933; // @[d_cache.scala 171:47]
  wire  _GEN_7524 = _GEN_1030 ? _GEN_3934 : _GEN_3934; // @[d_cache.scala 171:47]
  wire  _GEN_7525 = _GEN_1030 ? _GEN_3935 : _GEN_3935; // @[d_cache.scala 171:47]
  wire  _GEN_7526 = _GEN_1030 ? _GEN_3936 : _GEN_3936; // @[d_cache.scala 171:47]
  wire  _GEN_7527 = _GEN_1030 ? _GEN_3937 : _GEN_3937; // @[d_cache.scala 171:47]
  wire  _GEN_7528 = _GEN_1030 ? _GEN_3938 : _GEN_3938; // @[d_cache.scala 171:47]
  wire  _GEN_7529 = _GEN_1030 ? _GEN_3939 : _GEN_3939; // @[d_cache.scala 171:47]
  wire  _GEN_7530 = _GEN_1030 ? _GEN_3940 : _GEN_3940; // @[d_cache.scala 171:47]
  wire  _GEN_7531 = _GEN_1030 ? _GEN_3941 : _GEN_3941; // @[d_cache.scala 171:47]
  wire  _GEN_7532 = _GEN_1030 ? _GEN_3942 : _GEN_3942; // @[d_cache.scala 171:47]
  wire  _GEN_7533 = _GEN_1030 ? _GEN_3943 : _GEN_3943; // @[d_cache.scala 171:47]
  wire  _GEN_7534 = _GEN_1030 ? _GEN_3944 : _GEN_3944; // @[d_cache.scala 171:47]
  wire  _GEN_7535 = _GEN_1030 ? _GEN_3945 : _GEN_3945; // @[d_cache.scala 171:47]
  wire  _GEN_7536 = _GEN_1030 ? _GEN_3946 : _GEN_3946; // @[d_cache.scala 171:47]
  wire  _GEN_7537 = _GEN_1030 ? _GEN_3947 : _GEN_3947; // @[d_cache.scala 171:47]
  wire  _GEN_7538 = _GEN_1030 ? _GEN_3948 : _GEN_3948; // @[d_cache.scala 171:47]
  wire  _GEN_7539 = _GEN_1030 ? _GEN_3949 : _GEN_3949; // @[d_cache.scala 171:47]
  wire  _GEN_7540 = _GEN_1030 ? _GEN_3950 : _GEN_3950; // @[d_cache.scala 171:47]
  wire  _GEN_7541 = _GEN_1030 ? _GEN_3951 : _GEN_3951; // @[d_cache.scala 171:47]
  wire  _GEN_7542 = _GEN_1030 ? _GEN_3952 : _GEN_3952; // @[d_cache.scala 171:47]
  wire  _GEN_7543 = _GEN_1030 ? _GEN_3953 : _GEN_3953; // @[d_cache.scala 171:47]
  wire  _GEN_7544 = _GEN_1030 ? _GEN_3954 : _GEN_3954; // @[d_cache.scala 171:47]
  wire  _GEN_7545 = _GEN_1030 ? _GEN_3955 : _GEN_3955; // @[d_cache.scala 171:47]
  wire  _GEN_7546 = _GEN_1030 ? _GEN_3956 : _GEN_3956; // @[d_cache.scala 171:47]
  wire  _GEN_7547 = _GEN_1030 ? _GEN_3957 : _GEN_3957; // @[d_cache.scala 171:47]
  wire  _GEN_7548 = _GEN_1030 ? _GEN_3958 : _GEN_3958; // @[d_cache.scala 171:47]
  wire  _GEN_7549 = _GEN_1030 ? _GEN_3959 : _GEN_3959; // @[d_cache.scala 171:47]
  wire  _GEN_7550 = _GEN_1030 ? _GEN_3960 : _GEN_3960; // @[d_cache.scala 171:47]
  wire  _GEN_7551 = _GEN_1030 ? _GEN_3961 : _GEN_3961; // @[d_cache.scala 171:47]
  wire  _GEN_7552 = _GEN_1030 ? _GEN_3962 : _GEN_3962; // @[d_cache.scala 171:47]
  wire  _GEN_7553 = _GEN_1030 ? _GEN_3963 : _GEN_3963; // @[d_cache.scala 171:47]
  wire  _GEN_7554 = _GEN_1030 ? _GEN_3964 : _GEN_3964; // @[d_cache.scala 171:47]
  wire  _GEN_7555 = _GEN_1030 ? _GEN_3965 : _GEN_3965; // @[d_cache.scala 171:47]
  wire  _GEN_7556 = _GEN_1030 ? _GEN_3966 : _GEN_3966; // @[d_cache.scala 171:47]
  wire  _GEN_7557 = _GEN_1030 ? _GEN_3967 : _GEN_3967; // @[d_cache.scala 171:47]
  wire  _GEN_7558 = _GEN_1030 ? _GEN_3968 : _GEN_3968; // @[d_cache.scala 171:47]
  wire  _GEN_7559 = _GEN_1030 ? _GEN_3969 : _GEN_3969; // @[d_cache.scala 171:47]
  wire  _GEN_7560 = _GEN_1030 ? _GEN_3970 : _GEN_3970; // @[d_cache.scala 171:47]
  wire  _GEN_7561 = _GEN_1030 ? _GEN_3971 : _GEN_3971; // @[d_cache.scala 171:47]
  wire  _GEN_7562 = _GEN_1030 ? _GEN_3972 : _GEN_3972; // @[d_cache.scala 171:47]
  wire  _GEN_7563 = _GEN_1030 ? _GEN_3973 : _GEN_3973; // @[d_cache.scala 171:47]
  wire  _GEN_7564 = _GEN_1030 ? _GEN_3974 : _GEN_3974; // @[d_cache.scala 171:47]
  wire  _GEN_7565 = _GEN_1030 ? _GEN_3975 : _GEN_3975; // @[d_cache.scala 171:47]
  wire  _GEN_7566 = _GEN_1030 ? _GEN_3976 : _GEN_3976; // @[d_cache.scala 171:47]
  wire  _GEN_7567 = _GEN_1030 ? _GEN_3977 : _GEN_3977; // @[d_cache.scala 171:47]
  wire  _GEN_7568 = _GEN_1030 ? _GEN_3978 : _GEN_3978; // @[d_cache.scala 171:47]
  wire  _GEN_7569 = _GEN_1030 ? _GEN_3979 : _GEN_3979; // @[d_cache.scala 171:47]
  wire  _GEN_7570 = _GEN_1030 ? _GEN_3980 : _GEN_3980; // @[d_cache.scala 171:47]
  wire  _GEN_7571 = _GEN_1030 ? _GEN_3981 : _GEN_3981; // @[d_cache.scala 171:47]
  wire [2:0] _GEN_7572 = _GEN_1030 ? 3'h6 : 3'h7; // @[d_cache.scala 171:47 178:31 181:31]
  wire [63:0] _GEN_7574 = ~quene ? _GEN_5262 : _GEN_7058; // @[d_cache.scala 152:34]
  wire [41:0] _GEN_7575 = ~quene ? _GEN_5263 : _GEN_7059; // @[d_cache.scala 152:34]
  wire [63:0] _GEN_7576 = ~quene ? _GEN_5264 : ram_0_0; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7577 = ~quene ? _GEN_5265 : ram_0_1; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7578 = ~quene ? _GEN_5266 : ram_0_2; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7579 = ~quene ? _GEN_5267 : ram_0_3; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7580 = ~quene ? _GEN_5268 : ram_0_4; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7581 = ~quene ? _GEN_5269 : ram_0_5; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7582 = ~quene ? _GEN_5270 : ram_0_6; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7583 = ~quene ? _GEN_5271 : ram_0_7; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7584 = ~quene ? _GEN_5272 : ram_0_8; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7585 = ~quene ? _GEN_5273 : ram_0_9; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7586 = ~quene ? _GEN_5274 : ram_0_10; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7587 = ~quene ? _GEN_5275 : ram_0_11; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7588 = ~quene ? _GEN_5276 : ram_0_12; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7589 = ~quene ? _GEN_5277 : ram_0_13; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7590 = ~quene ? _GEN_5278 : ram_0_14; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7591 = ~quene ? _GEN_5279 : ram_0_15; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7592 = ~quene ? _GEN_5280 : ram_0_16; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7593 = ~quene ? _GEN_5281 : ram_0_17; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7594 = ~quene ? _GEN_5282 : ram_0_18; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7595 = ~quene ? _GEN_5283 : ram_0_19; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7596 = ~quene ? _GEN_5284 : ram_0_20; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7597 = ~quene ? _GEN_5285 : ram_0_21; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7598 = ~quene ? _GEN_5286 : ram_0_22; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7599 = ~quene ? _GEN_5287 : ram_0_23; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7600 = ~quene ? _GEN_5288 : ram_0_24; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7601 = ~quene ? _GEN_5289 : ram_0_25; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7602 = ~quene ? _GEN_5290 : ram_0_26; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7603 = ~quene ? _GEN_5291 : ram_0_27; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7604 = ~quene ? _GEN_5292 : ram_0_28; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7605 = ~quene ? _GEN_5293 : ram_0_29; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7606 = ~quene ? _GEN_5294 : ram_0_30; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7607 = ~quene ? _GEN_5295 : ram_0_31; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7608 = ~quene ? _GEN_5296 : ram_0_32; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7609 = ~quene ? _GEN_5297 : ram_0_33; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7610 = ~quene ? _GEN_5298 : ram_0_34; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7611 = ~quene ? _GEN_5299 : ram_0_35; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7612 = ~quene ? _GEN_5300 : ram_0_36; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7613 = ~quene ? _GEN_5301 : ram_0_37; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7614 = ~quene ? _GEN_5302 : ram_0_38; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7615 = ~quene ? _GEN_5303 : ram_0_39; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7616 = ~quene ? _GEN_5304 : ram_0_40; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7617 = ~quene ? _GEN_5305 : ram_0_41; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7618 = ~quene ? _GEN_5306 : ram_0_42; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7619 = ~quene ? _GEN_5307 : ram_0_43; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7620 = ~quene ? _GEN_5308 : ram_0_44; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7621 = ~quene ? _GEN_5309 : ram_0_45; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7622 = ~quene ? _GEN_5310 : ram_0_46; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7623 = ~quene ? _GEN_5311 : ram_0_47; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7624 = ~quene ? _GEN_5312 : ram_0_48; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7625 = ~quene ? _GEN_5313 : ram_0_49; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7626 = ~quene ? _GEN_5314 : ram_0_50; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7627 = ~quene ? _GEN_5315 : ram_0_51; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7628 = ~quene ? _GEN_5316 : ram_0_52; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7629 = ~quene ? _GEN_5317 : ram_0_53; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7630 = ~quene ? _GEN_5318 : ram_0_54; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7631 = ~quene ? _GEN_5319 : ram_0_55; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7632 = ~quene ? _GEN_5320 : ram_0_56; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7633 = ~quene ? _GEN_5321 : ram_0_57; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7634 = ~quene ? _GEN_5322 : ram_0_58; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7635 = ~quene ? _GEN_5323 : ram_0_59; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7636 = ~quene ? _GEN_5324 : ram_0_60; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7637 = ~quene ? _GEN_5325 : ram_0_61; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7638 = ~quene ? _GEN_5326 : ram_0_62; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7639 = ~quene ? _GEN_5327 : ram_0_63; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7640 = ~quene ? _GEN_5328 : ram_0_64; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7641 = ~quene ? _GEN_5329 : ram_0_65; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7642 = ~quene ? _GEN_5330 : ram_0_66; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7643 = ~quene ? _GEN_5331 : ram_0_67; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7644 = ~quene ? _GEN_5332 : ram_0_68; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7645 = ~quene ? _GEN_5333 : ram_0_69; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7646 = ~quene ? _GEN_5334 : ram_0_70; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7647 = ~quene ? _GEN_5335 : ram_0_71; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7648 = ~quene ? _GEN_5336 : ram_0_72; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7649 = ~quene ? _GEN_5337 : ram_0_73; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7650 = ~quene ? _GEN_5338 : ram_0_74; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7651 = ~quene ? _GEN_5339 : ram_0_75; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7652 = ~quene ? _GEN_5340 : ram_0_76; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7653 = ~quene ? _GEN_5341 : ram_0_77; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7654 = ~quene ? _GEN_5342 : ram_0_78; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7655 = ~quene ? _GEN_5343 : ram_0_79; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7656 = ~quene ? _GEN_5344 : ram_0_80; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7657 = ~quene ? _GEN_5345 : ram_0_81; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7658 = ~quene ? _GEN_5346 : ram_0_82; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7659 = ~quene ? _GEN_5347 : ram_0_83; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7660 = ~quene ? _GEN_5348 : ram_0_84; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7661 = ~quene ? _GEN_5349 : ram_0_85; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7662 = ~quene ? _GEN_5350 : ram_0_86; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7663 = ~quene ? _GEN_5351 : ram_0_87; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7664 = ~quene ? _GEN_5352 : ram_0_88; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7665 = ~quene ? _GEN_5353 : ram_0_89; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7666 = ~quene ? _GEN_5354 : ram_0_90; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7667 = ~quene ? _GEN_5355 : ram_0_91; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7668 = ~quene ? _GEN_5356 : ram_0_92; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7669 = ~quene ? _GEN_5357 : ram_0_93; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7670 = ~quene ? _GEN_5358 : ram_0_94; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7671 = ~quene ? _GEN_5359 : ram_0_95; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7672 = ~quene ? _GEN_5360 : ram_0_96; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7673 = ~quene ? _GEN_5361 : ram_0_97; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7674 = ~quene ? _GEN_5362 : ram_0_98; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7675 = ~quene ? _GEN_5363 : ram_0_99; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7676 = ~quene ? _GEN_5364 : ram_0_100; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7677 = ~quene ? _GEN_5365 : ram_0_101; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7678 = ~quene ? _GEN_5366 : ram_0_102; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7679 = ~quene ? _GEN_5367 : ram_0_103; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7680 = ~quene ? _GEN_5368 : ram_0_104; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7681 = ~quene ? _GEN_5369 : ram_0_105; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7682 = ~quene ? _GEN_5370 : ram_0_106; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7683 = ~quene ? _GEN_5371 : ram_0_107; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7684 = ~quene ? _GEN_5372 : ram_0_108; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7685 = ~quene ? _GEN_5373 : ram_0_109; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7686 = ~quene ? _GEN_5374 : ram_0_110; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7687 = ~quene ? _GEN_5375 : ram_0_111; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7688 = ~quene ? _GEN_5376 : ram_0_112; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7689 = ~quene ? _GEN_5377 : ram_0_113; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7690 = ~quene ? _GEN_5378 : ram_0_114; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7691 = ~quene ? _GEN_5379 : ram_0_115; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7692 = ~quene ? _GEN_5380 : ram_0_116; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7693 = ~quene ? _GEN_5381 : ram_0_117; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7694 = ~quene ? _GEN_5382 : ram_0_118; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7695 = ~quene ? _GEN_5383 : ram_0_119; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7696 = ~quene ? _GEN_5384 : ram_0_120; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7697 = ~quene ? _GEN_5385 : ram_0_121; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7698 = ~quene ? _GEN_5386 : ram_0_122; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7699 = ~quene ? _GEN_5387 : ram_0_123; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7700 = ~quene ? _GEN_5388 : ram_0_124; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7701 = ~quene ? _GEN_5389 : ram_0_125; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7702 = ~quene ? _GEN_5390 : ram_0_126; // @[d_cache.scala 152:34 18:24]
  wire [63:0] _GEN_7703 = ~quene ? _GEN_5391 : ram_0_127; // @[d_cache.scala 152:34 18:24]
  wire [31:0] _GEN_7704 = ~quene ? _GEN_5392 : tag_0_0; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7705 = ~quene ? _GEN_5393 : tag_0_1; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7706 = ~quene ? _GEN_5394 : tag_0_2; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7707 = ~quene ? _GEN_5395 : tag_0_3; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7708 = ~quene ? _GEN_5396 : tag_0_4; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7709 = ~quene ? _GEN_5397 : tag_0_5; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7710 = ~quene ? _GEN_5398 : tag_0_6; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7711 = ~quene ? _GEN_5399 : tag_0_7; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7712 = ~quene ? _GEN_5400 : tag_0_8; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7713 = ~quene ? _GEN_5401 : tag_0_9; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7714 = ~quene ? _GEN_5402 : tag_0_10; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7715 = ~quene ? _GEN_5403 : tag_0_11; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7716 = ~quene ? _GEN_5404 : tag_0_12; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7717 = ~quene ? _GEN_5405 : tag_0_13; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7718 = ~quene ? _GEN_5406 : tag_0_14; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7719 = ~quene ? _GEN_5407 : tag_0_15; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7720 = ~quene ? _GEN_5408 : tag_0_16; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7721 = ~quene ? _GEN_5409 : tag_0_17; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7722 = ~quene ? _GEN_5410 : tag_0_18; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7723 = ~quene ? _GEN_5411 : tag_0_19; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7724 = ~quene ? _GEN_5412 : tag_0_20; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7725 = ~quene ? _GEN_5413 : tag_0_21; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7726 = ~quene ? _GEN_5414 : tag_0_22; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7727 = ~quene ? _GEN_5415 : tag_0_23; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7728 = ~quene ? _GEN_5416 : tag_0_24; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7729 = ~quene ? _GEN_5417 : tag_0_25; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7730 = ~quene ? _GEN_5418 : tag_0_26; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7731 = ~quene ? _GEN_5419 : tag_0_27; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7732 = ~quene ? _GEN_5420 : tag_0_28; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7733 = ~quene ? _GEN_5421 : tag_0_29; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7734 = ~quene ? _GEN_5422 : tag_0_30; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7735 = ~quene ? _GEN_5423 : tag_0_31; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7736 = ~quene ? _GEN_5424 : tag_0_32; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7737 = ~quene ? _GEN_5425 : tag_0_33; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7738 = ~quene ? _GEN_5426 : tag_0_34; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7739 = ~quene ? _GEN_5427 : tag_0_35; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7740 = ~quene ? _GEN_5428 : tag_0_36; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7741 = ~quene ? _GEN_5429 : tag_0_37; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7742 = ~quene ? _GEN_5430 : tag_0_38; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7743 = ~quene ? _GEN_5431 : tag_0_39; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7744 = ~quene ? _GEN_5432 : tag_0_40; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7745 = ~quene ? _GEN_5433 : tag_0_41; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7746 = ~quene ? _GEN_5434 : tag_0_42; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7747 = ~quene ? _GEN_5435 : tag_0_43; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7748 = ~quene ? _GEN_5436 : tag_0_44; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7749 = ~quene ? _GEN_5437 : tag_0_45; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7750 = ~quene ? _GEN_5438 : tag_0_46; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7751 = ~quene ? _GEN_5439 : tag_0_47; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7752 = ~quene ? _GEN_5440 : tag_0_48; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7753 = ~quene ? _GEN_5441 : tag_0_49; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7754 = ~quene ? _GEN_5442 : tag_0_50; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7755 = ~quene ? _GEN_5443 : tag_0_51; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7756 = ~quene ? _GEN_5444 : tag_0_52; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7757 = ~quene ? _GEN_5445 : tag_0_53; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7758 = ~quene ? _GEN_5446 : tag_0_54; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7759 = ~quene ? _GEN_5447 : tag_0_55; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7760 = ~quene ? _GEN_5448 : tag_0_56; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7761 = ~quene ? _GEN_5449 : tag_0_57; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7762 = ~quene ? _GEN_5450 : tag_0_58; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7763 = ~quene ? _GEN_5451 : tag_0_59; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7764 = ~quene ? _GEN_5452 : tag_0_60; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7765 = ~quene ? _GEN_5453 : tag_0_61; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7766 = ~quene ? _GEN_5454 : tag_0_62; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7767 = ~quene ? _GEN_5455 : tag_0_63; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7768 = ~quene ? _GEN_5456 : tag_0_64; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7769 = ~quene ? _GEN_5457 : tag_0_65; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7770 = ~quene ? _GEN_5458 : tag_0_66; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7771 = ~quene ? _GEN_5459 : tag_0_67; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7772 = ~quene ? _GEN_5460 : tag_0_68; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7773 = ~quene ? _GEN_5461 : tag_0_69; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7774 = ~quene ? _GEN_5462 : tag_0_70; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7775 = ~quene ? _GEN_5463 : tag_0_71; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7776 = ~quene ? _GEN_5464 : tag_0_72; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7777 = ~quene ? _GEN_5465 : tag_0_73; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7778 = ~quene ? _GEN_5466 : tag_0_74; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7779 = ~quene ? _GEN_5467 : tag_0_75; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7780 = ~quene ? _GEN_5468 : tag_0_76; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7781 = ~quene ? _GEN_5469 : tag_0_77; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7782 = ~quene ? _GEN_5470 : tag_0_78; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7783 = ~quene ? _GEN_5471 : tag_0_79; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7784 = ~quene ? _GEN_5472 : tag_0_80; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7785 = ~quene ? _GEN_5473 : tag_0_81; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7786 = ~quene ? _GEN_5474 : tag_0_82; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7787 = ~quene ? _GEN_5475 : tag_0_83; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7788 = ~quene ? _GEN_5476 : tag_0_84; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7789 = ~quene ? _GEN_5477 : tag_0_85; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7790 = ~quene ? _GEN_5478 : tag_0_86; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7791 = ~quene ? _GEN_5479 : tag_0_87; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7792 = ~quene ? _GEN_5480 : tag_0_88; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7793 = ~quene ? _GEN_5481 : tag_0_89; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7794 = ~quene ? _GEN_5482 : tag_0_90; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7795 = ~quene ? _GEN_5483 : tag_0_91; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7796 = ~quene ? _GEN_5484 : tag_0_92; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7797 = ~quene ? _GEN_5485 : tag_0_93; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7798 = ~quene ? _GEN_5486 : tag_0_94; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7799 = ~quene ? _GEN_5487 : tag_0_95; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7800 = ~quene ? _GEN_5488 : tag_0_96; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7801 = ~quene ? _GEN_5489 : tag_0_97; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7802 = ~quene ? _GEN_5490 : tag_0_98; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7803 = ~quene ? _GEN_5491 : tag_0_99; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7804 = ~quene ? _GEN_5492 : tag_0_100; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7805 = ~quene ? _GEN_5493 : tag_0_101; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7806 = ~quene ? _GEN_5494 : tag_0_102; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7807 = ~quene ? _GEN_5495 : tag_0_103; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7808 = ~quene ? _GEN_5496 : tag_0_104; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7809 = ~quene ? _GEN_5497 : tag_0_105; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7810 = ~quene ? _GEN_5498 : tag_0_106; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7811 = ~quene ? _GEN_5499 : tag_0_107; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7812 = ~quene ? _GEN_5500 : tag_0_108; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7813 = ~quene ? _GEN_5501 : tag_0_109; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7814 = ~quene ? _GEN_5502 : tag_0_110; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7815 = ~quene ? _GEN_5503 : tag_0_111; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7816 = ~quene ? _GEN_5504 : tag_0_112; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7817 = ~quene ? _GEN_5505 : tag_0_113; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7818 = ~quene ? _GEN_5506 : tag_0_114; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7819 = ~quene ? _GEN_5507 : tag_0_115; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7820 = ~quene ? _GEN_5508 : tag_0_116; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7821 = ~quene ? _GEN_5509 : tag_0_117; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7822 = ~quene ? _GEN_5510 : tag_0_118; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7823 = ~quene ? _GEN_5511 : tag_0_119; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7824 = ~quene ? _GEN_5512 : tag_0_120; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7825 = ~quene ? _GEN_5513 : tag_0_121; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7826 = ~quene ? _GEN_5514 : tag_0_122; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7827 = ~quene ? _GEN_5515 : tag_0_123; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7828 = ~quene ? _GEN_5516 : tag_0_124; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7829 = ~quene ? _GEN_5517 : tag_0_125; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7830 = ~quene ? _GEN_5518 : tag_0_126; // @[d_cache.scala 152:34 22:24]
  wire [31:0] _GEN_7831 = ~quene ? _GEN_5519 : tag_0_127; // @[d_cache.scala 152:34 22:24]
  wire  _GEN_7832 = ~quene ? _GEN_5520 : dirty_0_0; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7833 = ~quene ? _GEN_5521 : dirty_0_1; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7834 = ~quene ? _GEN_5522 : dirty_0_2; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7835 = ~quene ? _GEN_5523 : dirty_0_3; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7836 = ~quene ? _GEN_5524 : dirty_0_4; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7837 = ~quene ? _GEN_5525 : dirty_0_5; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7838 = ~quene ? _GEN_5526 : dirty_0_6; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7839 = ~quene ? _GEN_5527 : dirty_0_7; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7840 = ~quene ? _GEN_5528 : dirty_0_8; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7841 = ~quene ? _GEN_5529 : dirty_0_9; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7842 = ~quene ? _GEN_5530 : dirty_0_10; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7843 = ~quene ? _GEN_5531 : dirty_0_11; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7844 = ~quene ? _GEN_5532 : dirty_0_12; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7845 = ~quene ? _GEN_5533 : dirty_0_13; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7846 = ~quene ? _GEN_5534 : dirty_0_14; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7847 = ~quene ? _GEN_5535 : dirty_0_15; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7848 = ~quene ? _GEN_5536 : dirty_0_16; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7849 = ~quene ? _GEN_5537 : dirty_0_17; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7850 = ~quene ? _GEN_5538 : dirty_0_18; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7851 = ~quene ? _GEN_5539 : dirty_0_19; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7852 = ~quene ? _GEN_5540 : dirty_0_20; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7853 = ~quene ? _GEN_5541 : dirty_0_21; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7854 = ~quene ? _GEN_5542 : dirty_0_22; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7855 = ~quene ? _GEN_5543 : dirty_0_23; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7856 = ~quene ? _GEN_5544 : dirty_0_24; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7857 = ~quene ? _GEN_5545 : dirty_0_25; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7858 = ~quene ? _GEN_5546 : dirty_0_26; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7859 = ~quene ? _GEN_5547 : dirty_0_27; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7860 = ~quene ? _GEN_5548 : dirty_0_28; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7861 = ~quene ? _GEN_5549 : dirty_0_29; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7862 = ~quene ? _GEN_5550 : dirty_0_30; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7863 = ~quene ? _GEN_5551 : dirty_0_31; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7864 = ~quene ? _GEN_5552 : dirty_0_32; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7865 = ~quene ? _GEN_5553 : dirty_0_33; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7866 = ~quene ? _GEN_5554 : dirty_0_34; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7867 = ~quene ? _GEN_5555 : dirty_0_35; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7868 = ~quene ? _GEN_5556 : dirty_0_36; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7869 = ~quene ? _GEN_5557 : dirty_0_37; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7870 = ~quene ? _GEN_5558 : dirty_0_38; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7871 = ~quene ? _GEN_5559 : dirty_0_39; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7872 = ~quene ? _GEN_5560 : dirty_0_40; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7873 = ~quene ? _GEN_5561 : dirty_0_41; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7874 = ~quene ? _GEN_5562 : dirty_0_42; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7875 = ~quene ? _GEN_5563 : dirty_0_43; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7876 = ~quene ? _GEN_5564 : dirty_0_44; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7877 = ~quene ? _GEN_5565 : dirty_0_45; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7878 = ~quene ? _GEN_5566 : dirty_0_46; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7879 = ~quene ? _GEN_5567 : dirty_0_47; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7880 = ~quene ? _GEN_5568 : dirty_0_48; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7881 = ~quene ? _GEN_5569 : dirty_0_49; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7882 = ~quene ? _GEN_5570 : dirty_0_50; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7883 = ~quene ? _GEN_5571 : dirty_0_51; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7884 = ~quene ? _GEN_5572 : dirty_0_52; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7885 = ~quene ? _GEN_5573 : dirty_0_53; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7886 = ~quene ? _GEN_5574 : dirty_0_54; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7887 = ~quene ? _GEN_5575 : dirty_0_55; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7888 = ~quene ? _GEN_5576 : dirty_0_56; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7889 = ~quene ? _GEN_5577 : dirty_0_57; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7890 = ~quene ? _GEN_5578 : dirty_0_58; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7891 = ~quene ? _GEN_5579 : dirty_0_59; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7892 = ~quene ? _GEN_5580 : dirty_0_60; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7893 = ~quene ? _GEN_5581 : dirty_0_61; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7894 = ~quene ? _GEN_5582 : dirty_0_62; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7895 = ~quene ? _GEN_5583 : dirty_0_63; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7896 = ~quene ? _GEN_5584 : dirty_0_64; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7897 = ~quene ? _GEN_5585 : dirty_0_65; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7898 = ~quene ? _GEN_5586 : dirty_0_66; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7899 = ~quene ? _GEN_5587 : dirty_0_67; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7900 = ~quene ? _GEN_5588 : dirty_0_68; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7901 = ~quene ? _GEN_5589 : dirty_0_69; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7902 = ~quene ? _GEN_5590 : dirty_0_70; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7903 = ~quene ? _GEN_5591 : dirty_0_71; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7904 = ~quene ? _GEN_5592 : dirty_0_72; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7905 = ~quene ? _GEN_5593 : dirty_0_73; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7906 = ~quene ? _GEN_5594 : dirty_0_74; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7907 = ~quene ? _GEN_5595 : dirty_0_75; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7908 = ~quene ? _GEN_5596 : dirty_0_76; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7909 = ~quene ? _GEN_5597 : dirty_0_77; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7910 = ~quene ? _GEN_5598 : dirty_0_78; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7911 = ~quene ? _GEN_5599 : dirty_0_79; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7912 = ~quene ? _GEN_5600 : dirty_0_80; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7913 = ~quene ? _GEN_5601 : dirty_0_81; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7914 = ~quene ? _GEN_5602 : dirty_0_82; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7915 = ~quene ? _GEN_5603 : dirty_0_83; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7916 = ~quene ? _GEN_5604 : dirty_0_84; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7917 = ~quene ? _GEN_5605 : dirty_0_85; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7918 = ~quene ? _GEN_5606 : dirty_0_86; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7919 = ~quene ? _GEN_5607 : dirty_0_87; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7920 = ~quene ? _GEN_5608 : dirty_0_88; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7921 = ~quene ? _GEN_5609 : dirty_0_89; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7922 = ~quene ? _GEN_5610 : dirty_0_90; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7923 = ~quene ? _GEN_5611 : dirty_0_91; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7924 = ~quene ? _GEN_5612 : dirty_0_92; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7925 = ~quene ? _GEN_5613 : dirty_0_93; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7926 = ~quene ? _GEN_5614 : dirty_0_94; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7927 = ~quene ? _GEN_5615 : dirty_0_95; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7928 = ~quene ? _GEN_5616 : dirty_0_96; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7929 = ~quene ? _GEN_5617 : dirty_0_97; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7930 = ~quene ? _GEN_5618 : dirty_0_98; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7931 = ~quene ? _GEN_5619 : dirty_0_99; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7932 = ~quene ? _GEN_5620 : dirty_0_100; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7933 = ~quene ? _GEN_5621 : dirty_0_101; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7934 = ~quene ? _GEN_5622 : dirty_0_102; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7935 = ~quene ? _GEN_5623 : dirty_0_103; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7936 = ~quene ? _GEN_5624 : dirty_0_104; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7937 = ~quene ? _GEN_5625 : dirty_0_105; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7938 = ~quene ? _GEN_5626 : dirty_0_106; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7939 = ~quene ? _GEN_5627 : dirty_0_107; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7940 = ~quene ? _GEN_5628 : dirty_0_108; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7941 = ~quene ? _GEN_5629 : dirty_0_109; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7942 = ~quene ? _GEN_5630 : dirty_0_110; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7943 = ~quene ? _GEN_5631 : dirty_0_111; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7944 = ~quene ? _GEN_5632 : dirty_0_112; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7945 = ~quene ? _GEN_5633 : dirty_0_113; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7946 = ~quene ? _GEN_5634 : dirty_0_114; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7947 = ~quene ? _GEN_5635 : dirty_0_115; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7948 = ~quene ? _GEN_5636 : dirty_0_116; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7949 = ~quene ? _GEN_5637 : dirty_0_117; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7950 = ~quene ? _GEN_5638 : dirty_0_118; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7951 = ~quene ? _GEN_5639 : dirty_0_119; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7952 = ~quene ? _GEN_5640 : dirty_0_120; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7953 = ~quene ? _GEN_5641 : dirty_0_121; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7954 = ~quene ? _GEN_5642 : dirty_0_122; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7955 = ~quene ? _GEN_5643 : dirty_0_123; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7956 = ~quene ? _GEN_5644 : dirty_0_124; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7957 = ~quene ? _GEN_5645 : dirty_0_125; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7958 = ~quene ? _GEN_5646 : dirty_0_126; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7959 = ~quene ? _GEN_5647 : dirty_0_127; // @[d_cache.scala 152:34 26:26]
  wire  _GEN_7960 = ~quene ? _GEN_5648 : valid_0_0; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7961 = ~quene ? _GEN_5649 : valid_0_1; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7962 = ~quene ? _GEN_5650 : valid_0_2; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7963 = ~quene ? _GEN_5651 : valid_0_3; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7964 = ~quene ? _GEN_5652 : valid_0_4; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7965 = ~quene ? _GEN_5653 : valid_0_5; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7966 = ~quene ? _GEN_5654 : valid_0_6; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7967 = ~quene ? _GEN_5655 : valid_0_7; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7968 = ~quene ? _GEN_5656 : valid_0_8; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7969 = ~quene ? _GEN_5657 : valid_0_9; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7970 = ~quene ? _GEN_5658 : valid_0_10; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7971 = ~quene ? _GEN_5659 : valid_0_11; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7972 = ~quene ? _GEN_5660 : valid_0_12; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7973 = ~quene ? _GEN_5661 : valid_0_13; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7974 = ~quene ? _GEN_5662 : valid_0_14; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7975 = ~quene ? _GEN_5663 : valid_0_15; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7976 = ~quene ? _GEN_5664 : valid_0_16; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7977 = ~quene ? _GEN_5665 : valid_0_17; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7978 = ~quene ? _GEN_5666 : valid_0_18; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7979 = ~quene ? _GEN_5667 : valid_0_19; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7980 = ~quene ? _GEN_5668 : valid_0_20; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7981 = ~quene ? _GEN_5669 : valid_0_21; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7982 = ~quene ? _GEN_5670 : valid_0_22; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7983 = ~quene ? _GEN_5671 : valid_0_23; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7984 = ~quene ? _GEN_5672 : valid_0_24; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7985 = ~quene ? _GEN_5673 : valid_0_25; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7986 = ~quene ? _GEN_5674 : valid_0_26; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7987 = ~quene ? _GEN_5675 : valid_0_27; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7988 = ~quene ? _GEN_5676 : valid_0_28; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7989 = ~quene ? _GEN_5677 : valid_0_29; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7990 = ~quene ? _GEN_5678 : valid_0_30; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7991 = ~quene ? _GEN_5679 : valid_0_31; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7992 = ~quene ? _GEN_5680 : valid_0_32; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7993 = ~quene ? _GEN_5681 : valid_0_33; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7994 = ~quene ? _GEN_5682 : valid_0_34; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7995 = ~quene ? _GEN_5683 : valid_0_35; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7996 = ~quene ? _GEN_5684 : valid_0_36; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7997 = ~quene ? _GEN_5685 : valid_0_37; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7998 = ~quene ? _GEN_5686 : valid_0_38; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_7999 = ~quene ? _GEN_5687 : valid_0_39; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8000 = ~quene ? _GEN_5688 : valid_0_40; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8001 = ~quene ? _GEN_5689 : valid_0_41; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8002 = ~quene ? _GEN_5690 : valid_0_42; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8003 = ~quene ? _GEN_5691 : valid_0_43; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8004 = ~quene ? _GEN_5692 : valid_0_44; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8005 = ~quene ? _GEN_5693 : valid_0_45; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8006 = ~quene ? _GEN_5694 : valid_0_46; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8007 = ~quene ? _GEN_5695 : valid_0_47; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8008 = ~quene ? _GEN_5696 : valid_0_48; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8009 = ~quene ? _GEN_5697 : valid_0_49; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8010 = ~quene ? _GEN_5698 : valid_0_50; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8011 = ~quene ? _GEN_5699 : valid_0_51; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8012 = ~quene ? _GEN_5700 : valid_0_52; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8013 = ~quene ? _GEN_5701 : valid_0_53; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8014 = ~quene ? _GEN_5702 : valid_0_54; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8015 = ~quene ? _GEN_5703 : valid_0_55; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8016 = ~quene ? _GEN_5704 : valid_0_56; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8017 = ~quene ? _GEN_5705 : valid_0_57; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8018 = ~quene ? _GEN_5706 : valid_0_58; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8019 = ~quene ? _GEN_5707 : valid_0_59; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8020 = ~quene ? _GEN_5708 : valid_0_60; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8021 = ~quene ? _GEN_5709 : valid_0_61; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8022 = ~quene ? _GEN_5710 : valid_0_62; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8023 = ~quene ? _GEN_5711 : valid_0_63; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8024 = ~quene ? _GEN_5712 : valid_0_64; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8025 = ~quene ? _GEN_5713 : valid_0_65; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8026 = ~quene ? _GEN_5714 : valid_0_66; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8027 = ~quene ? _GEN_5715 : valid_0_67; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8028 = ~quene ? _GEN_5716 : valid_0_68; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8029 = ~quene ? _GEN_5717 : valid_0_69; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8030 = ~quene ? _GEN_5718 : valid_0_70; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8031 = ~quene ? _GEN_5719 : valid_0_71; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8032 = ~quene ? _GEN_5720 : valid_0_72; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8033 = ~quene ? _GEN_5721 : valid_0_73; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8034 = ~quene ? _GEN_5722 : valid_0_74; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8035 = ~quene ? _GEN_5723 : valid_0_75; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8036 = ~quene ? _GEN_5724 : valid_0_76; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8037 = ~quene ? _GEN_5725 : valid_0_77; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8038 = ~quene ? _GEN_5726 : valid_0_78; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8039 = ~quene ? _GEN_5727 : valid_0_79; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8040 = ~quene ? _GEN_5728 : valid_0_80; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8041 = ~quene ? _GEN_5729 : valid_0_81; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8042 = ~quene ? _GEN_5730 : valid_0_82; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8043 = ~quene ? _GEN_5731 : valid_0_83; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8044 = ~quene ? _GEN_5732 : valid_0_84; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8045 = ~quene ? _GEN_5733 : valid_0_85; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8046 = ~quene ? _GEN_5734 : valid_0_86; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8047 = ~quene ? _GEN_5735 : valid_0_87; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8048 = ~quene ? _GEN_5736 : valid_0_88; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8049 = ~quene ? _GEN_5737 : valid_0_89; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8050 = ~quene ? _GEN_5738 : valid_0_90; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8051 = ~quene ? _GEN_5739 : valid_0_91; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8052 = ~quene ? _GEN_5740 : valid_0_92; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8053 = ~quene ? _GEN_5741 : valid_0_93; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8054 = ~quene ? _GEN_5742 : valid_0_94; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8055 = ~quene ? _GEN_5743 : valid_0_95; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8056 = ~quene ? _GEN_5744 : valid_0_96; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8057 = ~quene ? _GEN_5745 : valid_0_97; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8058 = ~quene ? _GEN_5746 : valid_0_98; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8059 = ~quene ? _GEN_5747 : valid_0_99; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8060 = ~quene ? _GEN_5748 : valid_0_100; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8061 = ~quene ? _GEN_5749 : valid_0_101; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8062 = ~quene ? _GEN_5750 : valid_0_102; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8063 = ~quene ? _GEN_5751 : valid_0_103; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8064 = ~quene ? _GEN_5752 : valid_0_104; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8065 = ~quene ? _GEN_5753 : valid_0_105; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8066 = ~quene ? _GEN_5754 : valid_0_106; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8067 = ~quene ? _GEN_5755 : valid_0_107; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8068 = ~quene ? _GEN_5756 : valid_0_108; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8069 = ~quene ? _GEN_5757 : valid_0_109; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8070 = ~quene ? _GEN_5758 : valid_0_110; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8071 = ~quene ? _GEN_5759 : valid_0_111; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8072 = ~quene ? _GEN_5760 : valid_0_112; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8073 = ~quene ? _GEN_5761 : valid_0_113; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8074 = ~quene ? _GEN_5762 : valid_0_114; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8075 = ~quene ? _GEN_5763 : valid_0_115; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8076 = ~quene ? _GEN_5764 : valid_0_116; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8077 = ~quene ? _GEN_5765 : valid_0_117; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8078 = ~quene ? _GEN_5766 : valid_0_118; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8079 = ~quene ? _GEN_5767 : valid_0_119; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8080 = ~quene ? _GEN_5768 : valid_0_120; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8081 = ~quene ? _GEN_5769 : valid_0_121; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8082 = ~quene ? _GEN_5770 : valid_0_122; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8083 = ~quene ? _GEN_5771 : valid_0_123; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8084 = ~quene ? _GEN_5772 : valid_0_124; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8085 = ~quene ? _GEN_5773 : valid_0_125; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8086 = ~quene ? _GEN_5774 : valid_0_126; // @[d_cache.scala 152:34 24:26]
  wire  _GEN_8087 = ~quene ? _GEN_5775 : valid_0_127; // @[d_cache.scala 152:34 24:26]
  wire [2:0] _GEN_8088 = ~quene ? _GEN_5776 : _GEN_7572; // @[d_cache.scala 152:34]
  wire [63:0] _GEN_8090 = ~quene ? ram_1_0 : _GEN_7060; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8091 = ~quene ? ram_1_1 : _GEN_7061; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8092 = ~quene ? ram_1_2 : _GEN_7062; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8093 = ~quene ? ram_1_3 : _GEN_7063; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8094 = ~quene ? ram_1_4 : _GEN_7064; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8095 = ~quene ? ram_1_5 : _GEN_7065; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8096 = ~quene ? ram_1_6 : _GEN_7066; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8097 = ~quene ? ram_1_7 : _GEN_7067; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8098 = ~quene ? ram_1_8 : _GEN_7068; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8099 = ~quene ? ram_1_9 : _GEN_7069; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8100 = ~quene ? ram_1_10 : _GEN_7070; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8101 = ~quene ? ram_1_11 : _GEN_7071; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8102 = ~quene ? ram_1_12 : _GEN_7072; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8103 = ~quene ? ram_1_13 : _GEN_7073; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8104 = ~quene ? ram_1_14 : _GEN_7074; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8105 = ~quene ? ram_1_15 : _GEN_7075; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8106 = ~quene ? ram_1_16 : _GEN_7076; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8107 = ~quene ? ram_1_17 : _GEN_7077; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8108 = ~quene ? ram_1_18 : _GEN_7078; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8109 = ~quene ? ram_1_19 : _GEN_7079; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8110 = ~quene ? ram_1_20 : _GEN_7080; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8111 = ~quene ? ram_1_21 : _GEN_7081; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8112 = ~quene ? ram_1_22 : _GEN_7082; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8113 = ~quene ? ram_1_23 : _GEN_7083; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8114 = ~quene ? ram_1_24 : _GEN_7084; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8115 = ~quene ? ram_1_25 : _GEN_7085; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8116 = ~quene ? ram_1_26 : _GEN_7086; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8117 = ~quene ? ram_1_27 : _GEN_7087; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8118 = ~quene ? ram_1_28 : _GEN_7088; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8119 = ~quene ? ram_1_29 : _GEN_7089; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8120 = ~quene ? ram_1_30 : _GEN_7090; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8121 = ~quene ? ram_1_31 : _GEN_7091; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8122 = ~quene ? ram_1_32 : _GEN_7092; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8123 = ~quene ? ram_1_33 : _GEN_7093; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8124 = ~quene ? ram_1_34 : _GEN_7094; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8125 = ~quene ? ram_1_35 : _GEN_7095; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8126 = ~quene ? ram_1_36 : _GEN_7096; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8127 = ~quene ? ram_1_37 : _GEN_7097; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8128 = ~quene ? ram_1_38 : _GEN_7098; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8129 = ~quene ? ram_1_39 : _GEN_7099; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8130 = ~quene ? ram_1_40 : _GEN_7100; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8131 = ~quene ? ram_1_41 : _GEN_7101; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8132 = ~quene ? ram_1_42 : _GEN_7102; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8133 = ~quene ? ram_1_43 : _GEN_7103; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8134 = ~quene ? ram_1_44 : _GEN_7104; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8135 = ~quene ? ram_1_45 : _GEN_7105; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8136 = ~quene ? ram_1_46 : _GEN_7106; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8137 = ~quene ? ram_1_47 : _GEN_7107; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8138 = ~quene ? ram_1_48 : _GEN_7108; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8139 = ~quene ? ram_1_49 : _GEN_7109; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8140 = ~quene ? ram_1_50 : _GEN_7110; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8141 = ~quene ? ram_1_51 : _GEN_7111; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8142 = ~quene ? ram_1_52 : _GEN_7112; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8143 = ~quene ? ram_1_53 : _GEN_7113; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8144 = ~quene ? ram_1_54 : _GEN_7114; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8145 = ~quene ? ram_1_55 : _GEN_7115; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8146 = ~quene ? ram_1_56 : _GEN_7116; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8147 = ~quene ? ram_1_57 : _GEN_7117; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8148 = ~quene ? ram_1_58 : _GEN_7118; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8149 = ~quene ? ram_1_59 : _GEN_7119; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8150 = ~quene ? ram_1_60 : _GEN_7120; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8151 = ~quene ? ram_1_61 : _GEN_7121; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8152 = ~quene ? ram_1_62 : _GEN_7122; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8153 = ~quene ? ram_1_63 : _GEN_7123; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8154 = ~quene ? ram_1_64 : _GEN_7124; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8155 = ~quene ? ram_1_65 : _GEN_7125; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8156 = ~quene ? ram_1_66 : _GEN_7126; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8157 = ~quene ? ram_1_67 : _GEN_7127; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8158 = ~quene ? ram_1_68 : _GEN_7128; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8159 = ~quene ? ram_1_69 : _GEN_7129; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8160 = ~quene ? ram_1_70 : _GEN_7130; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8161 = ~quene ? ram_1_71 : _GEN_7131; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8162 = ~quene ? ram_1_72 : _GEN_7132; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8163 = ~quene ? ram_1_73 : _GEN_7133; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8164 = ~quene ? ram_1_74 : _GEN_7134; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8165 = ~quene ? ram_1_75 : _GEN_7135; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8166 = ~quene ? ram_1_76 : _GEN_7136; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8167 = ~quene ? ram_1_77 : _GEN_7137; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8168 = ~quene ? ram_1_78 : _GEN_7138; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8169 = ~quene ? ram_1_79 : _GEN_7139; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8170 = ~quene ? ram_1_80 : _GEN_7140; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8171 = ~quene ? ram_1_81 : _GEN_7141; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8172 = ~quene ? ram_1_82 : _GEN_7142; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8173 = ~quene ? ram_1_83 : _GEN_7143; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8174 = ~quene ? ram_1_84 : _GEN_7144; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8175 = ~quene ? ram_1_85 : _GEN_7145; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8176 = ~quene ? ram_1_86 : _GEN_7146; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8177 = ~quene ? ram_1_87 : _GEN_7147; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8178 = ~quene ? ram_1_88 : _GEN_7148; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8179 = ~quene ? ram_1_89 : _GEN_7149; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8180 = ~quene ? ram_1_90 : _GEN_7150; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8181 = ~quene ? ram_1_91 : _GEN_7151; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8182 = ~quene ? ram_1_92 : _GEN_7152; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8183 = ~quene ? ram_1_93 : _GEN_7153; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8184 = ~quene ? ram_1_94 : _GEN_7154; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8185 = ~quene ? ram_1_95 : _GEN_7155; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8186 = ~quene ? ram_1_96 : _GEN_7156; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8187 = ~quene ? ram_1_97 : _GEN_7157; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8188 = ~quene ? ram_1_98 : _GEN_7158; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8189 = ~quene ? ram_1_99 : _GEN_7159; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8190 = ~quene ? ram_1_100 : _GEN_7160; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8191 = ~quene ? ram_1_101 : _GEN_7161; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8192 = ~quene ? ram_1_102 : _GEN_7162; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8193 = ~quene ? ram_1_103 : _GEN_7163; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8194 = ~quene ? ram_1_104 : _GEN_7164; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8195 = ~quene ? ram_1_105 : _GEN_7165; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8196 = ~quene ? ram_1_106 : _GEN_7166; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8197 = ~quene ? ram_1_107 : _GEN_7167; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8198 = ~quene ? ram_1_108 : _GEN_7168; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8199 = ~quene ? ram_1_109 : _GEN_7169; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8200 = ~quene ? ram_1_110 : _GEN_7170; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8201 = ~quene ? ram_1_111 : _GEN_7171; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8202 = ~quene ? ram_1_112 : _GEN_7172; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8203 = ~quene ? ram_1_113 : _GEN_7173; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8204 = ~quene ? ram_1_114 : _GEN_7174; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8205 = ~quene ? ram_1_115 : _GEN_7175; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8206 = ~quene ? ram_1_116 : _GEN_7176; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8207 = ~quene ? ram_1_117 : _GEN_7177; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8208 = ~quene ? ram_1_118 : _GEN_7178; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8209 = ~quene ? ram_1_119 : _GEN_7179; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8210 = ~quene ? ram_1_120 : _GEN_7180; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8211 = ~quene ? ram_1_121 : _GEN_7181; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8212 = ~quene ? ram_1_122 : _GEN_7182; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8213 = ~quene ? ram_1_123 : _GEN_7183; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8214 = ~quene ? ram_1_124 : _GEN_7184; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8215 = ~quene ? ram_1_125 : _GEN_7185; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8216 = ~quene ? ram_1_126 : _GEN_7186; // @[d_cache.scala 152:34 19:24]
  wire [63:0] _GEN_8217 = ~quene ? ram_1_127 : _GEN_7187; // @[d_cache.scala 152:34 19:24]
  wire [31:0] _GEN_8218 = ~quene ? tag_1_0 : _GEN_7188; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8219 = ~quene ? tag_1_1 : _GEN_7189; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8220 = ~quene ? tag_1_2 : _GEN_7190; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8221 = ~quene ? tag_1_3 : _GEN_7191; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8222 = ~quene ? tag_1_4 : _GEN_7192; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8223 = ~quene ? tag_1_5 : _GEN_7193; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8224 = ~quene ? tag_1_6 : _GEN_7194; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8225 = ~quene ? tag_1_7 : _GEN_7195; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8226 = ~quene ? tag_1_8 : _GEN_7196; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8227 = ~quene ? tag_1_9 : _GEN_7197; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8228 = ~quene ? tag_1_10 : _GEN_7198; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8229 = ~quene ? tag_1_11 : _GEN_7199; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8230 = ~quene ? tag_1_12 : _GEN_7200; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8231 = ~quene ? tag_1_13 : _GEN_7201; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8232 = ~quene ? tag_1_14 : _GEN_7202; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8233 = ~quene ? tag_1_15 : _GEN_7203; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8234 = ~quene ? tag_1_16 : _GEN_7204; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8235 = ~quene ? tag_1_17 : _GEN_7205; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8236 = ~quene ? tag_1_18 : _GEN_7206; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8237 = ~quene ? tag_1_19 : _GEN_7207; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8238 = ~quene ? tag_1_20 : _GEN_7208; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8239 = ~quene ? tag_1_21 : _GEN_7209; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8240 = ~quene ? tag_1_22 : _GEN_7210; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8241 = ~quene ? tag_1_23 : _GEN_7211; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8242 = ~quene ? tag_1_24 : _GEN_7212; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8243 = ~quene ? tag_1_25 : _GEN_7213; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8244 = ~quene ? tag_1_26 : _GEN_7214; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8245 = ~quene ? tag_1_27 : _GEN_7215; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8246 = ~quene ? tag_1_28 : _GEN_7216; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8247 = ~quene ? tag_1_29 : _GEN_7217; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8248 = ~quene ? tag_1_30 : _GEN_7218; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8249 = ~quene ? tag_1_31 : _GEN_7219; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8250 = ~quene ? tag_1_32 : _GEN_7220; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8251 = ~quene ? tag_1_33 : _GEN_7221; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8252 = ~quene ? tag_1_34 : _GEN_7222; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8253 = ~quene ? tag_1_35 : _GEN_7223; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8254 = ~quene ? tag_1_36 : _GEN_7224; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8255 = ~quene ? tag_1_37 : _GEN_7225; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8256 = ~quene ? tag_1_38 : _GEN_7226; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8257 = ~quene ? tag_1_39 : _GEN_7227; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8258 = ~quene ? tag_1_40 : _GEN_7228; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8259 = ~quene ? tag_1_41 : _GEN_7229; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8260 = ~quene ? tag_1_42 : _GEN_7230; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8261 = ~quene ? tag_1_43 : _GEN_7231; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8262 = ~quene ? tag_1_44 : _GEN_7232; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8263 = ~quene ? tag_1_45 : _GEN_7233; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8264 = ~quene ? tag_1_46 : _GEN_7234; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8265 = ~quene ? tag_1_47 : _GEN_7235; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8266 = ~quene ? tag_1_48 : _GEN_7236; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8267 = ~quene ? tag_1_49 : _GEN_7237; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8268 = ~quene ? tag_1_50 : _GEN_7238; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8269 = ~quene ? tag_1_51 : _GEN_7239; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8270 = ~quene ? tag_1_52 : _GEN_7240; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8271 = ~quene ? tag_1_53 : _GEN_7241; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8272 = ~quene ? tag_1_54 : _GEN_7242; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8273 = ~quene ? tag_1_55 : _GEN_7243; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8274 = ~quene ? tag_1_56 : _GEN_7244; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8275 = ~quene ? tag_1_57 : _GEN_7245; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8276 = ~quene ? tag_1_58 : _GEN_7246; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8277 = ~quene ? tag_1_59 : _GEN_7247; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8278 = ~quene ? tag_1_60 : _GEN_7248; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8279 = ~quene ? tag_1_61 : _GEN_7249; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8280 = ~quene ? tag_1_62 : _GEN_7250; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8281 = ~quene ? tag_1_63 : _GEN_7251; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8282 = ~quene ? tag_1_64 : _GEN_7252; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8283 = ~quene ? tag_1_65 : _GEN_7253; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8284 = ~quene ? tag_1_66 : _GEN_7254; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8285 = ~quene ? tag_1_67 : _GEN_7255; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8286 = ~quene ? tag_1_68 : _GEN_7256; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8287 = ~quene ? tag_1_69 : _GEN_7257; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8288 = ~quene ? tag_1_70 : _GEN_7258; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8289 = ~quene ? tag_1_71 : _GEN_7259; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8290 = ~quene ? tag_1_72 : _GEN_7260; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8291 = ~quene ? tag_1_73 : _GEN_7261; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8292 = ~quene ? tag_1_74 : _GEN_7262; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8293 = ~quene ? tag_1_75 : _GEN_7263; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8294 = ~quene ? tag_1_76 : _GEN_7264; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8295 = ~quene ? tag_1_77 : _GEN_7265; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8296 = ~quene ? tag_1_78 : _GEN_7266; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8297 = ~quene ? tag_1_79 : _GEN_7267; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8298 = ~quene ? tag_1_80 : _GEN_7268; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8299 = ~quene ? tag_1_81 : _GEN_7269; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8300 = ~quene ? tag_1_82 : _GEN_7270; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8301 = ~quene ? tag_1_83 : _GEN_7271; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8302 = ~quene ? tag_1_84 : _GEN_7272; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8303 = ~quene ? tag_1_85 : _GEN_7273; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8304 = ~quene ? tag_1_86 : _GEN_7274; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8305 = ~quene ? tag_1_87 : _GEN_7275; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8306 = ~quene ? tag_1_88 : _GEN_7276; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8307 = ~quene ? tag_1_89 : _GEN_7277; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8308 = ~quene ? tag_1_90 : _GEN_7278; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8309 = ~quene ? tag_1_91 : _GEN_7279; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8310 = ~quene ? tag_1_92 : _GEN_7280; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8311 = ~quene ? tag_1_93 : _GEN_7281; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8312 = ~quene ? tag_1_94 : _GEN_7282; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8313 = ~quene ? tag_1_95 : _GEN_7283; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8314 = ~quene ? tag_1_96 : _GEN_7284; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8315 = ~quene ? tag_1_97 : _GEN_7285; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8316 = ~quene ? tag_1_98 : _GEN_7286; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8317 = ~quene ? tag_1_99 : _GEN_7287; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8318 = ~quene ? tag_1_100 : _GEN_7288; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8319 = ~quene ? tag_1_101 : _GEN_7289; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8320 = ~quene ? tag_1_102 : _GEN_7290; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8321 = ~quene ? tag_1_103 : _GEN_7291; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8322 = ~quene ? tag_1_104 : _GEN_7292; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8323 = ~quene ? tag_1_105 : _GEN_7293; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8324 = ~quene ? tag_1_106 : _GEN_7294; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8325 = ~quene ? tag_1_107 : _GEN_7295; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8326 = ~quene ? tag_1_108 : _GEN_7296; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8327 = ~quene ? tag_1_109 : _GEN_7297; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8328 = ~quene ? tag_1_110 : _GEN_7298; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8329 = ~quene ? tag_1_111 : _GEN_7299; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8330 = ~quene ? tag_1_112 : _GEN_7300; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8331 = ~quene ? tag_1_113 : _GEN_7301; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8332 = ~quene ? tag_1_114 : _GEN_7302; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8333 = ~quene ? tag_1_115 : _GEN_7303; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8334 = ~quene ? tag_1_116 : _GEN_7304; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8335 = ~quene ? tag_1_117 : _GEN_7305; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8336 = ~quene ? tag_1_118 : _GEN_7306; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8337 = ~quene ? tag_1_119 : _GEN_7307; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8338 = ~quene ? tag_1_120 : _GEN_7308; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8339 = ~quene ? tag_1_121 : _GEN_7309; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8340 = ~quene ? tag_1_122 : _GEN_7310; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8341 = ~quene ? tag_1_123 : _GEN_7311; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8342 = ~quene ? tag_1_124 : _GEN_7312; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8343 = ~quene ? tag_1_125 : _GEN_7313; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8344 = ~quene ? tag_1_126 : _GEN_7314; // @[d_cache.scala 152:34 23:24]
  wire [31:0] _GEN_8345 = ~quene ? tag_1_127 : _GEN_7315; // @[d_cache.scala 152:34 23:24]
  wire  _GEN_8346 = ~quene ? dirty_1_0 : _GEN_7316; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8347 = ~quene ? dirty_1_1 : _GEN_7317; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8348 = ~quene ? dirty_1_2 : _GEN_7318; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8349 = ~quene ? dirty_1_3 : _GEN_7319; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8350 = ~quene ? dirty_1_4 : _GEN_7320; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8351 = ~quene ? dirty_1_5 : _GEN_7321; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8352 = ~quene ? dirty_1_6 : _GEN_7322; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8353 = ~quene ? dirty_1_7 : _GEN_7323; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8354 = ~quene ? dirty_1_8 : _GEN_7324; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8355 = ~quene ? dirty_1_9 : _GEN_7325; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8356 = ~quene ? dirty_1_10 : _GEN_7326; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8357 = ~quene ? dirty_1_11 : _GEN_7327; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8358 = ~quene ? dirty_1_12 : _GEN_7328; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8359 = ~quene ? dirty_1_13 : _GEN_7329; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8360 = ~quene ? dirty_1_14 : _GEN_7330; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8361 = ~quene ? dirty_1_15 : _GEN_7331; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8362 = ~quene ? dirty_1_16 : _GEN_7332; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8363 = ~quene ? dirty_1_17 : _GEN_7333; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8364 = ~quene ? dirty_1_18 : _GEN_7334; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8365 = ~quene ? dirty_1_19 : _GEN_7335; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8366 = ~quene ? dirty_1_20 : _GEN_7336; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8367 = ~quene ? dirty_1_21 : _GEN_7337; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8368 = ~quene ? dirty_1_22 : _GEN_7338; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8369 = ~quene ? dirty_1_23 : _GEN_7339; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8370 = ~quene ? dirty_1_24 : _GEN_7340; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8371 = ~quene ? dirty_1_25 : _GEN_7341; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8372 = ~quene ? dirty_1_26 : _GEN_7342; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8373 = ~quene ? dirty_1_27 : _GEN_7343; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8374 = ~quene ? dirty_1_28 : _GEN_7344; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8375 = ~quene ? dirty_1_29 : _GEN_7345; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8376 = ~quene ? dirty_1_30 : _GEN_7346; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8377 = ~quene ? dirty_1_31 : _GEN_7347; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8378 = ~quene ? dirty_1_32 : _GEN_7348; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8379 = ~quene ? dirty_1_33 : _GEN_7349; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8380 = ~quene ? dirty_1_34 : _GEN_7350; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8381 = ~quene ? dirty_1_35 : _GEN_7351; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8382 = ~quene ? dirty_1_36 : _GEN_7352; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8383 = ~quene ? dirty_1_37 : _GEN_7353; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8384 = ~quene ? dirty_1_38 : _GEN_7354; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8385 = ~quene ? dirty_1_39 : _GEN_7355; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8386 = ~quene ? dirty_1_40 : _GEN_7356; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8387 = ~quene ? dirty_1_41 : _GEN_7357; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8388 = ~quene ? dirty_1_42 : _GEN_7358; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8389 = ~quene ? dirty_1_43 : _GEN_7359; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8390 = ~quene ? dirty_1_44 : _GEN_7360; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8391 = ~quene ? dirty_1_45 : _GEN_7361; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8392 = ~quene ? dirty_1_46 : _GEN_7362; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8393 = ~quene ? dirty_1_47 : _GEN_7363; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8394 = ~quene ? dirty_1_48 : _GEN_7364; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8395 = ~quene ? dirty_1_49 : _GEN_7365; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8396 = ~quene ? dirty_1_50 : _GEN_7366; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8397 = ~quene ? dirty_1_51 : _GEN_7367; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8398 = ~quene ? dirty_1_52 : _GEN_7368; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8399 = ~quene ? dirty_1_53 : _GEN_7369; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8400 = ~quene ? dirty_1_54 : _GEN_7370; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8401 = ~quene ? dirty_1_55 : _GEN_7371; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8402 = ~quene ? dirty_1_56 : _GEN_7372; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8403 = ~quene ? dirty_1_57 : _GEN_7373; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8404 = ~quene ? dirty_1_58 : _GEN_7374; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8405 = ~quene ? dirty_1_59 : _GEN_7375; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8406 = ~quene ? dirty_1_60 : _GEN_7376; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8407 = ~quene ? dirty_1_61 : _GEN_7377; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8408 = ~quene ? dirty_1_62 : _GEN_7378; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8409 = ~quene ? dirty_1_63 : _GEN_7379; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8410 = ~quene ? dirty_1_64 : _GEN_7380; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8411 = ~quene ? dirty_1_65 : _GEN_7381; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8412 = ~quene ? dirty_1_66 : _GEN_7382; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8413 = ~quene ? dirty_1_67 : _GEN_7383; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8414 = ~quene ? dirty_1_68 : _GEN_7384; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8415 = ~quene ? dirty_1_69 : _GEN_7385; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8416 = ~quene ? dirty_1_70 : _GEN_7386; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8417 = ~quene ? dirty_1_71 : _GEN_7387; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8418 = ~quene ? dirty_1_72 : _GEN_7388; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8419 = ~quene ? dirty_1_73 : _GEN_7389; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8420 = ~quene ? dirty_1_74 : _GEN_7390; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8421 = ~quene ? dirty_1_75 : _GEN_7391; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8422 = ~quene ? dirty_1_76 : _GEN_7392; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8423 = ~quene ? dirty_1_77 : _GEN_7393; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8424 = ~quene ? dirty_1_78 : _GEN_7394; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8425 = ~quene ? dirty_1_79 : _GEN_7395; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8426 = ~quene ? dirty_1_80 : _GEN_7396; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8427 = ~quene ? dirty_1_81 : _GEN_7397; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8428 = ~quene ? dirty_1_82 : _GEN_7398; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8429 = ~quene ? dirty_1_83 : _GEN_7399; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8430 = ~quene ? dirty_1_84 : _GEN_7400; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8431 = ~quene ? dirty_1_85 : _GEN_7401; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8432 = ~quene ? dirty_1_86 : _GEN_7402; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8433 = ~quene ? dirty_1_87 : _GEN_7403; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8434 = ~quene ? dirty_1_88 : _GEN_7404; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8435 = ~quene ? dirty_1_89 : _GEN_7405; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8436 = ~quene ? dirty_1_90 : _GEN_7406; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8437 = ~quene ? dirty_1_91 : _GEN_7407; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8438 = ~quene ? dirty_1_92 : _GEN_7408; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8439 = ~quene ? dirty_1_93 : _GEN_7409; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8440 = ~quene ? dirty_1_94 : _GEN_7410; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8441 = ~quene ? dirty_1_95 : _GEN_7411; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8442 = ~quene ? dirty_1_96 : _GEN_7412; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8443 = ~quene ? dirty_1_97 : _GEN_7413; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8444 = ~quene ? dirty_1_98 : _GEN_7414; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8445 = ~quene ? dirty_1_99 : _GEN_7415; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8446 = ~quene ? dirty_1_100 : _GEN_7416; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8447 = ~quene ? dirty_1_101 : _GEN_7417; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8448 = ~quene ? dirty_1_102 : _GEN_7418; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8449 = ~quene ? dirty_1_103 : _GEN_7419; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8450 = ~quene ? dirty_1_104 : _GEN_7420; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8451 = ~quene ? dirty_1_105 : _GEN_7421; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8452 = ~quene ? dirty_1_106 : _GEN_7422; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8453 = ~quene ? dirty_1_107 : _GEN_7423; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8454 = ~quene ? dirty_1_108 : _GEN_7424; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8455 = ~quene ? dirty_1_109 : _GEN_7425; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8456 = ~quene ? dirty_1_110 : _GEN_7426; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8457 = ~quene ? dirty_1_111 : _GEN_7427; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8458 = ~quene ? dirty_1_112 : _GEN_7428; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8459 = ~quene ? dirty_1_113 : _GEN_7429; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8460 = ~quene ? dirty_1_114 : _GEN_7430; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8461 = ~quene ? dirty_1_115 : _GEN_7431; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8462 = ~quene ? dirty_1_116 : _GEN_7432; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8463 = ~quene ? dirty_1_117 : _GEN_7433; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8464 = ~quene ? dirty_1_118 : _GEN_7434; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8465 = ~quene ? dirty_1_119 : _GEN_7435; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8466 = ~quene ? dirty_1_120 : _GEN_7436; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8467 = ~quene ? dirty_1_121 : _GEN_7437; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8468 = ~quene ? dirty_1_122 : _GEN_7438; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8469 = ~quene ? dirty_1_123 : _GEN_7439; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8470 = ~quene ? dirty_1_124 : _GEN_7440; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8471 = ~quene ? dirty_1_125 : _GEN_7441; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8472 = ~quene ? dirty_1_126 : _GEN_7442; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8473 = ~quene ? dirty_1_127 : _GEN_7443; // @[d_cache.scala 152:34 27:26]
  wire  _GEN_8474 = ~quene ? valid_1_0 : _GEN_7444; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8475 = ~quene ? valid_1_1 : _GEN_7445; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8476 = ~quene ? valid_1_2 : _GEN_7446; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8477 = ~quene ? valid_1_3 : _GEN_7447; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8478 = ~quene ? valid_1_4 : _GEN_7448; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8479 = ~quene ? valid_1_5 : _GEN_7449; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8480 = ~quene ? valid_1_6 : _GEN_7450; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8481 = ~quene ? valid_1_7 : _GEN_7451; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8482 = ~quene ? valid_1_8 : _GEN_7452; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8483 = ~quene ? valid_1_9 : _GEN_7453; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8484 = ~quene ? valid_1_10 : _GEN_7454; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8485 = ~quene ? valid_1_11 : _GEN_7455; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8486 = ~quene ? valid_1_12 : _GEN_7456; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8487 = ~quene ? valid_1_13 : _GEN_7457; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8488 = ~quene ? valid_1_14 : _GEN_7458; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8489 = ~quene ? valid_1_15 : _GEN_7459; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8490 = ~quene ? valid_1_16 : _GEN_7460; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8491 = ~quene ? valid_1_17 : _GEN_7461; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8492 = ~quene ? valid_1_18 : _GEN_7462; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8493 = ~quene ? valid_1_19 : _GEN_7463; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8494 = ~quene ? valid_1_20 : _GEN_7464; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8495 = ~quene ? valid_1_21 : _GEN_7465; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8496 = ~quene ? valid_1_22 : _GEN_7466; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8497 = ~quene ? valid_1_23 : _GEN_7467; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8498 = ~quene ? valid_1_24 : _GEN_7468; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8499 = ~quene ? valid_1_25 : _GEN_7469; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8500 = ~quene ? valid_1_26 : _GEN_7470; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8501 = ~quene ? valid_1_27 : _GEN_7471; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8502 = ~quene ? valid_1_28 : _GEN_7472; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8503 = ~quene ? valid_1_29 : _GEN_7473; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8504 = ~quene ? valid_1_30 : _GEN_7474; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8505 = ~quene ? valid_1_31 : _GEN_7475; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8506 = ~quene ? valid_1_32 : _GEN_7476; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8507 = ~quene ? valid_1_33 : _GEN_7477; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8508 = ~quene ? valid_1_34 : _GEN_7478; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8509 = ~quene ? valid_1_35 : _GEN_7479; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8510 = ~quene ? valid_1_36 : _GEN_7480; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8511 = ~quene ? valid_1_37 : _GEN_7481; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8512 = ~quene ? valid_1_38 : _GEN_7482; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8513 = ~quene ? valid_1_39 : _GEN_7483; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8514 = ~quene ? valid_1_40 : _GEN_7484; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8515 = ~quene ? valid_1_41 : _GEN_7485; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8516 = ~quene ? valid_1_42 : _GEN_7486; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8517 = ~quene ? valid_1_43 : _GEN_7487; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8518 = ~quene ? valid_1_44 : _GEN_7488; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8519 = ~quene ? valid_1_45 : _GEN_7489; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8520 = ~quene ? valid_1_46 : _GEN_7490; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8521 = ~quene ? valid_1_47 : _GEN_7491; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8522 = ~quene ? valid_1_48 : _GEN_7492; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8523 = ~quene ? valid_1_49 : _GEN_7493; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8524 = ~quene ? valid_1_50 : _GEN_7494; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8525 = ~quene ? valid_1_51 : _GEN_7495; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8526 = ~quene ? valid_1_52 : _GEN_7496; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8527 = ~quene ? valid_1_53 : _GEN_7497; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8528 = ~quene ? valid_1_54 : _GEN_7498; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8529 = ~quene ? valid_1_55 : _GEN_7499; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8530 = ~quene ? valid_1_56 : _GEN_7500; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8531 = ~quene ? valid_1_57 : _GEN_7501; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8532 = ~quene ? valid_1_58 : _GEN_7502; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8533 = ~quene ? valid_1_59 : _GEN_7503; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8534 = ~quene ? valid_1_60 : _GEN_7504; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8535 = ~quene ? valid_1_61 : _GEN_7505; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8536 = ~quene ? valid_1_62 : _GEN_7506; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8537 = ~quene ? valid_1_63 : _GEN_7507; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8538 = ~quene ? valid_1_64 : _GEN_7508; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8539 = ~quene ? valid_1_65 : _GEN_7509; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8540 = ~quene ? valid_1_66 : _GEN_7510; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8541 = ~quene ? valid_1_67 : _GEN_7511; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8542 = ~quene ? valid_1_68 : _GEN_7512; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8543 = ~quene ? valid_1_69 : _GEN_7513; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8544 = ~quene ? valid_1_70 : _GEN_7514; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8545 = ~quene ? valid_1_71 : _GEN_7515; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8546 = ~quene ? valid_1_72 : _GEN_7516; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8547 = ~quene ? valid_1_73 : _GEN_7517; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8548 = ~quene ? valid_1_74 : _GEN_7518; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8549 = ~quene ? valid_1_75 : _GEN_7519; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8550 = ~quene ? valid_1_76 : _GEN_7520; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8551 = ~quene ? valid_1_77 : _GEN_7521; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8552 = ~quene ? valid_1_78 : _GEN_7522; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8553 = ~quene ? valid_1_79 : _GEN_7523; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8554 = ~quene ? valid_1_80 : _GEN_7524; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8555 = ~quene ? valid_1_81 : _GEN_7525; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8556 = ~quene ? valid_1_82 : _GEN_7526; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8557 = ~quene ? valid_1_83 : _GEN_7527; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8558 = ~quene ? valid_1_84 : _GEN_7528; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8559 = ~quene ? valid_1_85 : _GEN_7529; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8560 = ~quene ? valid_1_86 : _GEN_7530; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8561 = ~quene ? valid_1_87 : _GEN_7531; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8562 = ~quene ? valid_1_88 : _GEN_7532; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8563 = ~quene ? valid_1_89 : _GEN_7533; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8564 = ~quene ? valid_1_90 : _GEN_7534; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8565 = ~quene ? valid_1_91 : _GEN_7535; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8566 = ~quene ? valid_1_92 : _GEN_7536; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8567 = ~quene ? valid_1_93 : _GEN_7537; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8568 = ~quene ? valid_1_94 : _GEN_7538; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8569 = ~quene ? valid_1_95 : _GEN_7539; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8570 = ~quene ? valid_1_96 : _GEN_7540; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8571 = ~quene ? valid_1_97 : _GEN_7541; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8572 = ~quene ? valid_1_98 : _GEN_7542; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8573 = ~quene ? valid_1_99 : _GEN_7543; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8574 = ~quene ? valid_1_100 : _GEN_7544; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8575 = ~quene ? valid_1_101 : _GEN_7545; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8576 = ~quene ? valid_1_102 : _GEN_7546; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8577 = ~quene ? valid_1_103 : _GEN_7547; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8578 = ~quene ? valid_1_104 : _GEN_7548; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8579 = ~quene ? valid_1_105 : _GEN_7549; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8580 = ~quene ? valid_1_106 : _GEN_7550; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8581 = ~quene ? valid_1_107 : _GEN_7551; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8582 = ~quene ? valid_1_108 : _GEN_7552; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8583 = ~quene ? valid_1_109 : _GEN_7553; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8584 = ~quene ? valid_1_110 : _GEN_7554; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8585 = ~quene ? valid_1_111 : _GEN_7555; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8586 = ~quene ? valid_1_112 : _GEN_7556; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8587 = ~quene ? valid_1_113 : _GEN_7557; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8588 = ~quene ? valid_1_114 : _GEN_7558; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8589 = ~quene ? valid_1_115 : _GEN_7559; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8590 = ~quene ? valid_1_116 : _GEN_7560; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8591 = ~quene ? valid_1_117 : _GEN_7561; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8592 = ~quene ? valid_1_118 : _GEN_7562; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8593 = ~quene ? valid_1_119 : _GEN_7563; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8594 = ~quene ? valid_1_120 : _GEN_7564; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8595 = ~quene ? valid_1_121 : _GEN_7565; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8596 = ~quene ? valid_1_122 : _GEN_7566; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8597 = ~quene ? valid_1_123 : _GEN_7567; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8598 = ~quene ? valid_1_124 : _GEN_7568; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8599 = ~quene ? valid_1_125 : _GEN_7569; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8600 = ~quene ? valid_1_126 : _GEN_7570; // @[d_cache.scala 152:34 25:26]
  wire  _GEN_8601 = ~quene ? valid_1_127 : _GEN_7571; // @[d_cache.scala 152:34 25:26]
  wire [2:0] _GEN_8602 = unuse_way == 2'h2 ? 3'h7 : _GEN_8088; // @[d_cache.scala 145:40 146:23]
  wire [63:0] _GEN_8603 = unuse_way == 2'h2 ? _GEN_3598 : _GEN_8090; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8604 = unuse_way == 2'h2 ? _GEN_3599 : _GEN_8091; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8605 = unuse_way == 2'h2 ? _GEN_3600 : _GEN_8092; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8606 = unuse_way == 2'h2 ? _GEN_3601 : _GEN_8093; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8607 = unuse_way == 2'h2 ? _GEN_3602 : _GEN_8094; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8608 = unuse_way == 2'h2 ? _GEN_3603 : _GEN_8095; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8609 = unuse_way == 2'h2 ? _GEN_3604 : _GEN_8096; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8610 = unuse_way == 2'h2 ? _GEN_3605 : _GEN_8097; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8611 = unuse_way == 2'h2 ? _GEN_3606 : _GEN_8098; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8612 = unuse_way == 2'h2 ? _GEN_3607 : _GEN_8099; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8613 = unuse_way == 2'h2 ? _GEN_3608 : _GEN_8100; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8614 = unuse_way == 2'h2 ? _GEN_3609 : _GEN_8101; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8615 = unuse_way == 2'h2 ? _GEN_3610 : _GEN_8102; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8616 = unuse_way == 2'h2 ? _GEN_3611 : _GEN_8103; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8617 = unuse_way == 2'h2 ? _GEN_3612 : _GEN_8104; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8618 = unuse_way == 2'h2 ? _GEN_3613 : _GEN_8105; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8619 = unuse_way == 2'h2 ? _GEN_3614 : _GEN_8106; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8620 = unuse_way == 2'h2 ? _GEN_3615 : _GEN_8107; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8621 = unuse_way == 2'h2 ? _GEN_3616 : _GEN_8108; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8622 = unuse_way == 2'h2 ? _GEN_3617 : _GEN_8109; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8623 = unuse_way == 2'h2 ? _GEN_3618 : _GEN_8110; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8624 = unuse_way == 2'h2 ? _GEN_3619 : _GEN_8111; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8625 = unuse_way == 2'h2 ? _GEN_3620 : _GEN_8112; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8626 = unuse_way == 2'h2 ? _GEN_3621 : _GEN_8113; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8627 = unuse_way == 2'h2 ? _GEN_3622 : _GEN_8114; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8628 = unuse_way == 2'h2 ? _GEN_3623 : _GEN_8115; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8629 = unuse_way == 2'h2 ? _GEN_3624 : _GEN_8116; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8630 = unuse_way == 2'h2 ? _GEN_3625 : _GEN_8117; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8631 = unuse_way == 2'h2 ? _GEN_3626 : _GEN_8118; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8632 = unuse_way == 2'h2 ? _GEN_3627 : _GEN_8119; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8633 = unuse_way == 2'h2 ? _GEN_3628 : _GEN_8120; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8634 = unuse_way == 2'h2 ? _GEN_3629 : _GEN_8121; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8635 = unuse_way == 2'h2 ? _GEN_3630 : _GEN_8122; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8636 = unuse_way == 2'h2 ? _GEN_3631 : _GEN_8123; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8637 = unuse_way == 2'h2 ? _GEN_3632 : _GEN_8124; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8638 = unuse_way == 2'h2 ? _GEN_3633 : _GEN_8125; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8639 = unuse_way == 2'h2 ? _GEN_3634 : _GEN_8126; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8640 = unuse_way == 2'h2 ? _GEN_3635 : _GEN_8127; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8641 = unuse_way == 2'h2 ? _GEN_3636 : _GEN_8128; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8642 = unuse_way == 2'h2 ? _GEN_3637 : _GEN_8129; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8643 = unuse_way == 2'h2 ? _GEN_3638 : _GEN_8130; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8644 = unuse_way == 2'h2 ? _GEN_3639 : _GEN_8131; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8645 = unuse_way == 2'h2 ? _GEN_3640 : _GEN_8132; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8646 = unuse_way == 2'h2 ? _GEN_3641 : _GEN_8133; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8647 = unuse_way == 2'h2 ? _GEN_3642 : _GEN_8134; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8648 = unuse_way == 2'h2 ? _GEN_3643 : _GEN_8135; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8649 = unuse_way == 2'h2 ? _GEN_3644 : _GEN_8136; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8650 = unuse_way == 2'h2 ? _GEN_3645 : _GEN_8137; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8651 = unuse_way == 2'h2 ? _GEN_3646 : _GEN_8138; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8652 = unuse_way == 2'h2 ? _GEN_3647 : _GEN_8139; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8653 = unuse_way == 2'h2 ? _GEN_3648 : _GEN_8140; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8654 = unuse_way == 2'h2 ? _GEN_3649 : _GEN_8141; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8655 = unuse_way == 2'h2 ? _GEN_3650 : _GEN_8142; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8656 = unuse_way == 2'h2 ? _GEN_3651 : _GEN_8143; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8657 = unuse_way == 2'h2 ? _GEN_3652 : _GEN_8144; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8658 = unuse_way == 2'h2 ? _GEN_3653 : _GEN_8145; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8659 = unuse_way == 2'h2 ? _GEN_3654 : _GEN_8146; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8660 = unuse_way == 2'h2 ? _GEN_3655 : _GEN_8147; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8661 = unuse_way == 2'h2 ? _GEN_3656 : _GEN_8148; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8662 = unuse_way == 2'h2 ? _GEN_3657 : _GEN_8149; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8663 = unuse_way == 2'h2 ? _GEN_3658 : _GEN_8150; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8664 = unuse_way == 2'h2 ? _GEN_3659 : _GEN_8151; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8665 = unuse_way == 2'h2 ? _GEN_3660 : _GEN_8152; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8666 = unuse_way == 2'h2 ? _GEN_3661 : _GEN_8153; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8667 = unuse_way == 2'h2 ? _GEN_3662 : _GEN_8154; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8668 = unuse_way == 2'h2 ? _GEN_3663 : _GEN_8155; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8669 = unuse_way == 2'h2 ? _GEN_3664 : _GEN_8156; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8670 = unuse_way == 2'h2 ? _GEN_3665 : _GEN_8157; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8671 = unuse_way == 2'h2 ? _GEN_3666 : _GEN_8158; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8672 = unuse_way == 2'h2 ? _GEN_3667 : _GEN_8159; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8673 = unuse_way == 2'h2 ? _GEN_3668 : _GEN_8160; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8674 = unuse_way == 2'h2 ? _GEN_3669 : _GEN_8161; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8675 = unuse_way == 2'h2 ? _GEN_3670 : _GEN_8162; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8676 = unuse_way == 2'h2 ? _GEN_3671 : _GEN_8163; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8677 = unuse_way == 2'h2 ? _GEN_3672 : _GEN_8164; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8678 = unuse_way == 2'h2 ? _GEN_3673 : _GEN_8165; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8679 = unuse_way == 2'h2 ? _GEN_3674 : _GEN_8166; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8680 = unuse_way == 2'h2 ? _GEN_3675 : _GEN_8167; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8681 = unuse_way == 2'h2 ? _GEN_3676 : _GEN_8168; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8682 = unuse_way == 2'h2 ? _GEN_3677 : _GEN_8169; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8683 = unuse_way == 2'h2 ? _GEN_3678 : _GEN_8170; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8684 = unuse_way == 2'h2 ? _GEN_3679 : _GEN_8171; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8685 = unuse_way == 2'h2 ? _GEN_3680 : _GEN_8172; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8686 = unuse_way == 2'h2 ? _GEN_3681 : _GEN_8173; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8687 = unuse_way == 2'h2 ? _GEN_3682 : _GEN_8174; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8688 = unuse_way == 2'h2 ? _GEN_3683 : _GEN_8175; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8689 = unuse_way == 2'h2 ? _GEN_3684 : _GEN_8176; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8690 = unuse_way == 2'h2 ? _GEN_3685 : _GEN_8177; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8691 = unuse_way == 2'h2 ? _GEN_3686 : _GEN_8178; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8692 = unuse_way == 2'h2 ? _GEN_3687 : _GEN_8179; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8693 = unuse_way == 2'h2 ? _GEN_3688 : _GEN_8180; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8694 = unuse_way == 2'h2 ? _GEN_3689 : _GEN_8181; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8695 = unuse_way == 2'h2 ? _GEN_3690 : _GEN_8182; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8696 = unuse_way == 2'h2 ? _GEN_3691 : _GEN_8183; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8697 = unuse_way == 2'h2 ? _GEN_3692 : _GEN_8184; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8698 = unuse_way == 2'h2 ? _GEN_3693 : _GEN_8185; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8699 = unuse_way == 2'h2 ? _GEN_3694 : _GEN_8186; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8700 = unuse_way == 2'h2 ? _GEN_3695 : _GEN_8187; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8701 = unuse_way == 2'h2 ? _GEN_3696 : _GEN_8188; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8702 = unuse_way == 2'h2 ? _GEN_3697 : _GEN_8189; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8703 = unuse_way == 2'h2 ? _GEN_3698 : _GEN_8190; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8704 = unuse_way == 2'h2 ? _GEN_3699 : _GEN_8191; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8705 = unuse_way == 2'h2 ? _GEN_3700 : _GEN_8192; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8706 = unuse_way == 2'h2 ? _GEN_3701 : _GEN_8193; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8707 = unuse_way == 2'h2 ? _GEN_3702 : _GEN_8194; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8708 = unuse_way == 2'h2 ? _GEN_3703 : _GEN_8195; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8709 = unuse_way == 2'h2 ? _GEN_3704 : _GEN_8196; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8710 = unuse_way == 2'h2 ? _GEN_3705 : _GEN_8197; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8711 = unuse_way == 2'h2 ? _GEN_3706 : _GEN_8198; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8712 = unuse_way == 2'h2 ? _GEN_3707 : _GEN_8199; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8713 = unuse_way == 2'h2 ? _GEN_3708 : _GEN_8200; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8714 = unuse_way == 2'h2 ? _GEN_3709 : _GEN_8201; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8715 = unuse_way == 2'h2 ? _GEN_3710 : _GEN_8202; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8716 = unuse_way == 2'h2 ? _GEN_3711 : _GEN_8203; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8717 = unuse_way == 2'h2 ? _GEN_3712 : _GEN_8204; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8718 = unuse_way == 2'h2 ? _GEN_3713 : _GEN_8205; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8719 = unuse_way == 2'h2 ? _GEN_3714 : _GEN_8206; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8720 = unuse_way == 2'h2 ? _GEN_3715 : _GEN_8207; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8721 = unuse_way == 2'h2 ? _GEN_3716 : _GEN_8208; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8722 = unuse_way == 2'h2 ? _GEN_3717 : _GEN_8209; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8723 = unuse_way == 2'h2 ? _GEN_3718 : _GEN_8210; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8724 = unuse_way == 2'h2 ? _GEN_3719 : _GEN_8211; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8725 = unuse_way == 2'h2 ? _GEN_3720 : _GEN_8212; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8726 = unuse_way == 2'h2 ? _GEN_3721 : _GEN_8213; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8727 = unuse_way == 2'h2 ? _GEN_3722 : _GEN_8214; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8728 = unuse_way == 2'h2 ? _GEN_3723 : _GEN_8215; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8729 = unuse_way == 2'h2 ? _GEN_3724 : _GEN_8216; // @[d_cache.scala 145:40]
  wire [63:0] _GEN_8730 = unuse_way == 2'h2 ? _GEN_3725 : _GEN_8217; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8731 = unuse_way == 2'h2 ? _GEN_3726 : _GEN_8218; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8732 = unuse_way == 2'h2 ? _GEN_3727 : _GEN_8219; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8733 = unuse_way == 2'h2 ? _GEN_3728 : _GEN_8220; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8734 = unuse_way == 2'h2 ? _GEN_3729 : _GEN_8221; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8735 = unuse_way == 2'h2 ? _GEN_3730 : _GEN_8222; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8736 = unuse_way == 2'h2 ? _GEN_3731 : _GEN_8223; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8737 = unuse_way == 2'h2 ? _GEN_3732 : _GEN_8224; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8738 = unuse_way == 2'h2 ? _GEN_3733 : _GEN_8225; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8739 = unuse_way == 2'h2 ? _GEN_3734 : _GEN_8226; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8740 = unuse_way == 2'h2 ? _GEN_3735 : _GEN_8227; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8741 = unuse_way == 2'h2 ? _GEN_3736 : _GEN_8228; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8742 = unuse_way == 2'h2 ? _GEN_3737 : _GEN_8229; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8743 = unuse_way == 2'h2 ? _GEN_3738 : _GEN_8230; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8744 = unuse_way == 2'h2 ? _GEN_3739 : _GEN_8231; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8745 = unuse_way == 2'h2 ? _GEN_3740 : _GEN_8232; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8746 = unuse_way == 2'h2 ? _GEN_3741 : _GEN_8233; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8747 = unuse_way == 2'h2 ? _GEN_3742 : _GEN_8234; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8748 = unuse_way == 2'h2 ? _GEN_3743 : _GEN_8235; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8749 = unuse_way == 2'h2 ? _GEN_3744 : _GEN_8236; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8750 = unuse_way == 2'h2 ? _GEN_3745 : _GEN_8237; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8751 = unuse_way == 2'h2 ? _GEN_3746 : _GEN_8238; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8752 = unuse_way == 2'h2 ? _GEN_3747 : _GEN_8239; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8753 = unuse_way == 2'h2 ? _GEN_3748 : _GEN_8240; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8754 = unuse_way == 2'h2 ? _GEN_3749 : _GEN_8241; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8755 = unuse_way == 2'h2 ? _GEN_3750 : _GEN_8242; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8756 = unuse_way == 2'h2 ? _GEN_3751 : _GEN_8243; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8757 = unuse_way == 2'h2 ? _GEN_3752 : _GEN_8244; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8758 = unuse_way == 2'h2 ? _GEN_3753 : _GEN_8245; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8759 = unuse_way == 2'h2 ? _GEN_3754 : _GEN_8246; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8760 = unuse_way == 2'h2 ? _GEN_3755 : _GEN_8247; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8761 = unuse_way == 2'h2 ? _GEN_3756 : _GEN_8248; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8762 = unuse_way == 2'h2 ? _GEN_3757 : _GEN_8249; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8763 = unuse_way == 2'h2 ? _GEN_3758 : _GEN_8250; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8764 = unuse_way == 2'h2 ? _GEN_3759 : _GEN_8251; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8765 = unuse_way == 2'h2 ? _GEN_3760 : _GEN_8252; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8766 = unuse_way == 2'h2 ? _GEN_3761 : _GEN_8253; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8767 = unuse_way == 2'h2 ? _GEN_3762 : _GEN_8254; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8768 = unuse_way == 2'h2 ? _GEN_3763 : _GEN_8255; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8769 = unuse_way == 2'h2 ? _GEN_3764 : _GEN_8256; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8770 = unuse_way == 2'h2 ? _GEN_3765 : _GEN_8257; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8771 = unuse_way == 2'h2 ? _GEN_3766 : _GEN_8258; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8772 = unuse_way == 2'h2 ? _GEN_3767 : _GEN_8259; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8773 = unuse_way == 2'h2 ? _GEN_3768 : _GEN_8260; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8774 = unuse_way == 2'h2 ? _GEN_3769 : _GEN_8261; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8775 = unuse_way == 2'h2 ? _GEN_3770 : _GEN_8262; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8776 = unuse_way == 2'h2 ? _GEN_3771 : _GEN_8263; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8777 = unuse_way == 2'h2 ? _GEN_3772 : _GEN_8264; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8778 = unuse_way == 2'h2 ? _GEN_3773 : _GEN_8265; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8779 = unuse_way == 2'h2 ? _GEN_3774 : _GEN_8266; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8780 = unuse_way == 2'h2 ? _GEN_3775 : _GEN_8267; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8781 = unuse_way == 2'h2 ? _GEN_3776 : _GEN_8268; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8782 = unuse_way == 2'h2 ? _GEN_3777 : _GEN_8269; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8783 = unuse_way == 2'h2 ? _GEN_3778 : _GEN_8270; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8784 = unuse_way == 2'h2 ? _GEN_3779 : _GEN_8271; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8785 = unuse_way == 2'h2 ? _GEN_3780 : _GEN_8272; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8786 = unuse_way == 2'h2 ? _GEN_3781 : _GEN_8273; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8787 = unuse_way == 2'h2 ? _GEN_3782 : _GEN_8274; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8788 = unuse_way == 2'h2 ? _GEN_3783 : _GEN_8275; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8789 = unuse_way == 2'h2 ? _GEN_3784 : _GEN_8276; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8790 = unuse_way == 2'h2 ? _GEN_3785 : _GEN_8277; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8791 = unuse_way == 2'h2 ? _GEN_3786 : _GEN_8278; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8792 = unuse_way == 2'h2 ? _GEN_3787 : _GEN_8279; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8793 = unuse_way == 2'h2 ? _GEN_3788 : _GEN_8280; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8794 = unuse_way == 2'h2 ? _GEN_3789 : _GEN_8281; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8795 = unuse_way == 2'h2 ? _GEN_3790 : _GEN_8282; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8796 = unuse_way == 2'h2 ? _GEN_3791 : _GEN_8283; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8797 = unuse_way == 2'h2 ? _GEN_3792 : _GEN_8284; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8798 = unuse_way == 2'h2 ? _GEN_3793 : _GEN_8285; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8799 = unuse_way == 2'h2 ? _GEN_3794 : _GEN_8286; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8800 = unuse_way == 2'h2 ? _GEN_3795 : _GEN_8287; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8801 = unuse_way == 2'h2 ? _GEN_3796 : _GEN_8288; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8802 = unuse_way == 2'h2 ? _GEN_3797 : _GEN_8289; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8803 = unuse_way == 2'h2 ? _GEN_3798 : _GEN_8290; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8804 = unuse_way == 2'h2 ? _GEN_3799 : _GEN_8291; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8805 = unuse_way == 2'h2 ? _GEN_3800 : _GEN_8292; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8806 = unuse_way == 2'h2 ? _GEN_3801 : _GEN_8293; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8807 = unuse_way == 2'h2 ? _GEN_3802 : _GEN_8294; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8808 = unuse_way == 2'h2 ? _GEN_3803 : _GEN_8295; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8809 = unuse_way == 2'h2 ? _GEN_3804 : _GEN_8296; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8810 = unuse_way == 2'h2 ? _GEN_3805 : _GEN_8297; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8811 = unuse_way == 2'h2 ? _GEN_3806 : _GEN_8298; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8812 = unuse_way == 2'h2 ? _GEN_3807 : _GEN_8299; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8813 = unuse_way == 2'h2 ? _GEN_3808 : _GEN_8300; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8814 = unuse_way == 2'h2 ? _GEN_3809 : _GEN_8301; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8815 = unuse_way == 2'h2 ? _GEN_3810 : _GEN_8302; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8816 = unuse_way == 2'h2 ? _GEN_3811 : _GEN_8303; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8817 = unuse_way == 2'h2 ? _GEN_3812 : _GEN_8304; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8818 = unuse_way == 2'h2 ? _GEN_3813 : _GEN_8305; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8819 = unuse_way == 2'h2 ? _GEN_3814 : _GEN_8306; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8820 = unuse_way == 2'h2 ? _GEN_3815 : _GEN_8307; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8821 = unuse_way == 2'h2 ? _GEN_3816 : _GEN_8308; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8822 = unuse_way == 2'h2 ? _GEN_3817 : _GEN_8309; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8823 = unuse_way == 2'h2 ? _GEN_3818 : _GEN_8310; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8824 = unuse_way == 2'h2 ? _GEN_3819 : _GEN_8311; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8825 = unuse_way == 2'h2 ? _GEN_3820 : _GEN_8312; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8826 = unuse_way == 2'h2 ? _GEN_3821 : _GEN_8313; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8827 = unuse_way == 2'h2 ? _GEN_3822 : _GEN_8314; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8828 = unuse_way == 2'h2 ? _GEN_3823 : _GEN_8315; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8829 = unuse_way == 2'h2 ? _GEN_3824 : _GEN_8316; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8830 = unuse_way == 2'h2 ? _GEN_3825 : _GEN_8317; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8831 = unuse_way == 2'h2 ? _GEN_3826 : _GEN_8318; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8832 = unuse_way == 2'h2 ? _GEN_3827 : _GEN_8319; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8833 = unuse_way == 2'h2 ? _GEN_3828 : _GEN_8320; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8834 = unuse_way == 2'h2 ? _GEN_3829 : _GEN_8321; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8835 = unuse_way == 2'h2 ? _GEN_3830 : _GEN_8322; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8836 = unuse_way == 2'h2 ? _GEN_3831 : _GEN_8323; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8837 = unuse_way == 2'h2 ? _GEN_3832 : _GEN_8324; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8838 = unuse_way == 2'h2 ? _GEN_3833 : _GEN_8325; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8839 = unuse_way == 2'h2 ? _GEN_3834 : _GEN_8326; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8840 = unuse_way == 2'h2 ? _GEN_3835 : _GEN_8327; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8841 = unuse_way == 2'h2 ? _GEN_3836 : _GEN_8328; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8842 = unuse_way == 2'h2 ? _GEN_3837 : _GEN_8329; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8843 = unuse_way == 2'h2 ? _GEN_3838 : _GEN_8330; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8844 = unuse_way == 2'h2 ? _GEN_3839 : _GEN_8331; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8845 = unuse_way == 2'h2 ? _GEN_3840 : _GEN_8332; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8846 = unuse_way == 2'h2 ? _GEN_3841 : _GEN_8333; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8847 = unuse_way == 2'h2 ? _GEN_3842 : _GEN_8334; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8848 = unuse_way == 2'h2 ? _GEN_3843 : _GEN_8335; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8849 = unuse_way == 2'h2 ? _GEN_3844 : _GEN_8336; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8850 = unuse_way == 2'h2 ? _GEN_3845 : _GEN_8337; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8851 = unuse_way == 2'h2 ? _GEN_3846 : _GEN_8338; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8852 = unuse_way == 2'h2 ? _GEN_3847 : _GEN_8339; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8853 = unuse_way == 2'h2 ? _GEN_3848 : _GEN_8340; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8854 = unuse_way == 2'h2 ? _GEN_3849 : _GEN_8341; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8855 = unuse_way == 2'h2 ? _GEN_3850 : _GEN_8342; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8856 = unuse_way == 2'h2 ? _GEN_3851 : _GEN_8343; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8857 = unuse_way == 2'h2 ? _GEN_3852 : _GEN_8344; // @[d_cache.scala 145:40]
  wire [31:0] _GEN_8858 = unuse_way == 2'h2 ? _GEN_3853 : _GEN_8345; // @[d_cache.scala 145:40]
  wire  _GEN_8859 = unuse_way == 2'h2 ? _GEN_3854 : _GEN_8474; // @[d_cache.scala 145:40]
  wire  _GEN_8860 = unuse_way == 2'h2 ? _GEN_3855 : _GEN_8475; // @[d_cache.scala 145:40]
  wire  _GEN_8861 = unuse_way == 2'h2 ? _GEN_3856 : _GEN_8476; // @[d_cache.scala 145:40]
  wire  _GEN_8862 = unuse_way == 2'h2 ? _GEN_3857 : _GEN_8477; // @[d_cache.scala 145:40]
  wire  _GEN_8863 = unuse_way == 2'h2 ? _GEN_3858 : _GEN_8478; // @[d_cache.scala 145:40]
  wire  _GEN_8864 = unuse_way == 2'h2 ? _GEN_3859 : _GEN_8479; // @[d_cache.scala 145:40]
  wire  _GEN_8865 = unuse_way == 2'h2 ? _GEN_3860 : _GEN_8480; // @[d_cache.scala 145:40]
  wire  _GEN_8866 = unuse_way == 2'h2 ? _GEN_3861 : _GEN_8481; // @[d_cache.scala 145:40]
  wire  _GEN_8867 = unuse_way == 2'h2 ? _GEN_3862 : _GEN_8482; // @[d_cache.scala 145:40]
  wire  _GEN_8868 = unuse_way == 2'h2 ? _GEN_3863 : _GEN_8483; // @[d_cache.scala 145:40]
  wire  _GEN_8869 = unuse_way == 2'h2 ? _GEN_3864 : _GEN_8484; // @[d_cache.scala 145:40]
  wire  _GEN_8870 = unuse_way == 2'h2 ? _GEN_3865 : _GEN_8485; // @[d_cache.scala 145:40]
  wire  _GEN_8871 = unuse_way == 2'h2 ? _GEN_3866 : _GEN_8486; // @[d_cache.scala 145:40]
  wire  _GEN_8872 = unuse_way == 2'h2 ? _GEN_3867 : _GEN_8487; // @[d_cache.scala 145:40]
  wire  _GEN_8873 = unuse_way == 2'h2 ? _GEN_3868 : _GEN_8488; // @[d_cache.scala 145:40]
  wire  _GEN_8874 = unuse_way == 2'h2 ? _GEN_3869 : _GEN_8489; // @[d_cache.scala 145:40]
  wire  _GEN_8875 = unuse_way == 2'h2 ? _GEN_3870 : _GEN_8490; // @[d_cache.scala 145:40]
  wire  _GEN_8876 = unuse_way == 2'h2 ? _GEN_3871 : _GEN_8491; // @[d_cache.scala 145:40]
  wire  _GEN_8877 = unuse_way == 2'h2 ? _GEN_3872 : _GEN_8492; // @[d_cache.scala 145:40]
  wire  _GEN_8878 = unuse_way == 2'h2 ? _GEN_3873 : _GEN_8493; // @[d_cache.scala 145:40]
  wire  _GEN_8879 = unuse_way == 2'h2 ? _GEN_3874 : _GEN_8494; // @[d_cache.scala 145:40]
  wire  _GEN_8880 = unuse_way == 2'h2 ? _GEN_3875 : _GEN_8495; // @[d_cache.scala 145:40]
  wire  _GEN_8881 = unuse_way == 2'h2 ? _GEN_3876 : _GEN_8496; // @[d_cache.scala 145:40]
  wire  _GEN_8882 = unuse_way == 2'h2 ? _GEN_3877 : _GEN_8497; // @[d_cache.scala 145:40]
  wire  _GEN_8883 = unuse_way == 2'h2 ? _GEN_3878 : _GEN_8498; // @[d_cache.scala 145:40]
  wire  _GEN_8884 = unuse_way == 2'h2 ? _GEN_3879 : _GEN_8499; // @[d_cache.scala 145:40]
  wire  _GEN_8885 = unuse_way == 2'h2 ? _GEN_3880 : _GEN_8500; // @[d_cache.scala 145:40]
  wire  _GEN_8886 = unuse_way == 2'h2 ? _GEN_3881 : _GEN_8501; // @[d_cache.scala 145:40]
  wire  _GEN_8887 = unuse_way == 2'h2 ? _GEN_3882 : _GEN_8502; // @[d_cache.scala 145:40]
  wire  _GEN_8888 = unuse_way == 2'h2 ? _GEN_3883 : _GEN_8503; // @[d_cache.scala 145:40]
  wire  _GEN_8889 = unuse_way == 2'h2 ? _GEN_3884 : _GEN_8504; // @[d_cache.scala 145:40]
  wire  _GEN_8890 = unuse_way == 2'h2 ? _GEN_3885 : _GEN_8505; // @[d_cache.scala 145:40]
  wire  _GEN_8891 = unuse_way == 2'h2 ? _GEN_3886 : _GEN_8506; // @[d_cache.scala 145:40]
  wire  _GEN_8892 = unuse_way == 2'h2 ? _GEN_3887 : _GEN_8507; // @[d_cache.scala 145:40]
  wire  _GEN_8893 = unuse_way == 2'h2 ? _GEN_3888 : _GEN_8508; // @[d_cache.scala 145:40]
  wire  _GEN_8894 = unuse_way == 2'h2 ? _GEN_3889 : _GEN_8509; // @[d_cache.scala 145:40]
  wire  _GEN_8895 = unuse_way == 2'h2 ? _GEN_3890 : _GEN_8510; // @[d_cache.scala 145:40]
  wire  _GEN_8896 = unuse_way == 2'h2 ? _GEN_3891 : _GEN_8511; // @[d_cache.scala 145:40]
  wire  _GEN_8897 = unuse_way == 2'h2 ? _GEN_3892 : _GEN_8512; // @[d_cache.scala 145:40]
  wire  _GEN_8898 = unuse_way == 2'h2 ? _GEN_3893 : _GEN_8513; // @[d_cache.scala 145:40]
  wire  _GEN_8899 = unuse_way == 2'h2 ? _GEN_3894 : _GEN_8514; // @[d_cache.scala 145:40]
  wire  _GEN_8900 = unuse_way == 2'h2 ? _GEN_3895 : _GEN_8515; // @[d_cache.scala 145:40]
  wire  _GEN_8901 = unuse_way == 2'h2 ? _GEN_3896 : _GEN_8516; // @[d_cache.scala 145:40]
  wire  _GEN_8902 = unuse_way == 2'h2 ? _GEN_3897 : _GEN_8517; // @[d_cache.scala 145:40]
  wire  _GEN_8903 = unuse_way == 2'h2 ? _GEN_3898 : _GEN_8518; // @[d_cache.scala 145:40]
  wire  _GEN_8904 = unuse_way == 2'h2 ? _GEN_3899 : _GEN_8519; // @[d_cache.scala 145:40]
  wire  _GEN_8905 = unuse_way == 2'h2 ? _GEN_3900 : _GEN_8520; // @[d_cache.scala 145:40]
  wire  _GEN_8906 = unuse_way == 2'h2 ? _GEN_3901 : _GEN_8521; // @[d_cache.scala 145:40]
  wire  _GEN_8907 = unuse_way == 2'h2 ? _GEN_3902 : _GEN_8522; // @[d_cache.scala 145:40]
  wire  _GEN_8908 = unuse_way == 2'h2 ? _GEN_3903 : _GEN_8523; // @[d_cache.scala 145:40]
  wire  _GEN_8909 = unuse_way == 2'h2 ? _GEN_3904 : _GEN_8524; // @[d_cache.scala 145:40]
  wire  _GEN_8910 = unuse_way == 2'h2 ? _GEN_3905 : _GEN_8525; // @[d_cache.scala 145:40]
  wire  _GEN_8911 = unuse_way == 2'h2 ? _GEN_3906 : _GEN_8526; // @[d_cache.scala 145:40]
  wire  _GEN_8912 = unuse_way == 2'h2 ? _GEN_3907 : _GEN_8527; // @[d_cache.scala 145:40]
  wire  _GEN_8913 = unuse_way == 2'h2 ? _GEN_3908 : _GEN_8528; // @[d_cache.scala 145:40]
  wire  _GEN_8914 = unuse_way == 2'h2 ? _GEN_3909 : _GEN_8529; // @[d_cache.scala 145:40]
  wire  _GEN_8915 = unuse_way == 2'h2 ? _GEN_3910 : _GEN_8530; // @[d_cache.scala 145:40]
  wire  _GEN_8916 = unuse_way == 2'h2 ? _GEN_3911 : _GEN_8531; // @[d_cache.scala 145:40]
  wire  _GEN_8917 = unuse_way == 2'h2 ? _GEN_3912 : _GEN_8532; // @[d_cache.scala 145:40]
  wire  _GEN_8918 = unuse_way == 2'h2 ? _GEN_3913 : _GEN_8533; // @[d_cache.scala 145:40]
  wire  _GEN_8919 = unuse_way == 2'h2 ? _GEN_3914 : _GEN_8534; // @[d_cache.scala 145:40]
  wire  _GEN_8920 = unuse_way == 2'h2 ? _GEN_3915 : _GEN_8535; // @[d_cache.scala 145:40]
  wire  _GEN_8921 = unuse_way == 2'h2 ? _GEN_3916 : _GEN_8536; // @[d_cache.scala 145:40]
  wire  _GEN_8922 = unuse_way == 2'h2 ? _GEN_3917 : _GEN_8537; // @[d_cache.scala 145:40]
  wire  _GEN_8923 = unuse_way == 2'h2 ? _GEN_3918 : _GEN_8538; // @[d_cache.scala 145:40]
  wire  _GEN_8924 = unuse_way == 2'h2 ? _GEN_3919 : _GEN_8539; // @[d_cache.scala 145:40]
  wire  _GEN_8925 = unuse_way == 2'h2 ? _GEN_3920 : _GEN_8540; // @[d_cache.scala 145:40]
  wire  _GEN_8926 = unuse_way == 2'h2 ? _GEN_3921 : _GEN_8541; // @[d_cache.scala 145:40]
  wire  _GEN_8927 = unuse_way == 2'h2 ? _GEN_3922 : _GEN_8542; // @[d_cache.scala 145:40]
  wire  _GEN_8928 = unuse_way == 2'h2 ? _GEN_3923 : _GEN_8543; // @[d_cache.scala 145:40]
  wire  _GEN_8929 = unuse_way == 2'h2 ? _GEN_3924 : _GEN_8544; // @[d_cache.scala 145:40]
  wire  _GEN_8930 = unuse_way == 2'h2 ? _GEN_3925 : _GEN_8545; // @[d_cache.scala 145:40]
  wire  _GEN_8931 = unuse_way == 2'h2 ? _GEN_3926 : _GEN_8546; // @[d_cache.scala 145:40]
  wire  _GEN_8932 = unuse_way == 2'h2 ? _GEN_3927 : _GEN_8547; // @[d_cache.scala 145:40]
  wire  _GEN_8933 = unuse_way == 2'h2 ? _GEN_3928 : _GEN_8548; // @[d_cache.scala 145:40]
  wire  _GEN_8934 = unuse_way == 2'h2 ? _GEN_3929 : _GEN_8549; // @[d_cache.scala 145:40]
  wire  _GEN_8935 = unuse_way == 2'h2 ? _GEN_3930 : _GEN_8550; // @[d_cache.scala 145:40]
  wire  _GEN_8936 = unuse_way == 2'h2 ? _GEN_3931 : _GEN_8551; // @[d_cache.scala 145:40]
  wire  _GEN_8937 = unuse_way == 2'h2 ? _GEN_3932 : _GEN_8552; // @[d_cache.scala 145:40]
  wire  _GEN_8938 = unuse_way == 2'h2 ? _GEN_3933 : _GEN_8553; // @[d_cache.scala 145:40]
  wire  _GEN_8939 = unuse_way == 2'h2 ? _GEN_3934 : _GEN_8554; // @[d_cache.scala 145:40]
  wire  _GEN_8940 = unuse_way == 2'h2 ? _GEN_3935 : _GEN_8555; // @[d_cache.scala 145:40]
  wire  _GEN_8941 = unuse_way == 2'h2 ? _GEN_3936 : _GEN_8556; // @[d_cache.scala 145:40]
  wire  _GEN_8942 = unuse_way == 2'h2 ? _GEN_3937 : _GEN_8557; // @[d_cache.scala 145:40]
  wire  _GEN_8943 = unuse_way == 2'h2 ? _GEN_3938 : _GEN_8558; // @[d_cache.scala 145:40]
  wire  _GEN_8944 = unuse_way == 2'h2 ? _GEN_3939 : _GEN_8559; // @[d_cache.scala 145:40]
  wire  _GEN_8945 = unuse_way == 2'h2 ? _GEN_3940 : _GEN_8560; // @[d_cache.scala 145:40]
  wire  _GEN_8946 = unuse_way == 2'h2 ? _GEN_3941 : _GEN_8561; // @[d_cache.scala 145:40]
  wire  _GEN_8947 = unuse_way == 2'h2 ? _GEN_3942 : _GEN_8562; // @[d_cache.scala 145:40]
  wire  _GEN_8948 = unuse_way == 2'h2 ? _GEN_3943 : _GEN_8563; // @[d_cache.scala 145:40]
  wire  _GEN_8949 = unuse_way == 2'h2 ? _GEN_3944 : _GEN_8564; // @[d_cache.scala 145:40]
  wire  _GEN_8950 = unuse_way == 2'h2 ? _GEN_3945 : _GEN_8565; // @[d_cache.scala 145:40]
  wire  _GEN_8951 = unuse_way == 2'h2 ? _GEN_3946 : _GEN_8566; // @[d_cache.scala 145:40]
  wire  _GEN_8952 = unuse_way == 2'h2 ? _GEN_3947 : _GEN_8567; // @[d_cache.scala 145:40]
  wire  _GEN_8953 = unuse_way == 2'h2 ? _GEN_3948 : _GEN_8568; // @[d_cache.scala 145:40]
  wire  _GEN_8954 = unuse_way == 2'h2 ? _GEN_3949 : _GEN_8569; // @[d_cache.scala 145:40]
  wire  _GEN_8955 = unuse_way == 2'h2 ? _GEN_3950 : _GEN_8570; // @[d_cache.scala 145:40]
  wire  _GEN_8956 = unuse_way == 2'h2 ? _GEN_3951 : _GEN_8571; // @[d_cache.scala 145:40]
  wire  _GEN_8957 = unuse_way == 2'h2 ? _GEN_3952 : _GEN_8572; // @[d_cache.scala 145:40]
  wire  _GEN_8958 = unuse_way == 2'h2 ? _GEN_3953 : _GEN_8573; // @[d_cache.scala 145:40]
  wire  _GEN_8959 = unuse_way == 2'h2 ? _GEN_3954 : _GEN_8574; // @[d_cache.scala 145:40]
  wire  _GEN_8960 = unuse_way == 2'h2 ? _GEN_3955 : _GEN_8575; // @[d_cache.scala 145:40]
  wire  _GEN_8961 = unuse_way == 2'h2 ? _GEN_3956 : _GEN_8576; // @[d_cache.scala 145:40]
  wire  _GEN_8962 = unuse_way == 2'h2 ? _GEN_3957 : _GEN_8577; // @[d_cache.scala 145:40]
  wire  _GEN_8963 = unuse_way == 2'h2 ? _GEN_3958 : _GEN_8578; // @[d_cache.scala 145:40]
  wire  _GEN_8964 = unuse_way == 2'h2 ? _GEN_3959 : _GEN_8579; // @[d_cache.scala 145:40]
  wire  _GEN_8965 = unuse_way == 2'h2 ? _GEN_3960 : _GEN_8580; // @[d_cache.scala 145:40]
  wire  _GEN_8966 = unuse_way == 2'h2 ? _GEN_3961 : _GEN_8581; // @[d_cache.scala 145:40]
  wire  _GEN_8967 = unuse_way == 2'h2 ? _GEN_3962 : _GEN_8582; // @[d_cache.scala 145:40]
  wire  _GEN_8968 = unuse_way == 2'h2 ? _GEN_3963 : _GEN_8583; // @[d_cache.scala 145:40]
  wire  _GEN_8969 = unuse_way == 2'h2 ? _GEN_3964 : _GEN_8584; // @[d_cache.scala 145:40]
  wire  _GEN_8970 = unuse_way == 2'h2 ? _GEN_3965 : _GEN_8585; // @[d_cache.scala 145:40]
  wire  _GEN_8971 = unuse_way == 2'h2 ? _GEN_3966 : _GEN_8586; // @[d_cache.scala 145:40]
  wire  _GEN_8972 = unuse_way == 2'h2 ? _GEN_3967 : _GEN_8587; // @[d_cache.scala 145:40]
  wire  _GEN_8973 = unuse_way == 2'h2 ? _GEN_3968 : _GEN_8588; // @[d_cache.scala 145:40]
  wire  _GEN_8974 = unuse_way == 2'h2 ? _GEN_3969 : _GEN_8589; // @[d_cache.scala 145:40]
  wire  _GEN_8975 = unuse_way == 2'h2 ? _GEN_3970 : _GEN_8590; // @[d_cache.scala 145:40]
  wire  _GEN_8976 = unuse_way == 2'h2 ? _GEN_3971 : _GEN_8591; // @[d_cache.scala 145:40]
  wire  _GEN_8977 = unuse_way == 2'h2 ? _GEN_3972 : _GEN_8592; // @[d_cache.scala 145:40]
  wire  _GEN_8978 = unuse_way == 2'h2 ? _GEN_3973 : _GEN_8593; // @[d_cache.scala 145:40]
  wire  _GEN_8979 = unuse_way == 2'h2 ? _GEN_3974 : _GEN_8594; // @[d_cache.scala 145:40]
  wire  _GEN_8980 = unuse_way == 2'h2 ? _GEN_3975 : _GEN_8595; // @[d_cache.scala 145:40]
  wire  _GEN_8981 = unuse_way == 2'h2 ? _GEN_3976 : _GEN_8596; // @[d_cache.scala 145:40]
  wire  _GEN_8982 = unuse_way == 2'h2 ? _GEN_3977 : _GEN_8597; // @[d_cache.scala 145:40]
  wire  _GEN_8983 = unuse_way == 2'h2 ? _GEN_3978 : _GEN_8598; // @[d_cache.scala 145:40]
  wire  _GEN_8984 = unuse_way == 2'h2 ? _GEN_3979 : _GEN_8599; // @[d_cache.scala 145:40]
  wire  _GEN_8985 = unuse_way == 2'h2 ? _GEN_3980 : _GEN_8600; // @[d_cache.scala 145:40]
  wire  _GEN_8986 = unuse_way == 2'h2 ? _GEN_3981 : _GEN_8601; // @[d_cache.scala 145:40]
  wire  _GEN_8987 = unuse_way == 2'h2 ? 1'h0 : _T_46; // @[d_cache.scala 145:40 150:23]
  wire [63:0] _GEN_8988 = unuse_way == 2'h2 ? write_back_data : _GEN_7574; // @[d_cache.scala 145:40 31:34]
  wire [41:0] _GEN_8989 = unuse_way == 2'h2 ? {{10'd0}, write_back_addr} : _GEN_7575; // @[d_cache.scala 145:40 32:34]
  wire [63:0] _GEN_8990 = unuse_way == 2'h2 ? ram_0_0 : _GEN_7576; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_8991 = unuse_way == 2'h2 ? ram_0_1 : _GEN_7577; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_8992 = unuse_way == 2'h2 ? ram_0_2 : _GEN_7578; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_8993 = unuse_way == 2'h2 ? ram_0_3 : _GEN_7579; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_8994 = unuse_way == 2'h2 ? ram_0_4 : _GEN_7580; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_8995 = unuse_way == 2'h2 ? ram_0_5 : _GEN_7581; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_8996 = unuse_way == 2'h2 ? ram_0_6 : _GEN_7582; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_8997 = unuse_way == 2'h2 ? ram_0_7 : _GEN_7583; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_8998 = unuse_way == 2'h2 ? ram_0_8 : _GEN_7584; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_8999 = unuse_way == 2'h2 ? ram_0_9 : _GEN_7585; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9000 = unuse_way == 2'h2 ? ram_0_10 : _GEN_7586; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9001 = unuse_way == 2'h2 ? ram_0_11 : _GEN_7587; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9002 = unuse_way == 2'h2 ? ram_0_12 : _GEN_7588; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9003 = unuse_way == 2'h2 ? ram_0_13 : _GEN_7589; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9004 = unuse_way == 2'h2 ? ram_0_14 : _GEN_7590; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9005 = unuse_way == 2'h2 ? ram_0_15 : _GEN_7591; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9006 = unuse_way == 2'h2 ? ram_0_16 : _GEN_7592; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9007 = unuse_way == 2'h2 ? ram_0_17 : _GEN_7593; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9008 = unuse_way == 2'h2 ? ram_0_18 : _GEN_7594; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9009 = unuse_way == 2'h2 ? ram_0_19 : _GEN_7595; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9010 = unuse_way == 2'h2 ? ram_0_20 : _GEN_7596; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9011 = unuse_way == 2'h2 ? ram_0_21 : _GEN_7597; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9012 = unuse_way == 2'h2 ? ram_0_22 : _GEN_7598; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9013 = unuse_way == 2'h2 ? ram_0_23 : _GEN_7599; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9014 = unuse_way == 2'h2 ? ram_0_24 : _GEN_7600; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9015 = unuse_way == 2'h2 ? ram_0_25 : _GEN_7601; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9016 = unuse_way == 2'h2 ? ram_0_26 : _GEN_7602; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9017 = unuse_way == 2'h2 ? ram_0_27 : _GEN_7603; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9018 = unuse_way == 2'h2 ? ram_0_28 : _GEN_7604; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9019 = unuse_way == 2'h2 ? ram_0_29 : _GEN_7605; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9020 = unuse_way == 2'h2 ? ram_0_30 : _GEN_7606; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9021 = unuse_way == 2'h2 ? ram_0_31 : _GEN_7607; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9022 = unuse_way == 2'h2 ? ram_0_32 : _GEN_7608; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9023 = unuse_way == 2'h2 ? ram_0_33 : _GEN_7609; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9024 = unuse_way == 2'h2 ? ram_0_34 : _GEN_7610; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9025 = unuse_way == 2'h2 ? ram_0_35 : _GEN_7611; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9026 = unuse_way == 2'h2 ? ram_0_36 : _GEN_7612; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9027 = unuse_way == 2'h2 ? ram_0_37 : _GEN_7613; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9028 = unuse_way == 2'h2 ? ram_0_38 : _GEN_7614; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9029 = unuse_way == 2'h2 ? ram_0_39 : _GEN_7615; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9030 = unuse_way == 2'h2 ? ram_0_40 : _GEN_7616; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9031 = unuse_way == 2'h2 ? ram_0_41 : _GEN_7617; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9032 = unuse_way == 2'h2 ? ram_0_42 : _GEN_7618; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9033 = unuse_way == 2'h2 ? ram_0_43 : _GEN_7619; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9034 = unuse_way == 2'h2 ? ram_0_44 : _GEN_7620; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9035 = unuse_way == 2'h2 ? ram_0_45 : _GEN_7621; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9036 = unuse_way == 2'h2 ? ram_0_46 : _GEN_7622; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9037 = unuse_way == 2'h2 ? ram_0_47 : _GEN_7623; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9038 = unuse_way == 2'h2 ? ram_0_48 : _GEN_7624; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9039 = unuse_way == 2'h2 ? ram_0_49 : _GEN_7625; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9040 = unuse_way == 2'h2 ? ram_0_50 : _GEN_7626; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9041 = unuse_way == 2'h2 ? ram_0_51 : _GEN_7627; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9042 = unuse_way == 2'h2 ? ram_0_52 : _GEN_7628; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9043 = unuse_way == 2'h2 ? ram_0_53 : _GEN_7629; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9044 = unuse_way == 2'h2 ? ram_0_54 : _GEN_7630; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9045 = unuse_way == 2'h2 ? ram_0_55 : _GEN_7631; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9046 = unuse_way == 2'h2 ? ram_0_56 : _GEN_7632; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9047 = unuse_way == 2'h2 ? ram_0_57 : _GEN_7633; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9048 = unuse_way == 2'h2 ? ram_0_58 : _GEN_7634; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9049 = unuse_way == 2'h2 ? ram_0_59 : _GEN_7635; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9050 = unuse_way == 2'h2 ? ram_0_60 : _GEN_7636; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9051 = unuse_way == 2'h2 ? ram_0_61 : _GEN_7637; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9052 = unuse_way == 2'h2 ? ram_0_62 : _GEN_7638; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9053 = unuse_way == 2'h2 ? ram_0_63 : _GEN_7639; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9054 = unuse_way == 2'h2 ? ram_0_64 : _GEN_7640; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9055 = unuse_way == 2'h2 ? ram_0_65 : _GEN_7641; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9056 = unuse_way == 2'h2 ? ram_0_66 : _GEN_7642; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9057 = unuse_way == 2'h2 ? ram_0_67 : _GEN_7643; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9058 = unuse_way == 2'h2 ? ram_0_68 : _GEN_7644; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9059 = unuse_way == 2'h2 ? ram_0_69 : _GEN_7645; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9060 = unuse_way == 2'h2 ? ram_0_70 : _GEN_7646; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9061 = unuse_way == 2'h2 ? ram_0_71 : _GEN_7647; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9062 = unuse_way == 2'h2 ? ram_0_72 : _GEN_7648; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9063 = unuse_way == 2'h2 ? ram_0_73 : _GEN_7649; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9064 = unuse_way == 2'h2 ? ram_0_74 : _GEN_7650; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9065 = unuse_way == 2'h2 ? ram_0_75 : _GEN_7651; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9066 = unuse_way == 2'h2 ? ram_0_76 : _GEN_7652; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9067 = unuse_way == 2'h2 ? ram_0_77 : _GEN_7653; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9068 = unuse_way == 2'h2 ? ram_0_78 : _GEN_7654; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9069 = unuse_way == 2'h2 ? ram_0_79 : _GEN_7655; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9070 = unuse_way == 2'h2 ? ram_0_80 : _GEN_7656; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9071 = unuse_way == 2'h2 ? ram_0_81 : _GEN_7657; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9072 = unuse_way == 2'h2 ? ram_0_82 : _GEN_7658; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9073 = unuse_way == 2'h2 ? ram_0_83 : _GEN_7659; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9074 = unuse_way == 2'h2 ? ram_0_84 : _GEN_7660; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9075 = unuse_way == 2'h2 ? ram_0_85 : _GEN_7661; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9076 = unuse_way == 2'h2 ? ram_0_86 : _GEN_7662; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9077 = unuse_way == 2'h2 ? ram_0_87 : _GEN_7663; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9078 = unuse_way == 2'h2 ? ram_0_88 : _GEN_7664; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9079 = unuse_way == 2'h2 ? ram_0_89 : _GEN_7665; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9080 = unuse_way == 2'h2 ? ram_0_90 : _GEN_7666; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9081 = unuse_way == 2'h2 ? ram_0_91 : _GEN_7667; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9082 = unuse_way == 2'h2 ? ram_0_92 : _GEN_7668; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9083 = unuse_way == 2'h2 ? ram_0_93 : _GEN_7669; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9084 = unuse_way == 2'h2 ? ram_0_94 : _GEN_7670; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9085 = unuse_way == 2'h2 ? ram_0_95 : _GEN_7671; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9086 = unuse_way == 2'h2 ? ram_0_96 : _GEN_7672; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9087 = unuse_way == 2'h2 ? ram_0_97 : _GEN_7673; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9088 = unuse_way == 2'h2 ? ram_0_98 : _GEN_7674; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9089 = unuse_way == 2'h2 ? ram_0_99 : _GEN_7675; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9090 = unuse_way == 2'h2 ? ram_0_100 : _GEN_7676; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9091 = unuse_way == 2'h2 ? ram_0_101 : _GEN_7677; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9092 = unuse_way == 2'h2 ? ram_0_102 : _GEN_7678; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9093 = unuse_way == 2'h2 ? ram_0_103 : _GEN_7679; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9094 = unuse_way == 2'h2 ? ram_0_104 : _GEN_7680; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9095 = unuse_way == 2'h2 ? ram_0_105 : _GEN_7681; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9096 = unuse_way == 2'h2 ? ram_0_106 : _GEN_7682; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9097 = unuse_way == 2'h2 ? ram_0_107 : _GEN_7683; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9098 = unuse_way == 2'h2 ? ram_0_108 : _GEN_7684; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9099 = unuse_way == 2'h2 ? ram_0_109 : _GEN_7685; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9100 = unuse_way == 2'h2 ? ram_0_110 : _GEN_7686; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9101 = unuse_way == 2'h2 ? ram_0_111 : _GEN_7687; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9102 = unuse_way == 2'h2 ? ram_0_112 : _GEN_7688; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9103 = unuse_way == 2'h2 ? ram_0_113 : _GEN_7689; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9104 = unuse_way == 2'h2 ? ram_0_114 : _GEN_7690; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9105 = unuse_way == 2'h2 ? ram_0_115 : _GEN_7691; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9106 = unuse_way == 2'h2 ? ram_0_116 : _GEN_7692; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9107 = unuse_way == 2'h2 ? ram_0_117 : _GEN_7693; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9108 = unuse_way == 2'h2 ? ram_0_118 : _GEN_7694; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9109 = unuse_way == 2'h2 ? ram_0_119 : _GEN_7695; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9110 = unuse_way == 2'h2 ? ram_0_120 : _GEN_7696; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9111 = unuse_way == 2'h2 ? ram_0_121 : _GEN_7697; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9112 = unuse_way == 2'h2 ? ram_0_122 : _GEN_7698; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9113 = unuse_way == 2'h2 ? ram_0_123 : _GEN_7699; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9114 = unuse_way == 2'h2 ? ram_0_124 : _GEN_7700; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9115 = unuse_way == 2'h2 ? ram_0_125 : _GEN_7701; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9116 = unuse_way == 2'h2 ? ram_0_126 : _GEN_7702; // @[d_cache.scala 145:40 18:24]
  wire [63:0] _GEN_9117 = unuse_way == 2'h2 ? ram_0_127 : _GEN_7703; // @[d_cache.scala 145:40 18:24]
  wire [31:0] _GEN_9118 = unuse_way == 2'h2 ? tag_0_0 : _GEN_7704; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9119 = unuse_way == 2'h2 ? tag_0_1 : _GEN_7705; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9120 = unuse_way == 2'h2 ? tag_0_2 : _GEN_7706; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9121 = unuse_way == 2'h2 ? tag_0_3 : _GEN_7707; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9122 = unuse_way == 2'h2 ? tag_0_4 : _GEN_7708; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9123 = unuse_way == 2'h2 ? tag_0_5 : _GEN_7709; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9124 = unuse_way == 2'h2 ? tag_0_6 : _GEN_7710; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9125 = unuse_way == 2'h2 ? tag_0_7 : _GEN_7711; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9126 = unuse_way == 2'h2 ? tag_0_8 : _GEN_7712; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9127 = unuse_way == 2'h2 ? tag_0_9 : _GEN_7713; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9128 = unuse_way == 2'h2 ? tag_0_10 : _GEN_7714; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9129 = unuse_way == 2'h2 ? tag_0_11 : _GEN_7715; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9130 = unuse_way == 2'h2 ? tag_0_12 : _GEN_7716; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9131 = unuse_way == 2'h2 ? tag_0_13 : _GEN_7717; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9132 = unuse_way == 2'h2 ? tag_0_14 : _GEN_7718; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9133 = unuse_way == 2'h2 ? tag_0_15 : _GEN_7719; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9134 = unuse_way == 2'h2 ? tag_0_16 : _GEN_7720; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9135 = unuse_way == 2'h2 ? tag_0_17 : _GEN_7721; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9136 = unuse_way == 2'h2 ? tag_0_18 : _GEN_7722; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9137 = unuse_way == 2'h2 ? tag_0_19 : _GEN_7723; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9138 = unuse_way == 2'h2 ? tag_0_20 : _GEN_7724; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9139 = unuse_way == 2'h2 ? tag_0_21 : _GEN_7725; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9140 = unuse_way == 2'h2 ? tag_0_22 : _GEN_7726; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9141 = unuse_way == 2'h2 ? tag_0_23 : _GEN_7727; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9142 = unuse_way == 2'h2 ? tag_0_24 : _GEN_7728; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9143 = unuse_way == 2'h2 ? tag_0_25 : _GEN_7729; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9144 = unuse_way == 2'h2 ? tag_0_26 : _GEN_7730; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9145 = unuse_way == 2'h2 ? tag_0_27 : _GEN_7731; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9146 = unuse_way == 2'h2 ? tag_0_28 : _GEN_7732; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9147 = unuse_way == 2'h2 ? tag_0_29 : _GEN_7733; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9148 = unuse_way == 2'h2 ? tag_0_30 : _GEN_7734; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9149 = unuse_way == 2'h2 ? tag_0_31 : _GEN_7735; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9150 = unuse_way == 2'h2 ? tag_0_32 : _GEN_7736; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9151 = unuse_way == 2'h2 ? tag_0_33 : _GEN_7737; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9152 = unuse_way == 2'h2 ? tag_0_34 : _GEN_7738; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9153 = unuse_way == 2'h2 ? tag_0_35 : _GEN_7739; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9154 = unuse_way == 2'h2 ? tag_0_36 : _GEN_7740; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9155 = unuse_way == 2'h2 ? tag_0_37 : _GEN_7741; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9156 = unuse_way == 2'h2 ? tag_0_38 : _GEN_7742; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9157 = unuse_way == 2'h2 ? tag_0_39 : _GEN_7743; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9158 = unuse_way == 2'h2 ? tag_0_40 : _GEN_7744; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9159 = unuse_way == 2'h2 ? tag_0_41 : _GEN_7745; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9160 = unuse_way == 2'h2 ? tag_0_42 : _GEN_7746; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9161 = unuse_way == 2'h2 ? tag_0_43 : _GEN_7747; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9162 = unuse_way == 2'h2 ? tag_0_44 : _GEN_7748; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9163 = unuse_way == 2'h2 ? tag_0_45 : _GEN_7749; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9164 = unuse_way == 2'h2 ? tag_0_46 : _GEN_7750; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9165 = unuse_way == 2'h2 ? tag_0_47 : _GEN_7751; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9166 = unuse_way == 2'h2 ? tag_0_48 : _GEN_7752; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9167 = unuse_way == 2'h2 ? tag_0_49 : _GEN_7753; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9168 = unuse_way == 2'h2 ? tag_0_50 : _GEN_7754; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9169 = unuse_way == 2'h2 ? tag_0_51 : _GEN_7755; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9170 = unuse_way == 2'h2 ? tag_0_52 : _GEN_7756; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9171 = unuse_way == 2'h2 ? tag_0_53 : _GEN_7757; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9172 = unuse_way == 2'h2 ? tag_0_54 : _GEN_7758; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9173 = unuse_way == 2'h2 ? tag_0_55 : _GEN_7759; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9174 = unuse_way == 2'h2 ? tag_0_56 : _GEN_7760; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9175 = unuse_way == 2'h2 ? tag_0_57 : _GEN_7761; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9176 = unuse_way == 2'h2 ? tag_0_58 : _GEN_7762; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9177 = unuse_way == 2'h2 ? tag_0_59 : _GEN_7763; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9178 = unuse_way == 2'h2 ? tag_0_60 : _GEN_7764; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9179 = unuse_way == 2'h2 ? tag_0_61 : _GEN_7765; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9180 = unuse_way == 2'h2 ? tag_0_62 : _GEN_7766; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9181 = unuse_way == 2'h2 ? tag_0_63 : _GEN_7767; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9182 = unuse_way == 2'h2 ? tag_0_64 : _GEN_7768; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9183 = unuse_way == 2'h2 ? tag_0_65 : _GEN_7769; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9184 = unuse_way == 2'h2 ? tag_0_66 : _GEN_7770; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9185 = unuse_way == 2'h2 ? tag_0_67 : _GEN_7771; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9186 = unuse_way == 2'h2 ? tag_0_68 : _GEN_7772; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9187 = unuse_way == 2'h2 ? tag_0_69 : _GEN_7773; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9188 = unuse_way == 2'h2 ? tag_0_70 : _GEN_7774; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9189 = unuse_way == 2'h2 ? tag_0_71 : _GEN_7775; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9190 = unuse_way == 2'h2 ? tag_0_72 : _GEN_7776; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9191 = unuse_way == 2'h2 ? tag_0_73 : _GEN_7777; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9192 = unuse_way == 2'h2 ? tag_0_74 : _GEN_7778; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9193 = unuse_way == 2'h2 ? tag_0_75 : _GEN_7779; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9194 = unuse_way == 2'h2 ? tag_0_76 : _GEN_7780; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9195 = unuse_way == 2'h2 ? tag_0_77 : _GEN_7781; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9196 = unuse_way == 2'h2 ? tag_0_78 : _GEN_7782; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9197 = unuse_way == 2'h2 ? tag_0_79 : _GEN_7783; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9198 = unuse_way == 2'h2 ? tag_0_80 : _GEN_7784; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9199 = unuse_way == 2'h2 ? tag_0_81 : _GEN_7785; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9200 = unuse_way == 2'h2 ? tag_0_82 : _GEN_7786; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9201 = unuse_way == 2'h2 ? tag_0_83 : _GEN_7787; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9202 = unuse_way == 2'h2 ? tag_0_84 : _GEN_7788; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9203 = unuse_way == 2'h2 ? tag_0_85 : _GEN_7789; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9204 = unuse_way == 2'h2 ? tag_0_86 : _GEN_7790; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9205 = unuse_way == 2'h2 ? tag_0_87 : _GEN_7791; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9206 = unuse_way == 2'h2 ? tag_0_88 : _GEN_7792; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9207 = unuse_way == 2'h2 ? tag_0_89 : _GEN_7793; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9208 = unuse_way == 2'h2 ? tag_0_90 : _GEN_7794; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9209 = unuse_way == 2'h2 ? tag_0_91 : _GEN_7795; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9210 = unuse_way == 2'h2 ? tag_0_92 : _GEN_7796; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9211 = unuse_way == 2'h2 ? tag_0_93 : _GEN_7797; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9212 = unuse_way == 2'h2 ? tag_0_94 : _GEN_7798; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9213 = unuse_way == 2'h2 ? tag_0_95 : _GEN_7799; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9214 = unuse_way == 2'h2 ? tag_0_96 : _GEN_7800; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9215 = unuse_way == 2'h2 ? tag_0_97 : _GEN_7801; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9216 = unuse_way == 2'h2 ? tag_0_98 : _GEN_7802; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9217 = unuse_way == 2'h2 ? tag_0_99 : _GEN_7803; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9218 = unuse_way == 2'h2 ? tag_0_100 : _GEN_7804; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9219 = unuse_way == 2'h2 ? tag_0_101 : _GEN_7805; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9220 = unuse_way == 2'h2 ? tag_0_102 : _GEN_7806; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9221 = unuse_way == 2'h2 ? tag_0_103 : _GEN_7807; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9222 = unuse_way == 2'h2 ? tag_0_104 : _GEN_7808; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9223 = unuse_way == 2'h2 ? tag_0_105 : _GEN_7809; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9224 = unuse_way == 2'h2 ? tag_0_106 : _GEN_7810; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9225 = unuse_way == 2'h2 ? tag_0_107 : _GEN_7811; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9226 = unuse_way == 2'h2 ? tag_0_108 : _GEN_7812; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9227 = unuse_way == 2'h2 ? tag_0_109 : _GEN_7813; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9228 = unuse_way == 2'h2 ? tag_0_110 : _GEN_7814; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9229 = unuse_way == 2'h2 ? tag_0_111 : _GEN_7815; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9230 = unuse_way == 2'h2 ? tag_0_112 : _GEN_7816; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9231 = unuse_way == 2'h2 ? tag_0_113 : _GEN_7817; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9232 = unuse_way == 2'h2 ? tag_0_114 : _GEN_7818; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9233 = unuse_way == 2'h2 ? tag_0_115 : _GEN_7819; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9234 = unuse_way == 2'h2 ? tag_0_116 : _GEN_7820; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9235 = unuse_way == 2'h2 ? tag_0_117 : _GEN_7821; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9236 = unuse_way == 2'h2 ? tag_0_118 : _GEN_7822; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9237 = unuse_way == 2'h2 ? tag_0_119 : _GEN_7823; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9238 = unuse_way == 2'h2 ? tag_0_120 : _GEN_7824; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9239 = unuse_way == 2'h2 ? tag_0_121 : _GEN_7825; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9240 = unuse_way == 2'h2 ? tag_0_122 : _GEN_7826; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9241 = unuse_way == 2'h2 ? tag_0_123 : _GEN_7827; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9242 = unuse_way == 2'h2 ? tag_0_124 : _GEN_7828; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9243 = unuse_way == 2'h2 ? tag_0_125 : _GEN_7829; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9244 = unuse_way == 2'h2 ? tag_0_126 : _GEN_7830; // @[d_cache.scala 145:40 22:24]
  wire [31:0] _GEN_9245 = unuse_way == 2'h2 ? tag_0_127 : _GEN_7831; // @[d_cache.scala 145:40 22:24]
  wire  _GEN_9246 = unuse_way == 2'h2 ? dirty_0_0 : _GEN_7832; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9247 = unuse_way == 2'h2 ? dirty_0_1 : _GEN_7833; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9248 = unuse_way == 2'h2 ? dirty_0_2 : _GEN_7834; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9249 = unuse_way == 2'h2 ? dirty_0_3 : _GEN_7835; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9250 = unuse_way == 2'h2 ? dirty_0_4 : _GEN_7836; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9251 = unuse_way == 2'h2 ? dirty_0_5 : _GEN_7837; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9252 = unuse_way == 2'h2 ? dirty_0_6 : _GEN_7838; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9253 = unuse_way == 2'h2 ? dirty_0_7 : _GEN_7839; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9254 = unuse_way == 2'h2 ? dirty_0_8 : _GEN_7840; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9255 = unuse_way == 2'h2 ? dirty_0_9 : _GEN_7841; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9256 = unuse_way == 2'h2 ? dirty_0_10 : _GEN_7842; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9257 = unuse_way == 2'h2 ? dirty_0_11 : _GEN_7843; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9258 = unuse_way == 2'h2 ? dirty_0_12 : _GEN_7844; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9259 = unuse_way == 2'h2 ? dirty_0_13 : _GEN_7845; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9260 = unuse_way == 2'h2 ? dirty_0_14 : _GEN_7846; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9261 = unuse_way == 2'h2 ? dirty_0_15 : _GEN_7847; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9262 = unuse_way == 2'h2 ? dirty_0_16 : _GEN_7848; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9263 = unuse_way == 2'h2 ? dirty_0_17 : _GEN_7849; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9264 = unuse_way == 2'h2 ? dirty_0_18 : _GEN_7850; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9265 = unuse_way == 2'h2 ? dirty_0_19 : _GEN_7851; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9266 = unuse_way == 2'h2 ? dirty_0_20 : _GEN_7852; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9267 = unuse_way == 2'h2 ? dirty_0_21 : _GEN_7853; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9268 = unuse_way == 2'h2 ? dirty_0_22 : _GEN_7854; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9269 = unuse_way == 2'h2 ? dirty_0_23 : _GEN_7855; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9270 = unuse_way == 2'h2 ? dirty_0_24 : _GEN_7856; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9271 = unuse_way == 2'h2 ? dirty_0_25 : _GEN_7857; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9272 = unuse_way == 2'h2 ? dirty_0_26 : _GEN_7858; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9273 = unuse_way == 2'h2 ? dirty_0_27 : _GEN_7859; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9274 = unuse_way == 2'h2 ? dirty_0_28 : _GEN_7860; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9275 = unuse_way == 2'h2 ? dirty_0_29 : _GEN_7861; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9276 = unuse_way == 2'h2 ? dirty_0_30 : _GEN_7862; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9277 = unuse_way == 2'h2 ? dirty_0_31 : _GEN_7863; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9278 = unuse_way == 2'h2 ? dirty_0_32 : _GEN_7864; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9279 = unuse_way == 2'h2 ? dirty_0_33 : _GEN_7865; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9280 = unuse_way == 2'h2 ? dirty_0_34 : _GEN_7866; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9281 = unuse_way == 2'h2 ? dirty_0_35 : _GEN_7867; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9282 = unuse_way == 2'h2 ? dirty_0_36 : _GEN_7868; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9283 = unuse_way == 2'h2 ? dirty_0_37 : _GEN_7869; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9284 = unuse_way == 2'h2 ? dirty_0_38 : _GEN_7870; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9285 = unuse_way == 2'h2 ? dirty_0_39 : _GEN_7871; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9286 = unuse_way == 2'h2 ? dirty_0_40 : _GEN_7872; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9287 = unuse_way == 2'h2 ? dirty_0_41 : _GEN_7873; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9288 = unuse_way == 2'h2 ? dirty_0_42 : _GEN_7874; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9289 = unuse_way == 2'h2 ? dirty_0_43 : _GEN_7875; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9290 = unuse_way == 2'h2 ? dirty_0_44 : _GEN_7876; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9291 = unuse_way == 2'h2 ? dirty_0_45 : _GEN_7877; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9292 = unuse_way == 2'h2 ? dirty_0_46 : _GEN_7878; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9293 = unuse_way == 2'h2 ? dirty_0_47 : _GEN_7879; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9294 = unuse_way == 2'h2 ? dirty_0_48 : _GEN_7880; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9295 = unuse_way == 2'h2 ? dirty_0_49 : _GEN_7881; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9296 = unuse_way == 2'h2 ? dirty_0_50 : _GEN_7882; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9297 = unuse_way == 2'h2 ? dirty_0_51 : _GEN_7883; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9298 = unuse_way == 2'h2 ? dirty_0_52 : _GEN_7884; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9299 = unuse_way == 2'h2 ? dirty_0_53 : _GEN_7885; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9300 = unuse_way == 2'h2 ? dirty_0_54 : _GEN_7886; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9301 = unuse_way == 2'h2 ? dirty_0_55 : _GEN_7887; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9302 = unuse_way == 2'h2 ? dirty_0_56 : _GEN_7888; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9303 = unuse_way == 2'h2 ? dirty_0_57 : _GEN_7889; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9304 = unuse_way == 2'h2 ? dirty_0_58 : _GEN_7890; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9305 = unuse_way == 2'h2 ? dirty_0_59 : _GEN_7891; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9306 = unuse_way == 2'h2 ? dirty_0_60 : _GEN_7892; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9307 = unuse_way == 2'h2 ? dirty_0_61 : _GEN_7893; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9308 = unuse_way == 2'h2 ? dirty_0_62 : _GEN_7894; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9309 = unuse_way == 2'h2 ? dirty_0_63 : _GEN_7895; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9310 = unuse_way == 2'h2 ? dirty_0_64 : _GEN_7896; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9311 = unuse_way == 2'h2 ? dirty_0_65 : _GEN_7897; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9312 = unuse_way == 2'h2 ? dirty_0_66 : _GEN_7898; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9313 = unuse_way == 2'h2 ? dirty_0_67 : _GEN_7899; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9314 = unuse_way == 2'h2 ? dirty_0_68 : _GEN_7900; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9315 = unuse_way == 2'h2 ? dirty_0_69 : _GEN_7901; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9316 = unuse_way == 2'h2 ? dirty_0_70 : _GEN_7902; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9317 = unuse_way == 2'h2 ? dirty_0_71 : _GEN_7903; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9318 = unuse_way == 2'h2 ? dirty_0_72 : _GEN_7904; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9319 = unuse_way == 2'h2 ? dirty_0_73 : _GEN_7905; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9320 = unuse_way == 2'h2 ? dirty_0_74 : _GEN_7906; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9321 = unuse_way == 2'h2 ? dirty_0_75 : _GEN_7907; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9322 = unuse_way == 2'h2 ? dirty_0_76 : _GEN_7908; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9323 = unuse_way == 2'h2 ? dirty_0_77 : _GEN_7909; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9324 = unuse_way == 2'h2 ? dirty_0_78 : _GEN_7910; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9325 = unuse_way == 2'h2 ? dirty_0_79 : _GEN_7911; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9326 = unuse_way == 2'h2 ? dirty_0_80 : _GEN_7912; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9327 = unuse_way == 2'h2 ? dirty_0_81 : _GEN_7913; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9328 = unuse_way == 2'h2 ? dirty_0_82 : _GEN_7914; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9329 = unuse_way == 2'h2 ? dirty_0_83 : _GEN_7915; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9330 = unuse_way == 2'h2 ? dirty_0_84 : _GEN_7916; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9331 = unuse_way == 2'h2 ? dirty_0_85 : _GEN_7917; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9332 = unuse_way == 2'h2 ? dirty_0_86 : _GEN_7918; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9333 = unuse_way == 2'h2 ? dirty_0_87 : _GEN_7919; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9334 = unuse_way == 2'h2 ? dirty_0_88 : _GEN_7920; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9335 = unuse_way == 2'h2 ? dirty_0_89 : _GEN_7921; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9336 = unuse_way == 2'h2 ? dirty_0_90 : _GEN_7922; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9337 = unuse_way == 2'h2 ? dirty_0_91 : _GEN_7923; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9338 = unuse_way == 2'h2 ? dirty_0_92 : _GEN_7924; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9339 = unuse_way == 2'h2 ? dirty_0_93 : _GEN_7925; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9340 = unuse_way == 2'h2 ? dirty_0_94 : _GEN_7926; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9341 = unuse_way == 2'h2 ? dirty_0_95 : _GEN_7927; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9342 = unuse_way == 2'h2 ? dirty_0_96 : _GEN_7928; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9343 = unuse_way == 2'h2 ? dirty_0_97 : _GEN_7929; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9344 = unuse_way == 2'h2 ? dirty_0_98 : _GEN_7930; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9345 = unuse_way == 2'h2 ? dirty_0_99 : _GEN_7931; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9346 = unuse_way == 2'h2 ? dirty_0_100 : _GEN_7932; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9347 = unuse_way == 2'h2 ? dirty_0_101 : _GEN_7933; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9348 = unuse_way == 2'h2 ? dirty_0_102 : _GEN_7934; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9349 = unuse_way == 2'h2 ? dirty_0_103 : _GEN_7935; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9350 = unuse_way == 2'h2 ? dirty_0_104 : _GEN_7936; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9351 = unuse_way == 2'h2 ? dirty_0_105 : _GEN_7937; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9352 = unuse_way == 2'h2 ? dirty_0_106 : _GEN_7938; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9353 = unuse_way == 2'h2 ? dirty_0_107 : _GEN_7939; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9354 = unuse_way == 2'h2 ? dirty_0_108 : _GEN_7940; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9355 = unuse_way == 2'h2 ? dirty_0_109 : _GEN_7941; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9356 = unuse_way == 2'h2 ? dirty_0_110 : _GEN_7942; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9357 = unuse_way == 2'h2 ? dirty_0_111 : _GEN_7943; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9358 = unuse_way == 2'h2 ? dirty_0_112 : _GEN_7944; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9359 = unuse_way == 2'h2 ? dirty_0_113 : _GEN_7945; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9360 = unuse_way == 2'h2 ? dirty_0_114 : _GEN_7946; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9361 = unuse_way == 2'h2 ? dirty_0_115 : _GEN_7947; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9362 = unuse_way == 2'h2 ? dirty_0_116 : _GEN_7948; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9363 = unuse_way == 2'h2 ? dirty_0_117 : _GEN_7949; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9364 = unuse_way == 2'h2 ? dirty_0_118 : _GEN_7950; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9365 = unuse_way == 2'h2 ? dirty_0_119 : _GEN_7951; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9366 = unuse_way == 2'h2 ? dirty_0_120 : _GEN_7952; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9367 = unuse_way == 2'h2 ? dirty_0_121 : _GEN_7953; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9368 = unuse_way == 2'h2 ? dirty_0_122 : _GEN_7954; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9369 = unuse_way == 2'h2 ? dirty_0_123 : _GEN_7955; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9370 = unuse_way == 2'h2 ? dirty_0_124 : _GEN_7956; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9371 = unuse_way == 2'h2 ? dirty_0_125 : _GEN_7957; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9372 = unuse_way == 2'h2 ? dirty_0_126 : _GEN_7958; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9373 = unuse_way == 2'h2 ? dirty_0_127 : _GEN_7959; // @[d_cache.scala 145:40 26:26]
  wire  _GEN_9374 = unuse_way == 2'h2 ? valid_0_0 : _GEN_7960; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9375 = unuse_way == 2'h2 ? valid_0_1 : _GEN_7961; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9376 = unuse_way == 2'h2 ? valid_0_2 : _GEN_7962; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9377 = unuse_way == 2'h2 ? valid_0_3 : _GEN_7963; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9378 = unuse_way == 2'h2 ? valid_0_4 : _GEN_7964; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9379 = unuse_way == 2'h2 ? valid_0_5 : _GEN_7965; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9380 = unuse_way == 2'h2 ? valid_0_6 : _GEN_7966; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9381 = unuse_way == 2'h2 ? valid_0_7 : _GEN_7967; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9382 = unuse_way == 2'h2 ? valid_0_8 : _GEN_7968; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9383 = unuse_way == 2'h2 ? valid_0_9 : _GEN_7969; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9384 = unuse_way == 2'h2 ? valid_0_10 : _GEN_7970; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9385 = unuse_way == 2'h2 ? valid_0_11 : _GEN_7971; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9386 = unuse_way == 2'h2 ? valid_0_12 : _GEN_7972; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9387 = unuse_way == 2'h2 ? valid_0_13 : _GEN_7973; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9388 = unuse_way == 2'h2 ? valid_0_14 : _GEN_7974; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9389 = unuse_way == 2'h2 ? valid_0_15 : _GEN_7975; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9390 = unuse_way == 2'h2 ? valid_0_16 : _GEN_7976; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9391 = unuse_way == 2'h2 ? valid_0_17 : _GEN_7977; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9392 = unuse_way == 2'h2 ? valid_0_18 : _GEN_7978; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9393 = unuse_way == 2'h2 ? valid_0_19 : _GEN_7979; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9394 = unuse_way == 2'h2 ? valid_0_20 : _GEN_7980; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9395 = unuse_way == 2'h2 ? valid_0_21 : _GEN_7981; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9396 = unuse_way == 2'h2 ? valid_0_22 : _GEN_7982; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9397 = unuse_way == 2'h2 ? valid_0_23 : _GEN_7983; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9398 = unuse_way == 2'h2 ? valid_0_24 : _GEN_7984; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9399 = unuse_way == 2'h2 ? valid_0_25 : _GEN_7985; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9400 = unuse_way == 2'h2 ? valid_0_26 : _GEN_7986; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9401 = unuse_way == 2'h2 ? valid_0_27 : _GEN_7987; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9402 = unuse_way == 2'h2 ? valid_0_28 : _GEN_7988; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9403 = unuse_way == 2'h2 ? valid_0_29 : _GEN_7989; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9404 = unuse_way == 2'h2 ? valid_0_30 : _GEN_7990; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9405 = unuse_way == 2'h2 ? valid_0_31 : _GEN_7991; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9406 = unuse_way == 2'h2 ? valid_0_32 : _GEN_7992; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9407 = unuse_way == 2'h2 ? valid_0_33 : _GEN_7993; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9408 = unuse_way == 2'h2 ? valid_0_34 : _GEN_7994; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9409 = unuse_way == 2'h2 ? valid_0_35 : _GEN_7995; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9410 = unuse_way == 2'h2 ? valid_0_36 : _GEN_7996; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9411 = unuse_way == 2'h2 ? valid_0_37 : _GEN_7997; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9412 = unuse_way == 2'h2 ? valid_0_38 : _GEN_7998; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9413 = unuse_way == 2'h2 ? valid_0_39 : _GEN_7999; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9414 = unuse_way == 2'h2 ? valid_0_40 : _GEN_8000; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9415 = unuse_way == 2'h2 ? valid_0_41 : _GEN_8001; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9416 = unuse_way == 2'h2 ? valid_0_42 : _GEN_8002; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9417 = unuse_way == 2'h2 ? valid_0_43 : _GEN_8003; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9418 = unuse_way == 2'h2 ? valid_0_44 : _GEN_8004; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9419 = unuse_way == 2'h2 ? valid_0_45 : _GEN_8005; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9420 = unuse_way == 2'h2 ? valid_0_46 : _GEN_8006; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9421 = unuse_way == 2'h2 ? valid_0_47 : _GEN_8007; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9422 = unuse_way == 2'h2 ? valid_0_48 : _GEN_8008; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9423 = unuse_way == 2'h2 ? valid_0_49 : _GEN_8009; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9424 = unuse_way == 2'h2 ? valid_0_50 : _GEN_8010; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9425 = unuse_way == 2'h2 ? valid_0_51 : _GEN_8011; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9426 = unuse_way == 2'h2 ? valid_0_52 : _GEN_8012; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9427 = unuse_way == 2'h2 ? valid_0_53 : _GEN_8013; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9428 = unuse_way == 2'h2 ? valid_0_54 : _GEN_8014; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9429 = unuse_way == 2'h2 ? valid_0_55 : _GEN_8015; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9430 = unuse_way == 2'h2 ? valid_0_56 : _GEN_8016; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9431 = unuse_way == 2'h2 ? valid_0_57 : _GEN_8017; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9432 = unuse_way == 2'h2 ? valid_0_58 : _GEN_8018; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9433 = unuse_way == 2'h2 ? valid_0_59 : _GEN_8019; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9434 = unuse_way == 2'h2 ? valid_0_60 : _GEN_8020; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9435 = unuse_way == 2'h2 ? valid_0_61 : _GEN_8021; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9436 = unuse_way == 2'h2 ? valid_0_62 : _GEN_8022; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9437 = unuse_way == 2'h2 ? valid_0_63 : _GEN_8023; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9438 = unuse_way == 2'h2 ? valid_0_64 : _GEN_8024; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9439 = unuse_way == 2'h2 ? valid_0_65 : _GEN_8025; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9440 = unuse_way == 2'h2 ? valid_0_66 : _GEN_8026; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9441 = unuse_way == 2'h2 ? valid_0_67 : _GEN_8027; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9442 = unuse_way == 2'h2 ? valid_0_68 : _GEN_8028; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9443 = unuse_way == 2'h2 ? valid_0_69 : _GEN_8029; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9444 = unuse_way == 2'h2 ? valid_0_70 : _GEN_8030; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9445 = unuse_way == 2'h2 ? valid_0_71 : _GEN_8031; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9446 = unuse_way == 2'h2 ? valid_0_72 : _GEN_8032; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9447 = unuse_way == 2'h2 ? valid_0_73 : _GEN_8033; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9448 = unuse_way == 2'h2 ? valid_0_74 : _GEN_8034; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9449 = unuse_way == 2'h2 ? valid_0_75 : _GEN_8035; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9450 = unuse_way == 2'h2 ? valid_0_76 : _GEN_8036; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9451 = unuse_way == 2'h2 ? valid_0_77 : _GEN_8037; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9452 = unuse_way == 2'h2 ? valid_0_78 : _GEN_8038; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9453 = unuse_way == 2'h2 ? valid_0_79 : _GEN_8039; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9454 = unuse_way == 2'h2 ? valid_0_80 : _GEN_8040; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9455 = unuse_way == 2'h2 ? valid_0_81 : _GEN_8041; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9456 = unuse_way == 2'h2 ? valid_0_82 : _GEN_8042; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9457 = unuse_way == 2'h2 ? valid_0_83 : _GEN_8043; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9458 = unuse_way == 2'h2 ? valid_0_84 : _GEN_8044; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9459 = unuse_way == 2'h2 ? valid_0_85 : _GEN_8045; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9460 = unuse_way == 2'h2 ? valid_0_86 : _GEN_8046; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9461 = unuse_way == 2'h2 ? valid_0_87 : _GEN_8047; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9462 = unuse_way == 2'h2 ? valid_0_88 : _GEN_8048; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9463 = unuse_way == 2'h2 ? valid_0_89 : _GEN_8049; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9464 = unuse_way == 2'h2 ? valid_0_90 : _GEN_8050; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9465 = unuse_way == 2'h2 ? valid_0_91 : _GEN_8051; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9466 = unuse_way == 2'h2 ? valid_0_92 : _GEN_8052; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9467 = unuse_way == 2'h2 ? valid_0_93 : _GEN_8053; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9468 = unuse_way == 2'h2 ? valid_0_94 : _GEN_8054; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9469 = unuse_way == 2'h2 ? valid_0_95 : _GEN_8055; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9470 = unuse_way == 2'h2 ? valid_0_96 : _GEN_8056; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9471 = unuse_way == 2'h2 ? valid_0_97 : _GEN_8057; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9472 = unuse_way == 2'h2 ? valid_0_98 : _GEN_8058; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9473 = unuse_way == 2'h2 ? valid_0_99 : _GEN_8059; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9474 = unuse_way == 2'h2 ? valid_0_100 : _GEN_8060; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9475 = unuse_way == 2'h2 ? valid_0_101 : _GEN_8061; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9476 = unuse_way == 2'h2 ? valid_0_102 : _GEN_8062; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9477 = unuse_way == 2'h2 ? valid_0_103 : _GEN_8063; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9478 = unuse_way == 2'h2 ? valid_0_104 : _GEN_8064; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9479 = unuse_way == 2'h2 ? valid_0_105 : _GEN_8065; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9480 = unuse_way == 2'h2 ? valid_0_106 : _GEN_8066; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9481 = unuse_way == 2'h2 ? valid_0_107 : _GEN_8067; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9482 = unuse_way == 2'h2 ? valid_0_108 : _GEN_8068; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9483 = unuse_way == 2'h2 ? valid_0_109 : _GEN_8069; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9484 = unuse_way == 2'h2 ? valid_0_110 : _GEN_8070; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9485 = unuse_way == 2'h2 ? valid_0_111 : _GEN_8071; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9486 = unuse_way == 2'h2 ? valid_0_112 : _GEN_8072; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9487 = unuse_way == 2'h2 ? valid_0_113 : _GEN_8073; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9488 = unuse_way == 2'h2 ? valid_0_114 : _GEN_8074; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9489 = unuse_way == 2'h2 ? valid_0_115 : _GEN_8075; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9490 = unuse_way == 2'h2 ? valid_0_116 : _GEN_8076; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9491 = unuse_way == 2'h2 ? valid_0_117 : _GEN_8077; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9492 = unuse_way == 2'h2 ? valid_0_118 : _GEN_8078; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9493 = unuse_way == 2'h2 ? valid_0_119 : _GEN_8079; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9494 = unuse_way == 2'h2 ? valid_0_120 : _GEN_8080; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9495 = unuse_way == 2'h2 ? valid_0_121 : _GEN_8081; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9496 = unuse_way == 2'h2 ? valid_0_122 : _GEN_8082; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9497 = unuse_way == 2'h2 ? valid_0_123 : _GEN_8083; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9498 = unuse_way == 2'h2 ? valid_0_124 : _GEN_8084; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9499 = unuse_way == 2'h2 ? valid_0_125 : _GEN_8085; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9500 = unuse_way == 2'h2 ? valid_0_126 : _GEN_8086; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9501 = unuse_way == 2'h2 ? valid_0_127 : _GEN_8087; // @[d_cache.scala 145:40 24:26]
  wire  _GEN_9502 = unuse_way == 2'h2 ? dirty_1_0 : _GEN_8346; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9503 = unuse_way == 2'h2 ? dirty_1_1 : _GEN_8347; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9504 = unuse_way == 2'h2 ? dirty_1_2 : _GEN_8348; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9505 = unuse_way == 2'h2 ? dirty_1_3 : _GEN_8349; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9506 = unuse_way == 2'h2 ? dirty_1_4 : _GEN_8350; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9507 = unuse_way == 2'h2 ? dirty_1_5 : _GEN_8351; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9508 = unuse_way == 2'h2 ? dirty_1_6 : _GEN_8352; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9509 = unuse_way == 2'h2 ? dirty_1_7 : _GEN_8353; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9510 = unuse_way == 2'h2 ? dirty_1_8 : _GEN_8354; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9511 = unuse_way == 2'h2 ? dirty_1_9 : _GEN_8355; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9512 = unuse_way == 2'h2 ? dirty_1_10 : _GEN_8356; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9513 = unuse_way == 2'h2 ? dirty_1_11 : _GEN_8357; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9514 = unuse_way == 2'h2 ? dirty_1_12 : _GEN_8358; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9515 = unuse_way == 2'h2 ? dirty_1_13 : _GEN_8359; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9516 = unuse_way == 2'h2 ? dirty_1_14 : _GEN_8360; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9517 = unuse_way == 2'h2 ? dirty_1_15 : _GEN_8361; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9518 = unuse_way == 2'h2 ? dirty_1_16 : _GEN_8362; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9519 = unuse_way == 2'h2 ? dirty_1_17 : _GEN_8363; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9520 = unuse_way == 2'h2 ? dirty_1_18 : _GEN_8364; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9521 = unuse_way == 2'h2 ? dirty_1_19 : _GEN_8365; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9522 = unuse_way == 2'h2 ? dirty_1_20 : _GEN_8366; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9523 = unuse_way == 2'h2 ? dirty_1_21 : _GEN_8367; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9524 = unuse_way == 2'h2 ? dirty_1_22 : _GEN_8368; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9525 = unuse_way == 2'h2 ? dirty_1_23 : _GEN_8369; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9526 = unuse_way == 2'h2 ? dirty_1_24 : _GEN_8370; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9527 = unuse_way == 2'h2 ? dirty_1_25 : _GEN_8371; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9528 = unuse_way == 2'h2 ? dirty_1_26 : _GEN_8372; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9529 = unuse_way == 2'h2 ? dirty_1_27 : _GEN_8373; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9530 = unuse_way == 2'h2 ? dirty_1_28 : _GEN_8374; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9531 = unuse_way == 2'h2 ? dirty_1_29 : _GEN_8375; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9532 = unuse_way == 2'h2 ? dirty_1_30 : _GEN_8376; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9533 = unuse_way == 2'h2 ? dirty_1_31 : _GEN_8377; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9534 = unuse_way == 2'h2 ? dirty_1_32 : _GEN_8378; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9535 = unuse_way == 2'h2 ? dirty_1_33 : _GEN_8379; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9536 = unuse_way == 2'h2 ? dirty_1_34 : _GEN_8380; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9537 = unuse_way == 2'h2 ? dirty_1_35 : _GEN_8381; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9538 = unuse_way == 2'h2 ? dirty_1_36 : _GEN_8382; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9539 = unuse_way == 2'h2 ? dirty_1_37 : _GEN_8383; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9540 = unuse_way == 2'h2 ? dirty_1_38 : _GEN_8384; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9541 = unuse_way == 2'h2 ? dirty_1_39 : _GEN_8385; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9542 = unuse_way == 2'h2 ? dirty_1_40 : _GEN_8386; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9543 = unuse_way == 2'h2 ? dirty_1_41 : _GEN_8387; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9544 = unuse_way == 2'h2 ? dirty_1_42 : _GEN_8388; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9545 = unuse_way == 2'h2 ? dirty_1_43 : _GEN_8389; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9546 = unuse_way == 2'h2 ? dirty_1_44 : _GEN_8390; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9547 = unuse_way == 2'h2 ? dirty_1_45 : _GEN_8391; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9548 = unuse_way == 2'h2 ? dirty_1_46 : _GEN_8392; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9549 = unuse_way == 2'h2 ? dirty_1_47 : _GEN_8393; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9550 = unuse_way == 2'h2 ? dirty_1_48 : _GEN_8394; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9551 = unuse_way == 2'h2 ? dirty_1_49 : _GEN_8395; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9552 = unuse_way == 2'h2 ? dirty_1_50 : _GEN_8396; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9553 = unuse_way == 2'h2 ? dirty_1_51 : _GEN_8397; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9554 = unuse_way == 2'h2 ? dirty_1_52 : _GEN_8398; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9555 = unuse_way == 2'h2 ? dirty_1_53 : _GEN_8399; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9556 = unuse_way == 2'h2 ? dirty_1_54 : _GEN_8400; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9557 = unuse_way == 2'h2 ? dirty_1_55 : _GEN_8401; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9558 = unuse_way == 2'h2 ? dirty_1_56 : _GEN_8402; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9559 = unuse_way == 2'h2 ? dirty_1_57 : _GEN_8403; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9560 = unuse_way == 2'h2 ? dirty_1_58 : _GEN_8404; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9561 = unuse_way == 2'h2 ? dirty_1_59 : _GEN_8405; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9562 = unuse_way == 2'h2 ? dirty_1_60 : _GEN_8406; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9563 = unuse_way == 2'h2 ? dirty_1_61 : _GEN_8407; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9564 = unuse_way == 2'h2 ? dirty_1_62 : _GEN_8408; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9565 = unuse_way == 2'h2 ? dirty_1_63 : _GEN_8409; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9566 = unuse_way == 2'h2 ? dirty_1_64 : _GEN_8410; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9567 = unuse_way == 2'h2 ? dirty_1_65 : _GEN_8411; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9568 = unuse_way == 2'h2 ? dirty_1_66 : _GEN_8412; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9569 = unuse_way == 2'h2 ? dirty_1_67 : _GEN_8413; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9570 = unuse_way == 2'h2 ? dirty_1_68 : _GEN_8414; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9571 = unuse_way == 2'h2 ? dirty_1_69 : _GEN_8415; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9572 = unuse_way == 2'h2 ? dirty_1_70 : _GEN_8416; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9573 = unuse_way == 2'h2 ? dirty_1_71 : _GEN_8417; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9574 = unuse_way == 2'h2 ? dirty_1_72 : _GEN_8418; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9575 = unuse_way == 2'h2 ? dirty_1_73 : _GEN_8419; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9576 = unuse_way == 2'h2 ? dirty_1_74 : _GEN_8420; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9577 = unuse_way == 2'h2 ? dirty_1_75 : _GEN_8421; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9578 = unuse_way == 2'h2 ? dirty_1_76 : _GEN_8422; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9579 = unuse_way == 2'h2 ? dirty_1_77 : _GEN_8423; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9580 = unuse_way == 2'h2 ? dirty_1_78 : _GEN_8424; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9581 = unuse_way == 2'h2 ? dirty_1_79 : _GEN_8425; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9582 = unuse_way == 2'h2 ? dirty_1_80 : _GEN_8426; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9583 = unuse_way == 2'h2 ? dirty_1_81 : _GEN_8427; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9584 = unuse_way == 2'h2 ? dirty_1_82 : _GEN_8428; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9585 = unuse_way == 2'h2 ? dirty_1_83 : _GEN_8429; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9586 = unuse_way == 2'h2 ? dirty_1_84 : _GEN_8430; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9587 = unuse_way == 2'h2 ? dirty_1_85 : _GEN_8431; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9588 = unuse_way == 2'h2 ? dirty_1_86 : _GEN_8432; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9589 = unuse_way == 2'h2 ? dirty_1_87 : _GEN_8433; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9590 = unuse_way == 2'h2 ? dirty_1_88 : _GEN_8434; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9591 = unuse_way == 2'h2 ? dirty_1_89 : _GEN_8435; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9592 = unuse_way == 2'h2 ? dirty_1_90 : _GEN_8436; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9593 = unuse_way == 2'h2 ? dirty_1_91 : _GEN_8437; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9594 = unuse_way == 2'h2 ? dirty_1_92 : _GEN_8438; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9595 = unuse_way == 2'h2 ? dirty_1_93 : _GEN_8439; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9596 = unuse_way == 2'h2 ? dirty_1_94 : _GEN_8440; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9597 = unuse_way == 2'h2 ? dirty_1_95 : _GEN_8441; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9598 = unuse_way == 2'h2 ? dirty_1_96 : _GEN_8442; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9599 = unuse_way == 2'h2 ? dirty_1_97 : _GEN_8443; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9600 = unuse_way == 2'h2 ? dirty_1_98 : _GEN_8444; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9601 = unuse_way == 2'h2 ? dirty_1_99 : _GEN_8445; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9602 = unuse_way == 2'h2 ? dirty_1_100 : _GEN_8446; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9603 = unuse_way == 2'h2 ? dirty_1_101 : _GEN_8447; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9604 = unuse_way == 2'h2 ? dirty_1_102 : _GEN_8448; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9605 = unuse_way == 2'h2 ? dirty_1_103 : _GEN_8449; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9606 = unuse_way == 2'h2 ? dirty_1_104 : _GEN_8450; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9607 = unuse_way == 2'h2 ? dirty_1_105 : _GEN_8451; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9608 = unuse_way == 2'h2 ? dirty_1_106 : _GEN_8452; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9609 = unuse_way == 2'h2 ? dirty_1_107 : _GEN_8453; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9610 = unuse_way == 2'h2 ? dirty_1_108 : _GEN_8454; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9611 = unuse_way == 2'h2 ? dirty_1_109 : _GEN_8455; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9612 = unuse_way == 2'h2 ? dirty_1_110 : _GEN_8456; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9613 = unuse_way == 2'h2 ? dirty_1_111 : _GEN_8457; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9614 = unuse_way == 2'h2 ? dirty_1_112 : _GEN_8458; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9615 = unuse_way == 2'h2 ? dirty_1_113 : _GEN_8459; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9616 = unuse_way == 2'h2 ? dirty_1_114 : _GEN_8460; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9617 = unuse_way == 2'h2 ? dirty_1_115 : _GEN_8461; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9618 = unuse_way == 2'h2 ? dirty_1_116 : _GEN_8462; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9619 = unuse_way == 2'h2 ? dirty_1_117 : _GEN_8463; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9620 = unuse_way == 2'h2 ? dirty_1_118 : _GEN_8464; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9621 = unuse_way == 2'h2 ? dirty_1_119 : _GEN_8465; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9622 = unuse_way == 2'h2 ? dirty_1_120 : _GEN_8466; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9623 = unuse_way == 2'h2 ? dirty_1_121 : _GEN_8467; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9624 = unuse_way == 2'h2 ? dirty_1_122 : _GEN_8468; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9625 = unuse_way == 2'h2 ? dirty_1_123 : _GEN_8469; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9626 = unuse_way == 2'h2 ? dirty_1_124 : _GEN_8470; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9627 = unuse_way == 2'h2 ? dirty_1_125 : _GEN_8471; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9628 = unuse_way == 2'h2 ? dirty_1_126 : _GEN_8472; // @[d_cache.scala 145:40 27:26]
  wire  _GEN_9629 = unuse_way == 2'h2 ? dirty_1_127 : _GEN_8473; // @[d_cache.scala 145:40 27:26]
  wire [2:0] _GEN_9630 = unuse_way == 2'h1 ? 3'h7 : _GEN_8602; // @[d_cache.scala 139:34 140:23]
  wire [63:0] _GEN_9631 = unuse_way == 2'h1 ? _GEN_3214 : _GEN_8990; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9632 = unuse_way == 2'h1 ? _GEN_3215 : _GEN_8991; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9633 = unuse_way == 2'h1 ? _GEN_3216 : _GEN_8992; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9634 = unuse_way == 2'h1 ? _GEN_3217 : _GEN_8993; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9635 = unuse_way == 2'h1 ? _GEN_3218 : _GEN_8994; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9636 = unuse_way == 2'h1 ? _GEN_3219 : _GEN_8995; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9637 = unuse_way == 2'h1 ? _GEN_3220 : _GEN_8996; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9638 = unuse_way == 2'h1 ? _GEN_3221 : _GEN_8997; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9639 = unuse_way == 2'h1 ? _GEN_3222 : _GEN_8998; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9640 = unuse_way == 2'h1 ? _GEN_3223 : _GEN_8999; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9641 = unuse_way == 2'h1 ? _GEN_3224 : _GEN_9000; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9642 = unuse_way == 2'h1 ? _GEN_3225 : _GEN_9001; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9643 = unuse_way == 2'h1 ? _GEN_3226 : _GEN_9002; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9644 = unuse_way == 2'h1 ? _GEN_3227 : _GEN_9003; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9645 = unuse_way == 2'h1 ? _GEN_3228 : _GEN_9004; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9646 = unuse_way == 2'h1 ? _GEN_3229 : _GEN_9005; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9647 = unuse_way == 2'h1 ? _GEN_3230 : _GEN_9006; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9648 = unuse_way == 2'h1 ? _GEN_3231 : _GEN_9007; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9649 = unuse_way == 2'h1 ? _GEN_3232 : _GEN_9008; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9650 = unuse_way == 2'h1 ? _GEN_3233 : _GEN_9009; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9651 = unuse_way == 2'h1 ? _GEN_3234 : _GEN_9010; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9652 = unuse_way == 2'h1 ? _GEN_3235 : _GEN_9011; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9653 = unuse_way == 2'h1 ? _GEN_3236 : _GEN_9012; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9654 = unuse_way == 2'h1 ? _GEN_3237 : _GEN_9013; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9655 = unuse_way == 2'h1 ? _GEN_3238 : _GEN_9014; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9656 = unuse_way == 2'h1 ? _GEN_3239 : _GEN_9015; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9657 = unuse_way == 2'h1 ? _GEN_3240 : _GEN_9016; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9658 = unuse_way == 2'h1 ? _GEN_3241 : _GEN_9017; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9659 = unuse_way == 2'h1 ? _GEN_3242 : _GEN_9018; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9660 = unuse_way == 2'h1 ? _GEN_3243 : _GEN_9019; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9661 = unuse_way == 2'h1 ? _GEN_3244 : _GEN_9020; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9662 = unuse_way == 2'h1 ? _GEN_3245 : _GEN_9021; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9663 = unuse_way == 2'h1 ? _GEN_3246 : _GEN_9022; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9664 = unuse_way == 2'h1 ? _GEN_3247 : _GEN_9023; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9665 = unuse_way == 2'h1 ? _GEN_3248 : _GEN_9024; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9666 = unuse_way == 2'h1 ? _GEN_3249 : _GEN_9025; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9667 = unuse_way == 2'h1 ? _GEN_3250 : _GEN_9026; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9668 = unuse_way == 2'h1 ? _GEN_3251 : _GEN_9027; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9669 = unuse_way == 2'h1 ? _GEN_3252 : _GEN_9028; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9670 = unuse_way == 2'h1 ? _GEN_3253 : _GEN_9029; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9671 = unuse_way == 2'h1 ? _GEN_3254 : _GEN_9030; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9672 = unuse_way == 2'h1 ? _GEN_3255 : _GEN_9031; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9673 = unuse_way == 2'h1 ? _GEN_3256 : _GEN_9032; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9674 = unuse_way == 2'h1 ? _GEN_3257 : _GEN_9033; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9675 = unuse_way == 2'h1 ? _GEN_3258 : _GEN_9034; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9676 = unuse_way == 2'h1 ? _GEN_3259 : _GEN_9035; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9677 = unuse_way == 2'h1 ? _GEN_3260 : _GEN_9036; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9678 = unuse_way == 2'h1 ? _GEN_3261 : _GEN_9037; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9679 = unuse_way == 2'h1 ? _GEN_3262 : _GEN_9038; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9680 = unuse_way == 2'h1 ? _GEN_3263 : _GEN_9039; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9681 = unuse_way == 2'h1 ? _GEN_3264 : _GEN_9040; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9682 = unuse_way == 2'h1 ? _GEN_3265 : _GEN_9041; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9683 = unuse_way == 2'h1 ? _GEN_3266 : _GEN_9042; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9684 = unuse_way == 2'h1 ? _GEN_3267 : _GEN_9043; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9685 = unuse_way == 2'h1 ? _GEN_3268 : _GEN_9044; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9686 = unuse_way == 2'h1 ? _GEN_3269 : _GEN_9045; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9687 = unuse_way == 2'h1 ? _GEN_3270 : _GEN_9046; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9688 = unuse_way == 2'h1 ? _GEN_3271 : _GEN_9047; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9689 = unuse_way == 2'h1 ? _GEN_3272 : _GEN_9048; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9690 = unuse_way == 2'h1 ? _GEN_3273 : _GEN_9049; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9691 = unuse_way == 2'h1 ? _GEN_3274 : _GEN_9050; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9692 = unuse_way == 2'h1 ? _GEN_3275 : _GEN_9051; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9693 = unuse_way == 2'h1 ? _GEN_3276 : _GEN_9052; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9694 = unuse_way == 2'h1 ? _GEN_3277 : _GEN_9053; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9695 = unuse_way == 2'h1 ? _GEN_3278 : _GEN_9054; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9696 = unuse_way == 2'h1 ? _GEN_3279 : _GEN_9055; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9697 = unuse_way == 2'h1 ? _GEN_3280 : _GEN_9056; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9698 = unuse_way == 2'h1 ? _GEN_3281 : _GEN_9057; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9699 = unuse_way == 2'h1 ? _GEN_3282 : _GEN_9058; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9700 = unuse_way == 2'h1 ? _GEN_3283 : _GEN_9059; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9701 = unuse_way == 2'h1 ? _GEN_3284 : _GEN_9060; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9702 = unuse_way == 2'h1 ? _GEN_3285 : _GEN_9061; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9703 = unuse_way == 2'h1 ? _GEN_3286 : _GEN_9062; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9704 = unuse_way == 2'h1 ? _GEN_3287 : _GEN_9063; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9705 = unuse_way == 2'h1 ? _GEN_3288 : _GEN_9064; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9706 = unuse_way == 2'h1 ? _GEN_3289 : _GEN_9065; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9707 = unuse_way == 2'h1 ? _GEN_3290 : _GEN_9066; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9708 = unuse_way == 2'h1 ? _GEN_3291 : _GEN_9067; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9709 = unuse_way == 2'h1 ? _GEN_3292 : _GEN_9068; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9710 = unuse_way == 2'h1 ? _GEN_3293 : _GEN_9069; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9711 = unuse_way == 2'h1 ? _GEN_3294 : _GEN_9070; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9712 = unuse_way == 2'h1 ? _GEN_3295 : _GEN_9071; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9713 = unuse_way == 2'h1 ? _GEN_3296 : _GEN_9072; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9714 = unuse_way == 2'h1 ? _GEN_3297 : _GEN_9073; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9715 = unuse_way == 2'h1 ? _GEN_3298 : _GEN_9074; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9716 = unuse_way == 2'h1 ? _GEN_3299 : _GEN_9075; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9717 = unuse_way == 2'h1 ? _GEN_3300 : _GEN_9076; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9718 = unuse_way == 2'h1 ? _GEN_3301 : _GEN_9077; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9719 = unuse_way == 2'h1 ? _GEN_3302 : _GEN_9078; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9720 = unuse_way == 2'h1 ? _GEN_3303 : _GEN_9079; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9721 = unuse_way == 2'h1 ? _GEN_3304 : _GEN_9080; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9722 = unuse_way == 2'h1 ? _GEN_3305 : _GEN_9081; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9723 = unuse_way == 2'h1 ? _GEN_3306 : _GEN_9082; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9724 = unuse_way == 2'h1 ? _GEN_3307 : _GEN_9083; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9725 = unuse_way == 2'h1 ? _GEN_3308 : _GEN_9084; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9726 = unuse_way == 2'h1 ? _GEN_3309 : _GEN_9085; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9727 = unuse_way == 2'h1 ? _GEN_3310 : _GEN_9086; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9728 = unuse_way == 2'h1 ? _GEN_3311 : _GEN_9087; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9729 = unuse_way == 2'h1 ? _GEN_3312 : _GEN_9088; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9730 = unuse_way == 2'h1 ? _GEN_3313 : _GEN_9089; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9731 = unuse_way == 2'h1 ? _GEN_3314 : _GEN_9090; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9732 = unuse_way == 2'h1 ? _GEN_3315 : _GEN_9091; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9733 = unuse_way == 2'h1 ? _GEN_3316 : _GEN_9092; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9734 = unuse_way == 2'h1 ? _GEN_3317 : _GEN_9093; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9735 = unuse_way == 2'h1 ? _GEN_3318 : _GEN_9094; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9736 = unuse_way == 2'h1 ? _GEN_3319 : _GEN_9095; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9737 = unuse_way == 2'h1 ? _GEN_3320 : _GEN_9096; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9738 = unuse_way == 2'h1 ? _GEN_3321 : _GEN_9097; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9739 = unuse_way == 2'h1 ? _GEN_3322 : _GEN_9098; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9740 = unuse_way == 2'h1 ? _GEN_3323 : _GEN_9099; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9741 = unuse_way == 2'h1 ? _GEN_3324 : _GEN_9100; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9742 = unuse_way == 2'h1 ? _GEN_3325 : _GEN_9101; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9743 = unuse_way == 2'h1 ? _GEN_3326 : _GEN_9102; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9744 = unuse_way == 2'h1 ? _GEN_3327 : _GEN_9103; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9745 = unuse_way == 2'h1 ? _GEN_3328 : _GEN_9104; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9746 = unuse_way == 2'h1 ? _GEN_3329 : _GEN_9105; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9747 = unuse_way == 2'h1 ? _GEN_3330 : _GEN_9106; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9748 = unuse_way == 2'h1 ? _GEN_3331 : _GEN_9107; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9749 = unuse_way == 2'h1 ? _GEN_3332 : _GEN_9108; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9750 = unuse_way == 2'h1 ? _GEN_3333 : _GEN_9109; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9751 = unuse_way == 2'h1 ? _GEN_3334 : _GEN_9110; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9752 = unuse_way == 2'h1 ? _GEN_3335 : _GEN_9111; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9753 = unuse_way == 2'h1 ? _GEN_3336 : _GEN_9112; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9754 = unuse_way == 2'h1 ? _GEN_3337 : _GEN_9113; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9755 = unuse_way == 2'h1 ? _GEN_3338 : _GEN_9114; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9756 = unuse_way == 2'h1 ? _GEN_3339 : _GEN_9115; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9757 = unuse_way == 2'h1 ? _GEN_3340 : _GEN_9116; // @[d_cache.scala 139:34]
  wire [63:0] _GEN_9758 = unuse_way == 2'h1 ? _GEN_3341 : _GEN_9117; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9759 = unuse_way == 2'h1 ? _GEN_3342 : _GEN_9118; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9760 = unuse_way == 2'h1 ? _GEN_3343 : _GEN_9119; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9761 = unuse_way == 2'h1 ? _GEN_3344 : _GEN_9120; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9762 = unuse_way == 2'h1 ? _GEN_3345 : _GEN_9121; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9763 = unuse_way == 2'h1 ? _GEN_3346 : _GEN_9122; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9764 = unuse_way == 2'h1 ? _GEN_3347 : _GEN_9123; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9765 = unuse_way == 2'h1 ? _GEN_3348 : _GEN_9124; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9766 = unuse_way == 2'h1 ? _GEN_3349 : _GEN_9125; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9767 = unuse_way == 2'h1 ? _GEN_3350 : _GEN_9126; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9768 = unuse_way == 2'h1 ? _GEN_3351 : _GEN_9127; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9769 = unuse_way == 2'h1 ? _GEN_3352 : _GEN_9128; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9770 = unuse_way == 2'h1 ? _GEN_3353 : _GEN_9129; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9771 = unuse_way == 2'h1 ? _GEN_3354 : _GEN_9130; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9772 = unuse_way == 2'h1 ? _GEN_3355 : _GEN_9131; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9773 = unuse_way == 2'h1 ? _GEN_3356 : _GEN_9132; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9774 = unuse_way == 2'h1 ? _GEN_3357 : _GEN_9133; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9775 = unuse_way == 2'h1 ? _GEN_3358 : _GEN_9134; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9776 = unuse_way == 2'h1 ? _GEN_3359 : _GEN_9135; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9777 = unuse_way == 2'h1 ? _GEN_3360 : _GEN_9136; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9778 = unuse_way == 2'h1 ? _GEN_3361 : _GEN_9137; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9779 = unuse_way == 2'h1 ? _GEN_3362 : _GEN_9138; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9780 = unuse_way == 2'h1 ? _GEN_3363 : _GEN_9139; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9781 = unuse_way == 2'h1 ? _GEN_3364 : _GEN_9140; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9782 = unuse_way == 2'h1 ? _GEN_3365 : _GEN_9141; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9783 = unuse_way == 2'h1 ? _GEN_3366 : _GEN_9142; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9784 = unuse_way == 2'h1 ? _GEN_3367 : _GEN_9143; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9785 = unuse_way == 2'h1 ? _GEN_3368 : _GEN_9144; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9786 = unuse_way == 2'h1 ? _GEN_3369 : _GEN_9145; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9787 = unuse_way == 2'h1 ? _GEN_3370 : _GEN_9146; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9788 = unuse_way == 2'h1 ? _GEN_3371 : _GEN_9147; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9789 = unuse_way == 2'h1 ? _GEN_3372 : _GEN_9148; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9790 = unuse_way == 2'h1 ? _GEN_3373 : _GEN_9149; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9791 = unuse_way == 2'h1 ? _GEN_3374 : _GEN_9150; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9792 = unuse_way == 2'h1 ? _GEN_3375 : _GEN_9151; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9793 = unuse_way == 2'h1 ? _GEN_3376 : _GEN_9152; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9794 = unuse_way == 2'h1 ? _GEN_3377 : _GEN_9153; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9795 = unuse_way == 2'h1 ? _GEN_3378 : _GEN_9154; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9796 = unuse_way == 2'h1 ? _GEN_3379 : _GEN_9155; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9797 = unuse_way == 2'h1 ? _GEN_3380 : _GEN_9156; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9798 = unuse_way == 2'h1 ? _GEN_3381 : _GEN_9157; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9799 = unuse_way == 2'h1 ? _GEN_3382 : _GEN_9158; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9800 = unuse_way == 2'h1 ? _GEN_3383 : _GEN_9159; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9801 = unuse_way == 2'h1 ? _GEN_3384 : _GEN_9160; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9802 = unuse_way == 2'h1 ? _GEN_3385 : _GEN_9161; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9803 = unuse_way == 2'h1 ? _GEN_3386 : _GEN_9162; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9804 = unuse_way == 2'h1 ? _GEN_3387 : _GEN_9163; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9805 = unuse_way == 2'h1 ? _GEN_3388 : _GEN_9164; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9806 = unuse_way == 2'h1 ? _GEN_3389 : _GEN_9165; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9807 = unuse_way == 2'h1 ? _GEN_3390 : _GEN_9166; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9808 = unuse_way == 2'h1 ? _GEN_3391 : _GEN_9167; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9809 = unuse_way == 2'h1 ? _GEN_3392 : _GEN_9168; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9810 = unuse_way == 2'h1 ? _GEN_3393 : _GEN_9169; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9811 = unuse_way == 2'h1 ? _GEN_3394 : _GEN_9170; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9812 = unuse_way == 2'h1 ? _GEN_3395 : _GEN_9171; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9813 = unuse_way == 2'h1 ? _GEN_3396 : _GEN_9172; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9814 = unuse_way == 2'h1 ? _GEN_3397 : _GEN_9173; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9815 = unuse_way == 2'h1 ? _GEN_3398 : _GEN_9174; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9816 = unuse_way == 2'h1 ? _GEN_3399 : _GEN_9175; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9817 = unuse_way == 2'h1 ? _GEN_3400 : _GEN_9176; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9818 = unuse_way == 2'h1 ? _GEN_3401 : _GEN_9177; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9819 = unuse_way == 2'h1 ? _GEN_3402 : _GEN_9178; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9820 = unuse_way == 2'h1 ? _GEN_3403 : _GEN_9179; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9821 = unuse_way == 2'h1 ? _GEN_3404 : _GEN_9180; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9822 = unuse_way == 2'h1 ? _GEN_3405 : _GEN_9181; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9823 = unuse_way == 2'h1 ? _GEN_3406 : _GEN_9182; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9824 = unuse_way == 2'h1 ? _GEN_3407 : _GEN_9183; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9825 = unuse_way == 2'h1 ? _GEN_3408 : _GEN_9184; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9826 = unuse_way == 2'h1 ? _GEN_3409 : _GEN_9185; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9827 = unuse_way == 2'h1 ? _GEN_3410 : _GEN_9186; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9828 = unuse_way == 2'h1 ? _GEN_3411 : _GEN_9187; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9829 = unuse_way == 2'h1 ? _GEN_3412 : _GEN_9188; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9830 = unuse_way == 2'h1 ? _GEN_3413 : _GEN_9189; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9831 = unuse_way == 2'h1 ? _GEN_3414 : _GEN_9190; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9832 = unuse_way == 2'h1 ? _GEN_3415 : _GEN_9191; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9833 = unuse_way == 2'h1 ? _GEN_3416 : _GEN_9192; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9834 = unuse_way == 2'h1 ? _GEN_3417 : _GEN_9193; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9835 = unuse_way == 2'h1 ? _GEN_3418 : _GEN_9194; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9836 = unuse_way == 2'h1 ? _GEN_3419 : _GEN_9195; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9837 = unuse_way == 2'h1 ? _GEN_3420 : _GEN_9196; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9838 = unuse_way == 2'h1 ? _GEN_3421 : _GEN_9197; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9839 = unuse_way == 2'h1 ? _GEN_3422 : _GEN_9198; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9840 = unuse_way == 2'h1 ? _GEN_3423 : _GEN_9199; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9841 = unuse_way == 2'h1 ? _GEN_3424 : _GEN_9200; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9842 = unuse_way == 2'h1 ? _GEN_3425 : _GEN_9201; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9843 = unuse_way == 2'h1 ? _GEN_3426 : _GEN_9202; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9844 = unuse_way == 2'h1 ? _GEN_3427 : _GEN_9203; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9845 = unuse_way == 2'h1 ? _GEN_3428 : _GEN_9204; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9846 = unuse_way == 2'h1 ? _GEN_3429 : _GEN_9205; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9847 = unuse_way == 2'h1 ? _GEN_3430 : _GEN_9206; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9848 = unuse_way == 2'h1 ? _GEN_3431 : _GEN_9207; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9849 = unuse_way == 2'h1 ? _GEN_3432 : _GEN_9208; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9850 = unuse_way == 2'h1 ? _GEN_3433 : _GEN_9209; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9851 = unuse_way == 2'h1 ? _GEN_3434 : _GEN_9210; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9852 = unuse_way == 2'h1 ? _GEN_3435 : _GEN_9211; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9853 = unuse_way == 2'h1 ? _GEN_3436 : _GEN_9212; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9854 = unuse_way == 2'h1 ? _GEN_3437 : _GEN_9213; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9855 = unuse_way == 2'h1 ? _GEN_3438 : _GEN_9214; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9856 = unuse_way == 2'h1 ? _GEN_3439 : _GEN_9215; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9857 = unuse_way == 2'h1 ? _GEN_3440 : _GEN_9216; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9858 = unuse_way == 2'h1 ? _GEN_3441 : _GEN_9217; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9859 = unuse_way == 2'h1 ? _GEN_3442 : _GEN_9218; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9860 = unuse_way == 2'h1 ? _GEN_3443 : _GEN_9219; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9861 = unuse_way == 2'h1 ? _GEN_3444 : _GEN_9220; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9862 = unuse_way == 2'h1 ? _GEN_3445 : _GEN_9221; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9863 = unuse_way == 2'h1 ? _GEN_3446 : _GEN_9222; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9864 = unuse_way == 2'h1 ? _GEN_3447 : _GEN_9223; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9865 = unuse_way == 2'h1 ? _GEN_3448 : _GEN_9224; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9866 = unuse_way == 2'h1 ? _GEN_3449 : _GEN_9225; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9867 = unuse_way == 2'h1 ? _GEN_3450 : _GEN_9226; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9868 = unuse_way == 2'h1 ? _GEN_3451 : _GEN_9227; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9869 = unuse_way == 2'h1 ? _GEN_3452 : _GEN_9228; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9870 = unuse_way == 2'h1 ? _GEN_3453 : _GEN_9229; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9871 = unuse_way == 2'h1 ? _GEN_3454 : _GEN_9230; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9872 = unuse_way == 2'h1 ? _GEN_3455 : _GEN_9231; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9873 = unuse_way == 2'h1 ? _GEN_3456 : _GEN_9232; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9874 = unuse_way == 2'h1 ? _GEN_3457 : _GEN_9233; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9875 = unuse_way == 2'h1 ? _GEN_3458 : _GEN_9234; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9876 = unuse_way == 2'h1 ? _GEN_3459 : _GEN_9235; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9877 = unuse_way == 2'h1 ? _GEN_3460 : _GEN_9236; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9878 = unuse_way == 2'h1 ? _GEN_3461 : _GEN_9237; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9879 = unuse_way == 2'h1 ? _GEN_3462 : _GEN_9238; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9880 = unuse_way == 2'h1 ? _GEN_3463 : _GEN_9239; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9881 = unuse_way == 2'h1 ? _GEN_3464 : _GEN_9240; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9882 = unuse_way == 2'h1 ? _GEN_3465 : _GEN_9241; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9883 = unuse_way == 2'h1 ? _GEN_3466 : _GEN_9242; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9884 = unuse_way == 2'h1 ? _GEN_3467 : _GEN_9243; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9885 = unuse_way == 2'h1 ? _GEN_3468 : _GEN_9244; // @[d_cache.scala 139:34]
  wire [31:0] _GEN_9886 = unuse_way == 2'h1 ? _GEN_3469 : _GEN_9245; // @[d_cache.scala 139:34]
  wire  _GEN_9887 = unuse_way == 2'h1 ? _GEN_3470 : _GEN_9374; // @[d_cache.scala 139:34]
  wire  _GEN_9888 = unuse_way == 2'h1 ? _GEN_3471 : _GEN_9375; // @[d_cache.scala 139:34]
  wire  _GEN_9889 = unuse_way == 2'h1 ? _GEN_3472 : _GEN_9376; // @[d_cache.scala 139:34]
  wire  _GEN_9890 = unuse_way == 2'h1 ? _GEN_3473 : _GEN_9377; // @[d_cache.scala 139:34]
  wire  _GEN_9891 = unuse_way == 2'h1 ? _GEN_3474 : _GEN_9378; // @[d_cache.scala 139:34]
  wire  _GEN_9892 = unuse_way == 2'h1 ? _GEN_3475 : _GEN_9379; // @[d_cache.scala 139:34]
  wire  _GEN_9893 = unuse_way == 2'h1 ? _GEN_3476 : _GEN_9380; // @[d_cache.scala 139:34]
  wire  _GEN_9894 = unuse_way == 2'h1 ? _GEN_3477 : _GEN_9381; // @[d_cache.scala 139:34]
  wire  _GEN_9895 = unuse_way == 2'h1 ? _GEN_3478 : _GEN_9382; // @[d_cache.scala 139:34]
  wire  _GEN_9896 = unuse_way == 2'h1 ? _GEN_3479 : _GEN_9383; // @[d_cache.scala 139:34]
  wire  _GEN_9897 = unuse_way == 2'h1 ? _GEN_3480 : _GEN_9384; // @[d_cache.scala 139:34]
  wire  _GEN_9898 = unuse_way == 2'h1 ? _GEN_3481 : _GEN_9385; // @[d_cache.scala 139:34]
  wire  _GEN_9899 = unuse_way == 2'h1 ? _GEN_3482 : _GEN_9386; // @[d_cache.scala 139:34]
  wire  _GEN_9900 = unuse_way == 2'h1 ? _GEN_3483 : _GEN_9387; // @[d_cache.scala 139:34]
  wire  _GEN_9901 = unuse_way == 2'h1 ? _GEN_3484 : _GEN_9388; // @[d_cache.scala 139:34]
  wire  _GEN_9902 = unuse_way == 2'h1 ? _GEN_3485 : _GEN_9389; // @[d_cache.scala 139:34]
  wire  _GEN_9903 = unuse_way == 2'h1 ? _GEN_3486 : _GEN_9390; // @[d_cache.scala 139:34]
  wire  _GEN_9904 = unuse_way == 2'h1 ? _GEN_3487 : _GEN_9391; // @[d_cache.scala 139:34]
  wire  _GEN_9905 = unuse_way == 2'h1 ? _GEN_3488 : _GEN_9392; // @[d_cache.scala 139:34]
  wire  _GEN_9906 = unuse_way == 2'h1 ? _GEN_3489 : _GEN_9393; // @[d_cache.scala 139:34]
  wire  _GEN_9907 = unuse_way == 2'h1 ? _GEN_3490 : _GEN_9394; // @[d_cache.scala 139:34]
  wire  _GEN_9908 = unuse_way == 2'h1 ? _GEN_3491 : _GEN_9395; // @[d_cache.scala 139:34]
  wire  _GEN_9909 = unuse_way == 2'h1 ? _GEN_3492 : _GEN_9396; // @[d_cache.scala 139:34]
  wire  _GEN_9910 = unuse_way == 2'h1 ? _GEN_3493 : _GEN_9397; // @[d_cache.scala 139:34]
  wire  _GEN_9911 = unuse_way == 2'h1 ? _GEN_3494 : _GEN_9398; // @[d_cache.scala 139:34]
  wire  _GEN_9912 = unuse_way == 2'h1 ? _GEN_3495 : _GEN_9399; // @[d_cache.scala 139:34]
  wire  _GEN_9913 = unuse_way == 2'h1 ? _GEN_3496 : _GEN_9400; // @[d_cache.scala 139:34]
  wire  _GEN_9914 = unuse_way == 2'h1 ? _GEN_3497 : _GEN_9401; // @[d_cache.scala 139:34]
  wire  _GEN_9915 = unuse_way == 2'h1 ? _GEN_3498 : _GEN_9402; // @[d_cache.scala 139:34]
  wire  _GEN_9916 = unuse_way == 2'h1 ? _GEN_3499 : _GEN_9403; // @[d_cache.scala 139:34]
  wire  _GEN_9917 = unuse_way == 2'h1 ? _GEN_3500 : _GEN_9404; // @[d_cache.scala 139:34]
  wire  _GEN_9918 = unuse_way == 2'h1 ? _GEN_3501 : _GEN_9405; // @[d_cache.scala 139:34]
  wire  _GEN_9919 = unuse_way == 2'h1 ? _GEN_3502 : _GEN_9406; // @[d_cache.scala 139:34]
  wire  _GEN_9920 = unuse_way == 2'h1 ? _GEN_3503 : _GEN_9407; // @[d_cache.scala 139:34]
  wire  _GEN_9921 = unuse_way == 2'h1 ? _GEN_3504 : _GEN_9408; // @[d_cache.scala 139:34]
  wire  _GEN_9922 = unuse_way == 2'h1 ? _GEN_3505 : _GEN_9409; // @[d_cache.scala 139:34]
  wire  _GEN_9923 = unuse_way == 2'h1 ? _GEN_3506 : _GEN_9410; // @[d_cache.scala 139:34]
  wire  _GEN_9924 = unuse_way == 2'h1 ? _GEN_3507 : _GEN_9411; // @[d_cache.scala 139:34]
  wire  _GEN_9925 = unuse_way == 2'h1 ? _GEN_3508 : _GEN_9412; // @[d_cache.scala 139:34]
  wire  _GEN_9926 = unuse_way == 2'h1 ? _GEN_3509 : _GEN_9413; // @[d_cache.scala 139:34]
  wire  _GEN_9927 = unuse_way == 2'h1 ? _GEN_3510 : _GEN_9414; // @[d_cache.scala 139:34]
  wire  _GEN_9928 = unuse_way == 2'h1 ? _GEN_3511 : _GEN_9415; // @[d_cache.scala 139:34]
  wire  _GEN_9929 = unuse_way == 2'h1 ? _GEN_3512 : _GEN_9416; // @[d_cache.scala 139:34]
  wire  _GEN_9930 = unuse_way == 2'h1 ? _GEN_3513 : _GEN_9417; // @[d_cache.scala 139:34]
  wire  _GEN_9931 = unuse_way == 2'h1 ? _GEN_3514 : _GEN_9418; // @[d_cache.scala 139:34]
  wire  _GEN_9932 = unuse_way == 2'h1 ? _GEN_3515 : _GEN_9419; // @[d_cache.scala 139:34]
  wire  _GEN_9933 = unuse_way == 2'h1 ? _GEN_3516 : _GEN_9420; // @[d_cache.scala 139:34]
  wire  _GEN_9934 = unuse_way == 2'h1 ? _GEN_3517 : _GEN_9421; // @[d_cache.scala 139:34]
  wire  _GEN_9935 = unuse_way == 2'h1 ? _GEN_3518 : _GEN_9422; // @[d_cache.scala 139:34]
  wire  _GEN_9936 = unuse_way == 2'h1 ? _GEN_3519 : _GEN_9423; // @[d_cache.scala 139:34]
  wire  _GEN_9937 = unuse_way == 2'h1 ? _GEN_3520 : _GEN_9424; // @[d_cache.scala 139:34]
  wire  _GEN_9938 = unuse_way == 2'h1 ? _GEN_3521 : _GEN_9425; // @[d_cache.scala 139:34]
  wire  _GEN_9939 = unuse_way == 2'h1 ? _GEN_3522 : _GEN_9426; // @[d_cache.scala 139:34]
  wire  _GEN_9940 = unuse_way == 2'h1 ? _GEN_3523 : _GEN_9427; // @[d_cache.scala 139:34]
  wire  _GEN_9941 = unuse_way == 2'h1 ? _GEN_3524 : _GEN_9428; // @[d_cache.scala 139:34]
  wire  _GEN_9942 = unuse_way == 2'h1 ? _GEN_3525 : _GEN_9429; // @[d_cache.scala 139:34]
  wire  _GEN_9943 = unuse_way == 2'h1 ? _GEN_3526 : _GEN_9430; // @[d_cache.scala 139:34]
  wire  _GEN_9944 = unuse_way == 2'h1 ? _GEN_3527 : _GEN_9431; // @[d_cache.scala 139:34]
  wire  _GEN_9945 = unuse_way == 2'h1 ? _GEN_3528 : _GEN_9432; // @[d_cache.scala 139:34]
  wire  _GEN_9946 = unuse_way == 2'h1 ? _GEN_3529 : _GEN_9433; // @[d_cache.scala 139:34]
  wire  _GEN_9947 = unuse_way == 2'h1 ? _GEN_3530 : _GEN_9434; // @[d_cache.scala 139:34]
  wire  _GEN_9948 = unuse_way == 2'h1 ? _GEN_3531 : _GEN_9435; // @[d_cache.scala 139:34]
  wire  _GEN_9949 = unuse_way == 2'h1 ? _GEN_3532 : _GEN_9436; // @[d_cache.scala 139:34]
  wire  _GEN_9950 = unuse_way == 2'h1 ? _GEN_3533 : _GEN_9437; // @[d_cache.scala 139:34]
  wire  _GEN_9951 = unuse_way == 2'h1 ? _GEN_3534 : _GEN_9438; // @[d_cache.scala 139:34]
  wire  _GEN_9952 = unuse_way == 2'h1 ? _GEN_3535 : _GEN_9439; // @[d_cache.scala 139:34]
  wire  _GEN_9953 = unuse_way == 2'h1 ? _GEN_3536 : _GEN_9440; // @[d_cache.scala 139:34]
  wire  _GEN_9954 = unuse_way == 2'h1 ? _GEN_3537 : _GEN_9441; // @[d_cache.scala 139:34]
  wire  _GEN_9955 = unuse_way == 2'h1 ? _GEN_3538 : _GEN_9442; // @[d_cache.scala 139:34]
  wire  _GEN_9956 = unuse_way == 2'h1 ? _GEN_3539 : _GEN_9443; // @[d_cache.scala 139:34]
  wire  _GEN_9957 = unuse_way == 2'h1 ? _GEN_3540 : _GEN_9444; // @[d_cache.scala 139:34]
  wire  _GEN_9958 = unuse_way == 2'h1 ? _GEN_3541 : _GEN_9445; // @[d_cache.scala 139:34]
  wire  _GEN_9959 = unuse_way == 2'h1 ? _GEN_3542 : _GEN_9446; // @[d_cache.scala 139:34]
  wire  _GEN_9960 = unuse_way == 2'h1 ? _GEN_3543 : _GEN_9447; // @[d_cache.scala 139:34]
  wire  _GEN_9961 = unuse_way == 2'h1 ? _GEN_3544 : _GEN_9448; // @[d_cache.scala 139:34]
  wire  _GEN_9962 = unuse_way == 2'h1 ? _GEN_3545 : _GEN_9449; // @[d_cache.scala 139:34]
  wire  _GEN_9963 = unuse_way == 2'h1 ? _GEN_3546 : _GEN_9450; // @[d_cache.scala 139:34]
  wire  _GEN_9964 = unuse_way == 2'h1 ? _GEN_3547 : _GEN_9451; // @[d_cache.scala 139:34]
  wire  _GEN_9965 = unuse_way == 2'h1 ? _GEN_3548 : _GEN_9452; // @[d_cache.scala 139:34]
  wire  _GEN_9966 = unuse_way == 2'h1 ? _GEN_3549 : _GEN_9453; // @[d_cache.scala 139:34]
  wire  _GEN_9967 = unuse_way == 2'h1 ? _GEN_3550 : _GEN_9454; // @[d_cache.scala 139:34]
  wire  _GEN_9968 = unuse_way == 2'h1 ? _GEN_3551 : _GEN_9455; // @[d_cache.scala 139:34]
  wire  _GEN_9969 = unuse_way == 2'h1 ? _GEN_3552 : _GEN_9456; // @[d_cache.scala 139:34]
  wire  _GEN_9970 = unuse_way == 2'h1 ? _GEN_3553 : _GEN_9457; // @[d_cache.scala 139:34]
  wire  _GEN_9971 = unuse_way == 2'h1 ? _GEN_3554 : _GEN_9458; // @[d_cache.scala 139:34]
  wire  _GEN_9972 = unuse_way == 2'h1 ? _GEN_3555 : _GEN_9459; // @[d_cache.scala 139:34]
  wire  _GEN_9973 = unuse_way == 2'h1 ? _GEN_3556 : _GEN_9460; // @[d_cache.scala 139:34]
  wire  _GEN_9974 = unuse_way == 2'h1 ? _GEN_3557 : _GEN_9461; // @[d_cache.scala 139:34]
  wire  _GEN_9975 = unuse_way == 2'h1 ? _GEN_3558 : _GEN_9462; // @[d_cache.scala 139:34]
  wire  _GEN_9976 = unuse_way == 2'h1 ? _GEN_3559 : _GEN_9463; // @[d_cache.scala 139:34]
  wire  _GEN_9977 = unuse_way == 2'h1 ? _GEN_3560 : _GEN_9464; // @[d_cache.scala 139:34]
  wire  _GEN_9978 = unuse_way == 2'h1 ? _GEN_3561 : _GEN_9465; // @[d_cache.scala 139:34]
  wire  _GEN_9979 = unuse_way == 2'h1 ? _GEN_3562 : _GEN_9466; // @[d_cache.scala 139:34]
  wire  _GEN_9980 = unuse_way == 2'h1 ? _GEN_3563 : _GEN_9467; // @[d_cache.scala 139:34]
  wire  _GEN_9981 = unuse_way == 2'h1 ? _GEN_3564 : _GEN_9468; // @[d_cache.scala 139:34]
  wire  _GEN_9982 = unuse_way == 2'h1 ? _GEN_3565 : _GEN_9469; // @[d_cache.scala 139:34]
  wire  _GEN_9983 = unuse_way == 2'h1 ? _GEN_3566 : _GEN_9470; // @[d_cache.scala 139:34]
  wire  _GEN_9984 = unuse_way == 2'h1 ? _GEN_3567 : _GEN_9471; // @[d_cache.scala 139:34]
  wire  _GEN_9985 = unuse_way == 2'h1 ? _GEN_3568 : _GEN_9472; // @[d_cache.scala 139:34]
  wire  _GEN_9986 = unuse_way == 2'h1 ? _GEN_3569 : _GEN_9473; // @[d_cache.scala 139:34]
  wire  _GEN_9987 = unuse_way == 2'h1 ? _GEN_3570 : _GEN_9474; // @[d_cache.scala 139:34]
  wire  _GEN_9988 = unuse_way == 2'h1 ? _GEN_3571 : _GEN_9475; // @[d_cache.scala 139:34]
  wire  _GEN_9989 = unuse_way == 2'h1 ? _GEN_3572 : _GEN_9476; // @[d_cache.scala 139:34]
  wire  _GEN_9990 = unuse_way == 2'h1 ? _GEN_3573 : _GEN_9477; // @[d_cache.scala 139:34]
  wire  _GEN_9991 = unuse_way == 2'h1 ? _GEN_3574 : _GEN_9478; // @[d_cache.scala 139:34]
  wire  _GEN_9992 = unuse_way == 2'h1 ? _GEN_3575 : _GEN_9479; // @[d_cache.scala 139:34]
  wire  _GEN_9993 = unuse_way == 2'h1 ? _GEN_3576 : _GEN_9480; // @[d_cache.scala 139:34]
  wire  _GEN_9994 = unuse_way == 2'h1 ? _GEN_3577 : _GEN_9481; // @[d_cache.scala 139:34]
  wire  _GEN_9995 = unuse_way == 2'h1 ? _GEN_3578 : _GEN_9482; // @[d_cache.scala 139:34]
  wire  _GEN_9996 = unuse_way == 2'h1 ? _GEN_3579 : _GEN_9483; // @[d_cache.scala 139:34]
  wire  _GEN_9997 = unuse_way == 2'h1 ? _GEN_3580 : _GEN_9484; // @[d_cache.scala 139:34]
  wire  _GEN_9998 = unuse_way == 2'h1 ? _GEN_3581 : _GEN_9485; // @[d_cache.scala 139:34]
  wire  _GEN_9999 = unuse_way == 2'h1 ? _GEN_3582 : _GEN_9486; // @[d_cache.scala 139:34]
  wire  _GEN_10000 = unuse_way == 2'h1 ? _GEN_3583 : _GEN_9487; // @[d_cache.scala 139:34]
  wire  _GEN_10001 = unuse_way == 2'h1 ? _GEN_3584 : _GEN_9488; // @[d_cache.scala 139:34]
  wire  _GEN_10002 = unuse_way == 2'h1 ? _GEN_3585 : _GEN_9489; // @[d_cache.scala 139:34]
  wire  _GEN_10003 = unuse_way == 2'h1 ? _GEN_3586 : _GEN_9490; // @[d_cache.scala 139:34]
  wire  _GEN_10004 = unuse_way == 2'h1 ? _GEN_3587 : _GEN_9491; // @[d_cache.scala 139:34]
  wire  _GEN_10005 = unuse_way == 2'h1 ? _GEN_3588 : _GEN_9492; // @[d_cache.scala 139:34]
  wire  _GEN_10006 = unuse_way == 2'h1 ? _GEN_3589 : _GEN_9493; // @[d_cache.scala 139:34]
  wire  _GEN_10007 = unuse_way == 2'h1 ? _GEN_3590 : _GEN_9494; // @[d_cache.scala 139:34]
  wire  _GEN_10008 = unuse_way == 2'h1 ? _GEN_3591 : _GEN_9495; // @[d_cache.scala 139:34]
  wire  _GEN_10009 = unuse_way == 2'h1 ? _GEN_3592 : _GEN_9496; // @[d_cache.scala 139:34]
  wire  _GEN_10010 = unuse_way == 2'h1 ? _GEN_3593 : _GEN_9497; // @[d_cache.scala 139:34]
  wire  _GEN_10011 = unuse_way == 2'h1 ? _GEN_3594 : _GEN_9498; // @[d_cache.scala 139:34]
  wire  _GEN_10012 = unuse_way == 2'h1 ? _GEN_3595 : _GEN_9499; // @[d_cache.scala 139:34]
  wire  _GEN_10013 = unuse_way == 2'h1 ? _GEN_3596 : _GEN_9500; // @[d_cache.scala 139:34]
  wire  _GEN_10014 = unuse_way == 2'h1 ? _GEN_3597 : _GEN_9501; // @[d_cache.scala 139:34]
  wire  _GEN_10015 = unuse_way == 2'h1 | _GEN_8987; // @[d_cache.scala 139:34 144:23]
  wire [63:0] _GEN_10016 = unuse_way == 2'h1 ? ram_1_0 : _GEN_8603; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10017 = unuse_way == 2'h1 ? ram_1_1 : _GEN_8604; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10018 = unuse_way == 2'h1 ? ram_1_2 : _GEN_8605; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10019 = unuse_way == 2'h1 ? ram_1_3 : _GEN_8606; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10020 = unuse_way == 2'h1 ? ram_1_4 : _GEN_8607; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10021 = unuse_way == 2'h1 ? ram_1_5 : _GEN_8608; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10022 = unuse_way == 2'h1 ? ram_1_6 : _GEN_8609; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10023 = unuse_way == 2'h1 ? ram_1_7 : _GEN_8610; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10024 = unuse_way == 2'h1 ? ram_1_8 : _GEN_8611; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10025 = unuse_way == 2'h1 ? ram_1_9 : _GEN_8612; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10026 = unuse_way == 2'h1 ? ram_1_10 : _GEN_8613; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10027 = unuse_way == 2'h1 ? ram_1_11 : _GEN_8614; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10028 = unuse_way == 2'h1 ? ram_1_12 : _GEN_8615; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10029 = unuse_way == 2'h1 ? ram_1_13 : _GEN_8616; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10030 = unuse_way == 2'h1 ? ram_1_14 : _GEN_8617; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10031 = unuse_way == 2'h1 ? ram_1_15 : _GEN_8618; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10032 = unuse_way == 2'h1 ? ram_1_16 : _GEN_8619; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10033 = unuse_way == 2'h1 ? ram_1_17 : _GEN_8620; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10034 = unuse_way == 2'h1 ? ram_1_18 : _GEN_8621; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10035 = unuse_way == 2'h1 ? ram_1_19 : _GEN_8622; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10036 = unuse_way == 2'h1 ? ram_1_20 : _GEN_8623; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10037 = unuse_way == 2'h1 ? ram_1_21 : _GEN_8624; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10038 = unuse_way == 2'h1 ? ram_1_22 : _GEN_8625; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10039 = unuse_way == 2'h1 ? ram_1_23 : _GEN_8626; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10040 = unuse_way == 2'h1 ? ram_1_24 : _GEN_8627; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10041 = unuse_way == 2'h1 ? ram_1_25 : _GEN_8628; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10042 = unuse_way == 2'h1 ? ram_1_26 : _GEN_8629; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10043 = unuse_way == 2'h1 ? ram_1_27 : _GEN_8630; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10044 = unuse_way == 2'h1 ? ram_1_28 : _GEN_8631; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10045 = unuse_way == 2'h1 ? ram_1_29 : _GEN_8632; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10046 = unuse_way == 2'h1 ? ram_1_30 : _GEN_8633; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10047 = unuse_way == 2'h1 ? ram_1_31 : _GEN_8634; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10048 = unuse_way == 2'h1 ? ram_1_32 : _GEN_8635; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10049 = unuse_way == 2'h1 ? ram_1_33 : _GEN_8636; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10050 = unuse_way == 2'h1 ? ram_1_34 : _GEN_8637; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10051 = unuse_way == 2'h1 ? ram_1_35 : _GEN_8638; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10052 = unuse_way == 2'h1 ? ram_1_36 : _GEN_8639; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10053 = unuse_way == 2'h1 ? ram_1_37 : _GEN_8640; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10054 = unuse_way == 2'h1 ? ram_1_38 : _GEN_8641; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10055 = unuse_way == 2'h1 ? ram_1_39 : _GEN_8642; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10056 = unuse_way == 2'h1 ? ram_1_40 : _GEN_8643; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10057 = unuse_way == 2'h1 ? ram_1_41 : _GEN_8644; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10058 = unuse_way == 2'h1 ? ram_1_42 : _GEN_8645; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10059 = unuse_way == 2'h1 ? ram_1_43 : _GEN_8646; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10060 = unuse_way == 2'h1 ? ram_1_44 : _GEN_8647; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10061 = unuse_way == 2'h1 ? ram_1_45 : _GEN_8648; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10062 = unuse_way == 2'h1 ? ram_1_46 : _GEN_8649; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10063 = unuse_way == 2'h1 ? ram_1_47 : _GEN_8650; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10064 = unuse_way == 2'h1 ? ram_1_48 : _GEN_8651; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10065 = unuse_way == 2'h1 ? ram_1_49 : _GEN_8652; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10066 = unuse_way == 2'h1 ? ram_1_50 : _GEN_8653; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10067 = unuse_way == 2'h1 ? ram_1_51 : _GEN_8654; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10068 = unuse_way == 2'h1 ? ram_1_52 : _GEN_8655; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10069 = unuse_way == 2'h1 ? ram_1_53 : _GEN_8656; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10070 = unuse_way == 2'h1 ? ram_1_54 : _GEN_8657; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10071 = unuse_way == 2'h1 ? ram_1_55 : _GEN_8658; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10072 = unuse_way == 2'h1 ? ram_1_56 : _GEN_8659; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10073 = unuse_way == 2'h1 ? ram_1_57 : _GEN_8660; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10074 = unuse_way == 2'h1 ? ram_1_58 : _GEN_8661; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10075 = unuse_way == 2'h1 ? ram_1_59 : _GEN_8662; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10076 = unuse_way == 2'h1 ? ram_1_60 : _GEN_8663; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10077 = unuse_way == 2'h1 ? ram_1_61 : _GEN_8664; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10078 = unuse_way == 2'h1 ? ram_1_62 : _GEN_8665; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10079 = unuse_way == 2'h1 ? ram_1_63 : _GEN_8666; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10080 = unuse_way == 2'h1 ? ram_1_64 : _GEN_8667; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10081 = unuse_way == 2'h1 ? ram_1_65 : _GEN_8668; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10082 = unuse_way == 2'h1 ? ram_1_66 : _GEN_8669; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10083 = unuse_way == 2'h1 ? ram_1_67 : _GEN_8670; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10084 = unuse_way == 2'h1 ? ram_1_68 : _GEN_8671; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10085 = unuse_way == 2'h1 ? ram_1_69 : _GEN_8672; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10086 = unuse_way == 2'h1 ? ram_1_70 : _GEN_8673; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10087 = unuse_way == 2'h1 ? ram_1_71 : _GEN_8674; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10088 = unuse_way == 2'h1 ? ram_1_72 : _GEN_8675; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10089 = unuse_way == 2'h1 ? ram_1_73 : _GEN_8676; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10090 = unuse_way == 2'h1 ? ram_1_74 : _GEN_8677; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10091 = unuse_way == 2'h1 ? ram_1_75 : _GEN_8678; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10092 = unuse_way == 2'h1 ? ram_1_76 : _GEN_8679; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10093 = unuse_way == 2'h1 ? ram_1_77 : _GEN_8680; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10094 = unuse_way == 2'h1 ? ram_1_78 : _GEN_8681; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10095 = unuse_way == 2'h1 ? ram_1_79 : _GEN_8682; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10096 = unuse_way == 2'h1 ? ram_1_80 : _GEN_8683; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10097 = unuse_way == 2'h1 ? ram_1_81 : _GEN_8684; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10098 = unuse_way == 2'h1 ? ram_1_82 : _GEN_8685; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10099 = unuse_way == 2'h1 ? ram_1_83 : _GEN_8686; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10100 = unuse_way == 2'h1 ? ram_1_84 : _GEN_8687; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10101 = unuse_way == 2'h1 ? ram_1_85 : _GEN_8688; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10102 = unuse_way == 2'h1 ? ram_1_86 : _GEN_8689; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10103 = unuse_way == 2'h1 ? ram_1_87 : _GEN_8690; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10104 = unuse_way == 2'h1 ? ram_1_88 : _GEN_8691; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10105 = unuse_way == 2'h1 ? ram_1_89 : _GEN_8692; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10106 = unuse_way == 2'h1 ? ram_1_90 : _GEN_8693; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10107 = unuse_way == 2'h1 ? ram_1_91 : _GEN_8694; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10108 = unuse_way == 2'h1 ? ram_1_92 : _GEN_8695; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10109 = unuse_way == 2'h1 ? ram_1_93 : _GEN_8696; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10110 = unuse_way == 2'h1 ? ram_1_94 : _GEN_8697; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10111 = unuse_way == 2'h1 ? ram_1_95 : _GEN_8698; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10112 = unuse_way == 2'h1 ? ram_1_96 : _GEN_8699; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10113 = unuse_way == 2'h1 ? ram_1_97 : _GEN_8700; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10114 = unuse_way == 2'h1 ? ram_1_98 : _GEN_8701; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10115 = unuse_way == 2'h1 ? ram_1_99 : _GEN_8702; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10116 = unuse_way == 2'h1 ? ram_1_100 : _GEN_8703; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10117 = unuse_way == 2'h1 ? ram_1_101 : _GEN_8704; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10118 = unuse_way == 2'h1 ? ram_1_102 : _GEN_8705; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10119 = unuse_way == 2'h1 ? ram_1_103 : _GEN_8706; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10120 = unuse_way == 2'h1 ? ram_1_104 : _GEN_8707; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10121 = unuse_way == 2'h1 ? ram_1_105 : _GEN_8708; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10122 = unuse_way == 2'h1 ? ram_1_106 : _GEN_8709; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10123 = unuse_way == 2'h1 ? ram_1_107 : _GEN_8710; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10124 = unuse_way == 2'h1 ? ram_1_108 : _GEN_8711; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10125 = unuse_way == 2'h1 ? ram_1_109 : _GEN_8712; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10126 = unuse_way == 2'h1 ? ram_1_110 : _GEN_8713; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10127 = unuse_way == 2'h1 ? ram_1_111 : _GEN_8714; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10128 = unuse_way == 2'h1 ? ram_1_112 : _GEN_8715; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10129 = unuse_way == 2'h1 ? ram_1_113 : _GEN_8716; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10130 = unuse_way == 2'h1 ? ram_1_114 : _GEN_8717; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10131 = unuse_way == 2'h1 ? ram_1_115 : _GEN_8718; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10132 = unuse_way == 2'h1 ? ram_1_116 : _GEN_8719; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10133 = unuse_way == 2'h1 ? ram_1_117 : _GEN_8720; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10134 = unuse_way == 2'h1 ? ram_1_118 : _GEN_8721; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10135 = unuse_way == 2'h1 ? ram_1_119 : _GEN_8722; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10136 = unuse_way == 2'h1 ? ram_1_120 : _GEN_8723; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10137 = unuse_way == 2'h1 ? ram_1_121 : _GEN_8724; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10138 = unuse_way == 2'h1 ? ram_1_122 : _GEN_8725; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10139 = unuse_way == 2'h1 ? ram_1_123 : _GEN_8726; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10140 = unuse_way == 2'h1 ? ram_1_124 : _GEN_8727; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10141 = unuse_way == 2'h1 ? ram_1_125 : _GEN_8728; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10142 = unuse_way == 2'h1 ? ram_1_126 : _GEN_8729; // @[d_cache.scala 139:34 19:24]
  wire [63:0] _GEN_10143 = unuse_way == 2'h1 ? ram_1_127 : _GEN_8730; // @[d_cache.scala 139:34 19:24]
  wire [31:0] _GEN_10144 = unuse_way == 2'h1 ? tag_1_0 : _GEN_8731; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10145 = unuse_way == 2'h1 ? tag_1_1 : _GEN_8732; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10146 = unuse_way == 2'h1 ? tag_1_2 : _GEN_8733; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10147 = unuse_way == 2'h1 ? tag_1_3 : _GEN_8734; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10148 = unuse_way == 2'h1 ? tag_1_4 : _GEN_8735; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10149 = unuse_way == 2'h1 ? tag_1_5 : _GEN_8736; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10150 = unuse_way == 2'h1 ? tag_1_6 : _GEN_8737; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10151 = unuse_way == 2'h1 ? tag_1_7 : _GEN_8738; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10152 = unuse_way == 2'h1 ? tag_1_8 : _GEN_8739; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10153 = unuse_way == 2'h1 ? tag_1_9 : _GEN_8740; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10154 = unuse_way == 2'h1 ? tag_1_10 : _GEN_8741; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10155 = unuse_way == 2'h1 ? tag_1_11 : _GEN_8742; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10156 = unuse_way == 2'h1 ? tag_1_12 : _GEN_8743; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10157 = unuse_way == 2'h1 ? tag_1_13 : _GEN_8744; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10158 = unuse_way == 2'h1 ? tag_1_14 : _GEN_8745; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10159 = unuse_way == 2'h1 ? tag_1_15 : _GEN_8746; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10160 = unuse_way == 2'h1 ? tag_1_16 : _GEN_8747; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10161 = unuse_way == 2'h1 ? tag_1_17 : _GEN_8748; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10162 = unuse_way == 2'h1 ? tag_1_18 : _GEN_8749; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10163 = unuse_way == 2'h1 ? tag_1_19 : _GEN_8750; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10164 = unuse_way == 2'h1 ? tag_1_20 : _GEN_8751; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10165 = unuse_way == 2'h1 ? tag_1_21 : _GEN_8752; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10166 = unuse_way == 2'h1 ? tag_1_22 : _GEN_8753; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10167 = unuse_way == 2'h1 ? tag_1_23 : _GEN_8754; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10168 = unuse_way == 2'h1 ? tag_1_24 : _GEN_8755; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10169 = unuse_way == 2'h1 ? tag_1_25 : _GEN_8756; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10170 = unuse_way == 2'h1 ? tag_1_26 : _GEN_8757; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10171 = unuse_way == 2'h1 ? tag_1_27 : _GEN_8758; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10172 = unuse_way == 2'h1 ? tag_1_28 : _GEN_8759; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10173 = unuse_way == 2'h1 ? tag_1_29 : _GEN_8760; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10174 = unuse_way == 2'h1 ? tag_1_30 : _GEN_8761; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10175 = unuse_way == 2'h1 ? tag_1_31 : _GEN_8762; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10176 = unuse_way == 2'h1 ? tag_1_32 : _GEN_8763; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10177 = unuse_way == 2'h1 ? tag_1_33 : _GEN_8764; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10178 = unuse_way == 2'h1 ? tag_1_34 : _GEN_8765; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10179 = unuse_way == 2'h1 ? tag_1_35 : _GEN_8766; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10180 = unuse_way == 2'h1 ? tag_1_36 : _GEN_8767; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10181 = unuse_way == 2'h1 ? tag_1_37 : _GEN_8768; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10182 = unuse_way == 2'h1 ? tag_1_38 : _GEN_8769; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10183 = unuse_way == 2'h1 ? tag_1_39 : _GEN_8770; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10184 = unuse_way == 2'h1 ? tag_1_40 : _GEN_8771; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10185 = unuse_way == 2'h1 ? tag_1_41 : _GEN_8772; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10186 = unuse_way == 2'h1 ? tag_1_42 : _GEN_8773; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10187 = unuse_way == 2'h1 ? tag_1_43 : _GEN_8774; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10188 = unuse_way == 2'h1 ? tag_1_44 : _GEN_8775; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10189 = unuse_way == 2'h1 ? tag_1_45 : _GEN_8776; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10190 = unuse_way == 2'h1 ? tag_1_46 : _GEN_8777; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10191 = unuse_way == 2'h1 ? tag_1_47 : _GEN_8778; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10192 = unuse_way == 2'h1 ? tag_1_48 : _GEN_8779; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10193 = unuse_way == 2'h1 ? tag_1_49 : _GEN_8780; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10194 = unuse_way == 2'h1 ? tag_1_50 : _GEN_8781; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10195 = unuse_way == 2'h1 ? tag_1_51 : _GEN_8782; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10196 = unuse_way == 2'h1 ? tag_1_52 : _GEN_8783; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10197 = unuse_way == 2'h1 ? tag_1_53 : _GEN_8784; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10198 = unuse_way == 2'h1 ? tag_1_54 : _GEN_8785; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10199 = unuse_way == 2'h1 ? tag_1_55 : _GEN_8786; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10200 = unuse_way == 2'h1 ? tag_1_56 : _GEN_8787; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10201 = unuse_way == 2'h1 ? tag_1_57 : _GEN_8788; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10202 = unuse_way == 2'h1 ? tag_1_58 : _GEN_8789; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10203 = unuse_way == 2'h1 ? tag_1_59 : _GEN_8790; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10204 = unuse_way == 2'h1 ? tag_1_60 : _GEN_8791; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10205 = unuse_way == 2'h1 ? tag_1_61 : _GEN_8792; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10206 = unuse_way == 2'h1 ? tag_1_62 : _GEN_8793; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10207 = unuse_way == 2'h1 ? tag_1_63 : _GEN_8794; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10208 = unuse_way == 2'h1 ? tag_1_64 : _GEN_8795; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10209 = unuse_way == 2'h1 ? tag_1_65 : _GEN_8796; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10210 = unuse_way == 2'h1 ? tag_1_66 : _GEN_8797; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10211 = unuse_way == 2'h1 ? tag_1_67 : _GEN_8798; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10212 = unuse_way == 2'h1 ? tag_1_68 : _GEN_8799; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10213 = unuse_way == 2'h1 ? tag_1_69 : _GEN_8800; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10214 = unuse_way == 2'h1 ? tag_1_70 : _GEN_8801; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10215 = unuse_way == 2'h1 ? tag_1_71 : _GEN_8802; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10216 = unuse_way == 2'h1 ? tag_1_72 : _GEN_8803; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10217 = unuse_way == 2'h1 ? tag_1_73 : _GEN_8804; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10218 = unuse_way == 2'h1 ? tag_1_74 : _GEN_8805; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10219 = unuse_way == 2'h1 ? tag_1_75 : _GEN_8806; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10220 = unuse_way == 2'h1 ? tag_1_76 : _GEN_8807; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10221 = unuse_way == 2'h1 ? tag_1_77 : _GEN_8808; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10222 = unuse_way == 2'h1 ? tag_1_78 : _GEN_8809; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10223 = unuse_way == 2'h1 ? tag_1_79 : _GEN_8810; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10224 = unuse_way == 2'h1 ? tag_1_80 : _GEN_8811; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10225 = unuse_way == 2'h1 ? tag_1_81 : _GEN_8812; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10226 = unuse_way == 2'h1 ? tag_1_82 : _GEN_8813; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10227 = unuse_way == 2'h1 ? tag_1_83 : _GEN_8814; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10228 = unuse_way == 2'h1 ? tag_1_84 : _GEN_8815; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10229 = unuse_way == 2'h1 ? tag_1_85 : _GEN_8816; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10230 = unuse_way == 2'h1 ? tag_1_86 : _GEN_8817; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10231 = unuse_way == 2'h1 ? tag_1_87 : _GEN_8818; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10232 = unuse_way == 2'h1 ? tag_1_88 : _GEN_8819; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10233 = unuse_way == 2'h1 ? tag_1_89 : _GEN_8820; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10234 = unuse_way == 2'h1 ? tag_1_90 : _GEN_8821; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10235 = unuse_way == 2'h1 ? tag_1_91 : _GEN_8822; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10236 = unuse_way == 2'h1 ? tag_1_92 : _GEN_8823; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10237 = unuse_way == 2'h1 ? tag_1_93 : _GEN_8824; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10238 = unuse_way == 2'h1 ? tag_1_94 : _GEN_8825; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10239 = unuse_way == 2'h1 ? tag_1_95 : _GEN_8826; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10240 = unuse_way == 2'h1 ? tag_1_96 : _GEN_8827; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10241 = unuse_way == 2'h1 ? tag_1_97 : _GEN_8828; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10242 = unuse_way == 2'h1 ? tag_1_98 : _GEN_8829; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10243 = unuse_way == 2'h1 ? tag_1_99 : _GEN_8830; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10244 = unuse_way == 2'h1 ? tag_1_100 : _GEN_8831; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10245 = unuse_way == 2'h1 ? tag_1_101 : _GEN_8832; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10246 = unuse_way == 2'h1 ? tag_1_102 : _GEN_8833; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10247 = unuse_way == 2'h1 ? tag_1_103 : _GEN_8834; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10248 = unuse_way == 2'h1 ? tag_1_104 : _GEN_8835; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10249 = unuse_way == 2'h1 ? tag_1_105 : _GEN_8836; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10250 = unuse_way == 2'h1 ? tag_1_106 : _GEN_8837; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10251 = unuse_way == 2'h1 ? tag_1_107 : _GEN_8838; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10252 = unuse_way == 2'h1 ? tag_1_108 : _GEN_8839; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10253 = unuse_way == 2'h1 ? tag_1_109 : _GEN_8840; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10254 = unuse_way == 2'h1 ? tag_1_110 : _GEN_8841; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10255 = unuse_way == 2'h1 ? tag_1_111 : _GEN_8842; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10256 = unuse_way == 2'h1 ? tag_1_112 : _GEN_8843; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10257 = unuse_way == 2'h1 ? tag_1_113 : _GEN_8844; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10258 = unuse_way == 2'h1 ? tag_1_114 : _GEN_8845; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10259 = unuse_way == 2'h1 ? tag_1_115 : _GEN_8846; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10260 = unuse_way == 2'h1 ? tag_1_116 : _GEN_8847; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10261 = unuse_way == 2'h1 ? tag_1_117 : _GEN_8848; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10262 = unuse_way == 2'h1 ? tag_1_118 : _GEN_8849; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10263 = unuse_way == 2'h1 ? tag_1_119 : _GEN_8850; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10264 = unuse_way == 2'h1 ? tag_1_120 : _GEN_8851; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10265 = unuse_way == 2'h1 ? tag_1_121 : _GEN_8852; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10266 = unuse_way == 2'h1 ? tag_1_122 : _GEN_8853; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10267 = unuse_way == 2'h1 ? tag_1_123 : _GEN_8854; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10268 = unuse_way == 2'h1 ? tag_1_124 : _GEN_8855; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10269 = unuse_way == 2'h1 ? tag_1_125 : _GEN_8856; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10270 = unuse_way == 2'h1 ? tag_1_126 : _GEN_8857; // @[d_cache.scala 139:34 23:24]
  wire [31:0] _GEN_10271 = unuse_way == 2'h1 ? tag_1_127 : _GEN_8858; // @[d_cache.scala 139:34 23:24]
  wire  _GEN_10272 = unuse_way == 2'h1 ? valid_1_0 : _GEN_8859; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10273 = unuse_way == 2'h1 ? valid_1_1 : _GEN_8860; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10274 = unuse_way == 2'h1 ? valid_1_2 : _GEN_8861; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10275 = unuse_way == 2'h1 ? valid_1_3 : _GEN_8862; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10276 = unuse_way == 2'h1 ? valid_1_4 : _GEN_8863; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10277 = unuse_way == 2'h1 ? valid_1_5 : _GEN_8864; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10278 = unuse_way == 2'h1 ? valid_1_6 : _GEN_8865; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10279 = unuse_way == 2'h1 ? valid_1_7 : _GEN_8866; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10280 = unuse_way == 2'h1 ? valid_1_8 : _GEN_8867; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10281 = unuse_way == 2'h1 ? valid_1_9 : _GEN_8868; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10282 = unuse_way == 2'h1 ? valid_1_10 : _GEN_8869; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10283 = unuse_way == 2'h1 ? valid_1_11 : _GEN_8870; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10284 = unuse_way == 2'h1 ? valid_1_12 : _GEN_8871; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10285 = unuse_way == 2'h1 ? valid_1_13 : _GEN_8872; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10286 = unuse_way == 2'h1 ? valid_1_14 : _GEN_8873; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10287 = unuse_way == 2'h1 ? valid_1_15 : _GEN_8874; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10288 = unuse_way == 2'h1 ? valid_1_16 : _GEN_8875; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10289 = unuse_way == 2'h1 ? valid_1_17 : _GEN_8876; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10290 = unuse_way == 2'h1 ? valid_1_18 : _GEN_8877; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10291 = unuse_way == 2'h1 ? valid_1_19 : _GEN_8878; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10292 = unuse_way == 2'h1 ? valid_1_20 : _GEN_8879; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10293 = unuse_way == 2'h1 ? valid_1_21 : _GEN_8880; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10294 = unuse_way == 2'h1 ? valid_1_22 : _GEN_8881; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10295 = unuse_way == 2'h1 ? valid_1_23 : _GEN_8882; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10296 = unuse_way == 2'h1 ? valid_1_24 : _GEN_8883; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10297 = unuse_way == 2'h1 ? valid_1_25 : _GEN_8884; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10298 = unuse_way == 2'h1 ? valid_1_26 : _GEN_8885; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10299 = unuse_way == 2'h1 ? valid_1_27 : _GEN_8886; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10300 = unuse_way == 2'h1 ? valid_1_28 : _GEN_8887; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10301 = unuse_way == 2'h1 ? valid_1_29 : _GEN_8888; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10302 = unuse_way == 2'h1 ? valid_1_30 : _GEN_8889; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10303 = unuse_way == 2'h1 ? valid_1_31 : _GEN_8890; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10304 = unuse_way == 2'h1 ? valid_1_32 : _GEN_8891; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10305 = unuse_way == 2'h1 ? valid_1_33 : _GEN_8892; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10306 = unuse_way == 2'h1 ? valid_1_34 : _GEN_8893; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10307 = unuse_way == 2'h1 ? valid_1_35 : _GEN_8894; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10308 = unuse_way == 2'h1 ? valid_1_36 : _GEN_8895; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10309 = unuse_way == 2'h1 ? valid_1_37 : _GEN_8896; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10310 = unuse_way == 2'h1 ? valid_1_38 : _GEN_8897; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10311 = unuse_way == 2'h1 ? valid_1_39 : _GEN_8898; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10312 = unuse_way == 2'h1 ? valid_1_40 : _GEN_8899; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10313 = unuse_way == 2'h1 ? valid_1_41 : _GEN_8900; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10314 = unuse_way == 2'h1 ? valid_1_42 : _GEN_8901; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10315 = unuse_way == 2'h1 ? valid_1_43 : _GEN_8902; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10316 = unuse_way == 2'h1 ? valid_1_44 : _GEN_8903; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10317 = unuse_way == 2'h1 ? valid_1_45 : _GEN_8904; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10318 = unuse_way == 2'h1 ? valid_1_46 : _GEN_8905; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10319 = unuse_way == 2'h1 ? valid_1_47 : _GEN_8906; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10320 = unuse_way == 2'h1 ? valid_1_48 : _GEN_8907; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10321 = unuse_way == 2'h1 ? valid_1_49 : _GEN_8908; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10322 = unuse_way == 2'h1 ? valid_1_50 : _GEN_8909; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10323 = unuse_way == 2'h1 ? valid_1_51 : _GEN_8910; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10324 = unuse_way == 2'h1 ? valid_1_52 : _GEN_8911; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10325 = unuse_way == 2'h1 ? valid_1_53 : _GEN_8912; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10326 = unuse_way == 2'h1 ? valid_1_54 : _GEN_8913; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10327 = unuse_way == 2'h1 ? valid_1_55 : _GEN_8914; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10328 = unuse_way == 2'h1 ? valid_1_56 : _GEN_8915; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10329 = unuse_way == 2'h1 ? valid_1_57 : _GEN_8916; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10330 = unuse_way == 2'h1 ? valid_1_58 : _GEN_8917; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10331 = unuse_way == 2'h1 ? valid_1_59 : _GEN_8918; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10332 = unuse_way == 2'h1 ? valid_1_60 : _GEN_8919; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10333 = unuse_way == 2'h1 ? valid_1_61 : _GEN_8920; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10334 = unuse_way == 2'h1 ? valid_1_62 : _GEN_8921; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10335 = unuse_way == 2'h1 ? valid_1_63 : _GEN_8922; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10336 = unuse_way == 2'h1 ? valid_1_64 : _GEN_8923; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10337 = unuse_way == 2'h1 ? valid_1_65 : _GEN_8924; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10338 = unuse_way == 2'h1 ? valid_1_66 : _GEN_8925; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10339 = unuse_way == 2'h1 ? valid_1_67 : _GEN_8926; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10340 = unuse_way == 2'h1 ? valid_1_68 : _GEN_8927; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10341 = unuse_way == 2'h1 ? valid_1_69 : _GEN_8928; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10342 = unuse_way == 2'h1 ? valid_1_70 : _GEN_8929; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10343 = unuse_way == 2'h1 ? valid_1_71 : _GEN_8930; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10344 = unuse_way == 2'h1 ? valid_1_72 : _GEN_8931; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10345 = unuse_way == 2'h1 ? valid_1_73 : _GEN_8932; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10346 = unuse_way == 2'h1 ? valid_1_74 : _GEN_8933; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10347 = unuse_way == 2'h1 ? valid_1_75 : _GEN_8934; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10348 = unuse_way == 2'h1 ? valid_1_76 : _GEN_8935; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10349 = unuse_way == 2'h1 ? valid_1_77 : _GEN_8936; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10350 = unuse_way == 2'h1 ? valid_1_78 : _GEN_8937; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10351 = unuse_way == 2'h1 ? valid_1_79 : _GEN_8938; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10352 = unuse_way == 2'h1 ? valid_1_80 : _GEN_8939; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10353 = unuse_way == 2'h1 ? valid_1_81 : _GEN_8940; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10354 = unuse_way == 2'h1 ? valid_1_82 : _GEN_8941; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10355 = unuse_way == 2'h1 ? valid_1_83 : _GEN_8942; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10356 = unuse_way == 2'h1 ? valid_1_84 : _GEN_8943; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10357 = unuse_way == 2'h1 ? valid_1_85 : _GEN_8944; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10358 = unuse_way == 2'h1 ? valid_1_86 : _GEN_8945; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10359 = unuse_way == 2'h1 ? valid_1_87 : _GEN_8946; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10360 = unuse_way == 2'h1 ? valid_1_88 : _GEN_8947; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10361 = unuse_way == 2'h1 ? valid_1_89 : _GEN_8948; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10362 = unuse_way == 2'h1 ? valid_1_90 : _GEN_8949; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10363 = unuse_way == 2'h1 ? valid_1_91 : _GEN_8950; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10364 = unuse_way == 2'h1 ? valid_1_92 : _GEN_8951; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10365 = unuse_way == 2'h1 ? valid_1_93 : _GEN_8952; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10366 = unuse_way == 2'h1 ? valid_1_94 : _GEN_8953; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10367 = unuse_way == 2'h1 ? valid_1_95 : _GEN_8954; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10368 = unuse_way == 2'h1 ? valid_1_96 : _GEN_8955; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10369 = unuse_way == 2'h1 ? valid_1_97 : _GEN_8956; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10370 = unuse_way == 2'h1 ? valid_1_98 : _GEN_8957; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10371 = unuse_way == 2'h1 ? valid_1_99 : _GEN_8958; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10372 = unuse_way == 2'h1 ? valid_1_100 : _GEN_8959; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10373 = unuse_way == 2'h1 ? valid_1_101 : _GEN_8960; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10374 = unuse_way == 2'h1 ? valid_1_102 : _GEN_8961; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10375 = unuse_way == 2'h1 ? valid_1_103 : _GEN_8962; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10376 = unuse_way == 2'h1 ? valid_1_104 : _GEN_8963; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10377 = unuse_way == 2'h1 ? valid_1_105 : _GEN_8964; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10378 = unuse_way == 2'h1 ? valid_1_106 : _GEN_8965; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10379 = unuse_way == 2'h1 ? valid_1_107 : _GEN_8966; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10380 = unuse_way == 2'h1 ? valid_1_108 : _GEN_8967; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10381 = unuse_way == 2'h1 ? valid_1_109 : _GEN_8968; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10382 = unuse_way == 2'h1 ? valid_1_110 : _GEN_8969; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10383 = unuse_way == 2'h1 ? valid_1_111 : _GEN_8970; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10384 = unuse_way == 2'h1 ? valid_1_112 : _GEN_8971; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10385 = unuse_way == 2'h1 ? valid_1_113 : _GEN_8972; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10386 = unuse_way == 2'h1 ? valid_1_114 : _GEN_8973; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10387 = unuse_way == 2'h1 ? valid_1_115 : _GEN_8974; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10388 = unuse_way == 2'h1 ? valid_1_116 : _GEN_8975; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10389 = unuse_way == 2'h1 ? valid_1_117 : _GEN_8976; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10390 = unuse_way == 2'h1 ? valid_1_118 : _GEN_8977; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10391 = unuse_way == 2'h1 ? valid_1_119 : _GEN_8978; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10392 = unuse_way == 2'h1 ? valid_1_120 : _GEN_8979; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10393 = unuse_way == 2'h1 ? valid_1_121 : _GEN_8980; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10394 = unuse_way == 2'h1 ? valid_1_122 : _GEN_8981; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10395 = unuse_way == 2'h1 ? valid_1_123 : _GEN_8982; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10396 = unuse_way == 2'h1 ? valid_1_124 : _GEN_8983; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10397 = unuse_way == 2'h1 ? valid_1_125 : _GEN_8984; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10398 = unuse_way == 2'h1 ? valid_1_126 : _GEN_8985; // @[d_cache.scala 139:34 25:26]
  wire  _GEN_10399 = unuse_way == 2'h1 ? valid_1_127 : _GEN_8986; // @[d_cache.scala 139:34 25:26]
  wire [63:0] _GEN_10400 = unuse_way == 2'h1 ? write_back_data : _GEN_8988; // @[d_cache.scala 139:34 31:34]
  wire [41:0] _GEN_10401 = unuse_way == 2'h1 ? {{10'd0}, write_back_addr} : _GEN_8989; // @[d_cache.scala 139:34 32:34]
  wire  _GEN_10402 = unuse_way == 2'h1 ? dirty_0_0 : _GEN_9246; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10403 = unuse_way == 2'h1 ? dirty_0_1 : _GEN_9247; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10404 = unuse_way == 2'h1 ? dirty_0_2 : _GEN_9248; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10405 = unuse_way == 2'h1 ? dirty_0_3 : _GEN_9249; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10406 = unuse_way == 2'h1 ? dirty_0_4 : _GEN_9250; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10407 = unuse_way == 2'h1 ? dirty_0_5 : _GEN_9251; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10408 = unuse_way == 2'h1 ? dirty_0_6 : _GEN_9252; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10409 = unuse_way == 2'h1 ? dirty_0_7 : _GEN_9253; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10410 = unuse_way == 2'h1 ? dirty_0_8 : _GEN_9254; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10411 = unuse_way == 2'h1 ? dirty_0_9 : _GEN_9255; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10412 = unuse_way == 2'h1 ? dirty_0_10 : _GEN_9256; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10413 = unuse_way == 2'h1 ? dirty_0_11 : _GEN_9257; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10414 = unuse_way == 2'h1 ? dirty_0_12 : _GEN_9258; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10415 = unuse_way == 2'h1 ? dirty_0_13 : _GEN_9259; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10416 = unuse_way == 2'h1 ? dirty_0_14 : _GEN_9260; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10417 = unuse_way == 2'h1 ? dirty_0_15 : _GEN_9261; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10418 = unuse_way == 2'h1 ? dirty_0_16 : _GEN_9262; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10419 = unuse_way == 2'h1 ? dirty_0_17 : _GEN_9263; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10420 = unuse_way == 2'h1 ? dirty_0_18 : _GEN_9264; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10421 = unuse_way == 2'h1 ? dirty_0_19 : _GEN_9265; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10422 = unuse_way == 2'h1 ? dirty_0_20 : _GEN_9266; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10423 = unuse_way == 2'h1 ? dirty_0_21 : _GEN_9267; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10424 = unuse_way == 2'h1 ? dirty_0_22 : _GEN_9268; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10425 = unuse_way == 2'h1 ? dirty_0_23 : _GEN_9269; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10426 = unuse_way == 2'h1 ? dirty_0_24 : _GEN_9270; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10427 = unuse_way == 2'h1 ? dirty_0_25 : _GEN_9271; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10428 = unuse_way == 2'h1 ? dirty_0_26 : _GEN_9272; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10429 = unuse_way == 2'h1 ? dirty_0_27 : _GEN_9273; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10430 = unuse_way == 2'h1 ? dirty_0_28 : _GEN_9274; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10431 = unuse_way == 2'h1 ? dirty_0_29 : _GEN_9275; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10432 = unuse_way == 2'h1 ? dirty_0_30 : _GEN_9276; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10433 = unuse_way == 2'h1 ? dirty_0_31 : _GEN_9277; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10434 = unuse_way == 2'h1 ? dirty_0_32 : _GEN_9278; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10435 = unuse_way == 2'h1 ? dirty_0_33 : _GEN_9279; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10436 = unuse_way == 2'h1 ? dirty_0_34 : _GEN_9280; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10437 = unuse_way == 2'h1 ? dirty_0_35 : _GEN_9281; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10438 = unuse_way == 2'h1 ? dirty_0_36 : _GEN_9282; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10439 = unuse_way == 2'h1 ? dirty_0_37 : _GEN_9283; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10440 = unuse_way == 2'h1 ? dirty_0_38 : _GEN_9284; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10441 = unuse_way == 2'h1 ? dirty_0_39 : _GEN_9285; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10442 = unuse_way == 2'h1 ? dirty_0_40 : _GEN_9286; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10443 = unuse_way == 2'h1 ? dirty_0_41 : _GEN_9287; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10444 = unuse_way == 2'h1 ? dirty_0_42 : _GEN_9288; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10445 = unuse_way == 2'h1 ? dirty_0_43 : _GEN_9289; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10446 = unuse_way == 2'h1 ? dirty_0_44 : _GEN_9290; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10447 = unuse_way == 2'h1 ? dirty_0_45 : _GEN_9291; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10448 = unuse_way == 2'h1 ? dirty_0_46 : _GEN_9292; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10449 = unuse_way == 2'h1 ? dirty_0_47 : _GEN_9293; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10450 = unuse_way == 2'h1 ? dirty_0_48 : _GEN_9294; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10451 = unuse_way == 2'h1 ? dirty_0_49 : _GEN_9295; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10452 = unuse_way == 2'h1 ? dirty_0_50 : _GEN_9296; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10453 = unuse_way == 2'h1 ? dirty_0_51 : _GEN_9297; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10454 = unuse_way == 2'h1 ? dirty_0_52 : _GEN_9298; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10455 = unuse_way == 2'h1 ? dirty_0_53 : _GEN_9299; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10456 = unuse_way == 2'h1 ? dirty_0_54 : _GEN_9300; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10457 = unuse_way == 2'h1 ? dirty_0_55 : _GEN_9301; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10458 = unuse_way == 2'h1 ? dirty_0_56 : _GEN_9302; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10459 = unuse_way == 2'h1 ? dirty_0_57 : _GEN_9303; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10460 = unuse_way == 2'h1 ? dirty_0_58 : _GEN_9304; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10461 = unuse_way == 2'h1 ? dirty_0_59 : _GEN_9305; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10462 = unuse_way == 2'h1 ? dirty_0_60 : _GEN_9306; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10463 = unuse_way == 2'h1 ? dirty_0_61 : _GEN_9307; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10464 = unuse_way == 2'h1 ? dirty_0_62 : _GEN_9308; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10465 = unuse_way == 2'h1 ? dirty_0_63 : _GEN_9309; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10466 = unuse_way == 2'h1 ? dirty_0_64 : _GEN_9310; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10467 = unuse_way == 2'h1 ? dirty_0_65 : _GEN_9311; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10468 = unuse_way == 2'h1 ? dirty_0_66 : _GEN_9312; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10469 = unuse_way == 2'h1 ? dirty_0_67 : _GEN_9313; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10470 = unuse_way == 2'h1 ? dirty_0_68 : _GEN_9314; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10471 = unuse_way == 2'h1 ? dirty_0_69 : _GEN_9315; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10472 = unuse_way == 2'h1 ? dirty_0_70 : _GEN_9316; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10473 = unuse_way == 2'h1 ? dirty_0_71 : _GEN_9317; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10474 = unuse_way == 2'h1 ? dirty_0_72 : _GEN_9318; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10475 = unuse_way == 2'h1 ? dirty_0_73 : _GEN_9319; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10476 = unuse_way == 2'h1 ? dirty_0_74 : _GEN_9320; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10477 = unuse_way == 2'h1 ? dirty_0_75 : _GEN_9321; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10478 = unuse_way == 2'h1 ? dirty_0_76 : _GEN_9322; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10479 = unuse_way == 2'h1 ? dirty_0_77 : _GEN_9323; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10480 = unuse_way == 2'h1 ? dirty_0_78 : _GEN_9324; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10481 = unuse_way == 2'h1 ? dirty_0_79 : _GEN_9325; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10482 = unuse_way == 2'h1 ? dirty_0_80 : _GEN_9326; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10483 = unuse_way == 2'h1 ? dirty_0_81 : _GEN_9327; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10484 = unuse_way == 2'h1 ? dirty_0_82 : _GEN_9328; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10485 = unuse_way == 2'h1 ? dirty_0_83 : _GEN_9329; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10486 = unuse_way == 2'h1 ? dirty_0_84 : _GEN_9330; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10487 = unuse_way == 2'h1 ? dirty_0_85 : _GEN_9331; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10488 = unuse_way == 2'h1 ? dirty_0_86 : _GEN_9332; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10489 = unuse_way == 2'h1 ? dirty_0_87 : _GEN_9333; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10490 = unuse_way == 2'h1 ? dirty_0_88 : _GEN_9334; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10491 = unuse_way == 2'h1 ? dirty_0_89 : _GEN_9335; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10492 = unuse_way == 2'h1 ? dirty_0_90 : _GEN_9336; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10493 = unuse_way == 2'h1 ? dirty_0_91 : _GEN_9337; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10494 = unuse_way == 2'h1 ? dirty_0_92 : _GEN_9338; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10495 = unuse_way == 2'h1 ? dirty_0_93 : _GEN_9339; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10496 = unuse_way == 2'h1 ? dirty_0_94 : _GEN_9340; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10497 = unuse_way == 2'h1 ? dirty_0_95 : _GEN_9341; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10498 = unuse_way == 2'h1 ? dirty_0_96 : _GEN_9342; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10499 = unuse_way == 2'h1 ? dirty_0_97 : _GEN_9343; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10500 = unuse_way == 2'h1 ? dirty_0_98 : _GEN_9344; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10501 = unuse_way == 2'h1 ? dirty_0_99 : _GEN_9345; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10502 = unuse_way == 2'h1 ? dirty_0_100 : _GEN_9346; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10503 = unuse_way == 2'h1 ? dirty_0_101 : _GEN_9347; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10504 = unuse_way == 2'h1 ? dirty_0_102 : _GEN_9348; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10505 = unuse_way == 2'h1 ? dirty_0_103 : _GEN_9349; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10506 = unuse_way == 2'h1 ? dirty_0_104 : _GEN_9350; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10507 = unuse_way == 2'h1 ? dirty_0_105 : _GEN_9351; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10508 = unuse_way == 2'h1 ? dirty_0_106 : _GEN_9352; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10509 = unuse_way == 2'h1 ? dirty_0_107 : _GEN_9353; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10510 = unuse_way == 2'h1 ? dirty_0_108 : _GEN_9354; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10511 = unuse_way == 2'h1 ? dirty_0_109 : _GEN_9355; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10512 = unuse_way == 2'h1 ? dirty_0_110 : _GEN_9356; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10513 = unuse_way == 2'h1 ? dirty_0_111 : _GEN_9357; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10514 = unuse_way == 2'h1 ? dirty_0_112 : _GEN_9358; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10515 = unuse_way == 2'h1 ? dirty_0_113 : _GEN_9359; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10516 = unuse_way == 2'h1 ? dirty_0_114 : _GEN_9360; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10517 = unuse_way == 2'h1 ? dirty_0_115 : _GEN_9361; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10518 = unuse_way == 2'h1 ? dirty_0_116 : _GEN_9362; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10519 = unuse_way == 2'h1 ? dirty_0_117 : _GEN_9363; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10520 = unuse_way == 2'h1 ? dirty_0_118 : _GEN_9364; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10521 = unuse_way == 2'h1 ? dirty_0_119 : _GEN_9365; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10522 = unuse_way == 2'h1 ? dirty_0_120 : _GEN_9366; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10523 = unuse_way == 2'h1 ? dirty_0_121 : _GEN_9367; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10524 = unuse_way == 2'h1 ? dirty_0_122 : _GEN_9368; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10525 = unuse_way == 2'h1 ? dirty_0_123 : _GEN_9369; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10526 = unuse_way == 2'h1 ? dirty_0_124 : _GEN_9370; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10527 = unuse_way == 2'h1 ? dirty_0_125 : _GEN_9371; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10528 = unuse_way == 2'h1 ? dirty_0_126 : _GEN_9372; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10529 = unuse_way == 2'h1 ? dirty_0_127 : _GEN_9373; // @[d_cache.scala 139:34 26:26]
  wire  _GEN_10530 = unuse_way == 2'h1 ? dirty_1_0 : _GEN_9502; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10531 = unuse_way == 2'h1 ? dirty_1_1 : _GEN_9503; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10532 = unuse_way == 2'h1 ? dirty_1_2 : _GEN_9504; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10533 = unuse_way == 2'h1 ? dirty_1_3 : _GEN_9505; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10534 = unuse_way == 2'h1 ? dirty_1_4 : _GEN_9506; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10535 = unuse_way == 2'h1 ? dirty_1_5 : _GEN_9507; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10536 = unuse_way == 2'h1 ? dirty_1_6 : _GEN_9508; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10537 = unuse_way == 2'h1 ? dirty_1_7 : _GEN_9509; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10538 = unuse_way == 2'h1 ? dirty_1_8 : _GEN_9510; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10539 = unuse_way == 2'h1 ? dirty_1_9 : _GEN_9511; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10540 = unuse_way == 2'h1 ? dirty_1_10 : _GEN_9512; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10541 = unuse_way == 2'h1 ? dirty_1_11 : _GEN_9513; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10542 = unuse_way == 2'h1 ? dirty_1_12 : _GEN_9514; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10543 = unuse_way == 2'h1 ? dirty_1_13 : _GEN_9515; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10544 = unuse_way == 2'h1 ? dirty_1_14 : _GEN_9516; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10545 = unuse_way == 2'h1 ? dirty_1_15 : _GEN_9517; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10546 = unuse_way == 2'h1 ? dirty_1_16 : _GEN_9518; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10547 = unuse_way == 2'h1 ? dirty_1_17 : _GEN_9519; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10548 = unuse_way == 2'h1 ? dirty_1_18 : _GEN_9520; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10549 = unuse_way == 2'h1 ? dirty_1_19 : _GEN_9521; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10550 = unuse_way == 2'h1 ? dirty_1_20 : _GEN_9522; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10551 = unuse_way == 2'h1 ? dirty_1_21 : _GEN_9523; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10552 = unuse_way == 2'h1 ? dirty_1_22 : _GEN_9524; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10553 = unuse_way == 2'h1 ? dirty_1_23 : _GEN_9525; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10554 = unuse_way == 2'h1 ? dirty_1_24 : _GEN_9526; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10555 = unuse_way == 2'h1 ? dirty_1_25 : _GEN_9527; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10556 = unuse_way == 2'h1 ? dirty_1_26 : _GEN_9528; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10557 = unuse_way == 2'h1 ? dirty_1_27 : _GEN_9529; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10558 = unuse_way == 2'h1 ? dirty_1_28 : _GEN_9530; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10559 = unuse_way == 2'h1 ? dirty_1_29 : _GEN_9531; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10560 = unuse_way == 2'h1 ? dirty_1_30 : _GEN_9532; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10561 = unuse_way == 2'h1 ? dirty_1_31 : _GEN_9533; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10562 = unuse_way == 2'h1 ? dirty_1_32 : _GEN_9534; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10563 = unuse_way == 2'h1 ? dirty_1_33 : _GEN_9535; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10564 = unuse_way == 2'h1 ? dirty_1_34 : _GEN_9536; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10565 = unuse_way == 2'h1 ? dirty_1_35 : _GEN_9537; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10566 = unuse_way == 2'h1 ? dirty_1_36 : _GEN_9538; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10567 = unuse_way == 2'h1 ? dirty_1_37 : _GEN_9539; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10568 = unuse_way == 2'h1 ? dirty_1_38 : _GEN_9540; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10569 = unuse_way == 2'h1 ? dirty_1_39 : _GEN_9541; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10570 = unuse_way == 2'h1 ? dirty_1_40 : _GEN_9542; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10571 = unuse_way == 2'h1 ? dirty_1_41 : _GEN_9543; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10572 = unuse_way == 2'h1 ? dirty_1_42 : _GEN_9544; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10573 = unuse_way == 2'h1 ? dirty_1_43 : _GEN_9545; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10574 = unuse_way == 2'h1 ? dirty_1_44 : _GEN_9546; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10575 = unuse_way == 2'h1 ? dirty_1_45 : _GEN_9547; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10576 = unuse_way == 2'h1 ? dirty_1_46 : _GEN_9548; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10577 = unuse_way == 2'h1 ? dirty_1_47 : _GEN_9549; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10578 = unuse_way == 2'h1 ? dirty_1_48 : _GEN_9550; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10579 = unuse_way == 2'h1 ? dirty_1_49 : _GEN_9551; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10580 = unuse_way == 2'h1 ? dirty_1_50 : _GEN_9552; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10581 = unuse_way == 2'h1 ? dirty_1_51 : _GEN_9553; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10582 = unuse_way == 2'h1 ? dirty_1_52 : _GEN_9554; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10583 = unuse_way == 2'h1 ? dirty_1_53 : _GEN_9555; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10584 = unuse_way == 2'h1 ? dirty_1_54 : _GEN_9556; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10585 = unuse_way == 2'h1 ? dirty_1_55 : _GEN_9557; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10586 = unuse_way == 2'h1 ? dirty_1_56 : _GEN_9558; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10587 = unuse_way == 2'h1 ? dirty_1_57 : _GEN_9559; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10588 = unuse_way == 2'h1 ? dirty_1_58 : _GEN_9560; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10589 = unuse_way == 2'h1 ? dirty_1_59 : _GEN_9561; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10590 = unuse_way == 2'h1 ? dirty_1_60 : _GEN_9562; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10591 = unuse_way == 2'h1 ? dirty_1_61 : _GEN_9563; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10592 = unuse_way == 2'h1 ? dirty_1_62 : _GEN_9564; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10593 = unuse_way == 2'h1 ? dirty_1_63 : _GEN_9565; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10594 = unuse_way == 2'h1 ? dirty_1_64 : _GEN_9566; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10595 = unuse_way == 2'h1 ? dirty_1_65 : _GEN_9567; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10596 = unuse_way == 2'h1 ? dirty_1_66 : _GEN_9568; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10597 = unuse_way == 2'h1 ? dirty_1_67 : _GEN_9569; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10598 = unuse_way == 2'h1 ? dirty_1_68 : _GEN_9570; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10599 = unuse_way == 2'h1 ? dirty_1_69 : _GEN_9571; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10600 = unuse_way == 2'h1 ? dirty_1_70 : _GEN_9572; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10601 = unuse_way == 2'h1 ? dirty_1_71 : _GEN_9573; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10602 = unuse_way == 2'h1 ? dirty_1_72 : _GEN_9574; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10603 = unuse_way == 2'h1 ? dirty_1_73 : _GEN_9575; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10604 = unuse_way == 2'h1 ? dirty_1_74 : _GEN_9576; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10605 = unuse_way == 2'h1 ? dirty_1_75 : _GEN_9577; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10606 = unuse_way == 2'h1 ? dirty_1_76 : _GEN_9578; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10607 = unuse_way == 2'h1 ? dirty_1_77 : _GEN_9579; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10608 = unuse_way == 2'h1 ? dirty_1_78 : _GEN_9580; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10609 = unuse_way == 2'h1 ? dirty_1_79 : _GEN_9581; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10610 = unuse_way == 2'h1 ? dirty_1_80 : _GEN_9582; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10611 = unuse_way == 2'h1 ? dirty_1_81 : _GEN_9583; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10612 = unuse_way == 2'h1 ? dirty_1_82 : _GEN_9584; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10613 = unuse_way == 2'h1 ? dirty_1_83 : _GEN_9585; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10614 = unuse_way == 2'h1 ? dirty_1_84 : _GEN_9586; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10615 = unuse_way == 2'h1 ? dirty_1_85 : _GEN_9587; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10616 = unuse_way == 2'h1 ? dirty_1_86 : _GEN_9588; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10617 = unuse_way == 2'h1 ? dirty_1_87 : _GEN_9589; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10618 = unuse_way == 2'h1 ? dirty_1_88 : _GEN_9590; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10619 = unuse_way == 2'h1 ? dirty_1_89 : _GEN_9591; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10620 = unuse_way == 2'h1 ? dirty_1_90 : _GEN_9592; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10621 = unuse_way == 2'h1 ? dirty_1_91 : _GEN_9593; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10622 = unuse_way == 2'h1 ? dirty_1_92 : _GEN_9594; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10623 = unuse_way == 2'h1 ? dirty_1_93 : _GEN_9595; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10624 = unuse_way == 2'h1 ? dirty_1_94 : _GEN_9596; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10625 = unuse_way == 2'h1 ? dirty_1_95 : _GEN_9597; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10626 = unuse_way == 2'h1 ? dirty_1_96 : _GEN_9598; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10627 = unuse_way == 2'h1 ? dirty_1_97 : _GEN_9599; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10628 = unuse_way == 2'h1 ? dirty_1_98 : _GEN_9600; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10629 = unuse_way == 2'h1 ? dirty_1_99 : _GEN_9601; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10630 = unuse_way == 2'h1 ? dirty_1_100 : _GEN_9602; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10631 = unuse_way == 2'h1 ? dirty_1_101 : _GEN_9603; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10632 = unuse_way == 2'h1 ? dirty_1_102 : _GEN_9604; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10633 = unuse_way == 2'h1 ? dirty_1_103 : _GEN_9605; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10634 = unuse_way == 2'h1 ? dirty_1_104 : _GEN_9606; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10635 = unuse_way == 2'h1 ? dirty_1_105 : _GEN_9607; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10636 = unuse_way == 2'h1 ? dirty_1_106 : _GEN_9608; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10637 = unuse_way == 2'h1 ? dirty_1_107 : _GEN_9609; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10638 = unuse_way == 2'h1 ? dirty_1_108 : _GEN_9610; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10639 = unuse_way == 2'h1 ? dirty_1_109 : _GEN_9611; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10640 = unuse_way == 2'h1 ? dirty_1_110 : _GEN_9612; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10641 = unuse_way == 2'h1 ? dirty_1_111 : _GEN_9613; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10642 = unuse_way == 2'h1 ? dirty_1_112 : _GEN_9614; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10643 = unuse_way == 2'h1 ? dirty_1_113 : _GEN_9615; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10644 = unuse_way == 2'h1 ? dirty_1_114 : _GEN_9616; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10645 = unuse_way == 2'h1 ? dirty_1_115 : _GEN_9617; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10646 = unuse_way == 2'h1 ? dirty_1_116 : _GEN_9618; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10647 = unuse_way == 2'h1 ? dirty_1_117 : _GEN_9619; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10648 = unuse_way == 2'h1 ? dirty_1_118 : _GEN_9620; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10649 = unuse_way == 2'h1 ? dirty_1_119 : _GEN_9621; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10650 = unuse_way == 2'h1 ? dirty_1_120 : _GEN_9622; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10651 = unuse_way == 2'h1 ? dirty_1_121 : _GEN_9623; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10652 = unuse_way == 2'h1 ? dirty_1_122 : _GEN_9624; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10653 = unuse_way == 2'h1 ? dirty_1_123 : _GEN_9625; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10654 = unuse_way == 2'h1 ? dirty_1_124 : _GEN_9626; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10655 = unuse_way == 2'h1 ? dirty_1_125 : _GEN_9627; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10656 = unuse_way == 2'h1 ? dirty_1_126 : _GEN_9628; // @[d_cache.scala 139:34 27:26]
  wire  _GEN_10657 = unuse_way == 2'h1 ? dirty_1_127 : _GEN_9629; // @[d_cache.scala 139:34 27:26]
  wire [2:0] _GEN_10658 = io_from_axi_bvalid ? 3'h7 : state; // @[d_cache.scala 191:37 192:23 76:24]
  wire [2:0] _GEN_10659 = 3'h7 == state ? 3'h1 : state; // @[d_cache.scala 81:18 196:19 76:24]
  wire [2:0] _GEN_10660 = 3'h6 == state ? _GEN_10658 : _GEN_10659; // @[d_cache.scala 81:18]
  wire [2:0] _GEN_10661 = 3'h5 == state ? _GEN_9630 : _GEN_10660; // @[d_cache.scala 81:18]
  wire [63:0] _GEN_10662 = 3'h5 == state ? _GEN_9631 : ram_0_0; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10663 = 3'h5 == state ? _GEN_9632 : ram_0_1; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10664 = 3'h5 == state ? _GEN_9633 : ram_0_2; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10665 = 3'h5 == state ? _GEN_9634 : ram_0_3; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10666 = 3'h5 == state ? _GEN_9635 : ram_0_4; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10667 = 3'h5 == state ? _GEN_9636 : ram_0_5; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10668 = 3'h5 == state ? _GEN_9637 : ram_0_6; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10669 = 3'h5 == state ? _GEN_9638 : ram_0_7; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10670 = 3'h5 == state ? _GEN_9639 : ram_0_8; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10671 = 3'h5 == state ? _GEN_9640 : ram_0_9; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10672 = 3'h5 == state ? _GEN_9641 : ram_0_10; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10673 = 3'h5 == state ? _GEN_9642 : ram_0_11; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10674 = 3'h5 == state ? _GEN_9643 : ram_0_12; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10675 = 3'h5 == state ? _GEN_9644 : ram_0_13; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10676 = 3'h5 == state ? _GEN_9645 : ram_0_14; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10677 = 3'h5 == state ? _GEN_9646 : ram_0_15; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10678 = 3'h5 == state ? _GEN_9647 : ram_0_16; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10679 = 3'h5 == state ? _GEN_9648 : ram_0_17; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10680 = 3'h5 == state ? _GEN_9649 : ram_0_18; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10681 = 3'h5 == state ? _GEN_9650 : ram_0_19; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10682 = 3'h5 == state ? _GEN_9651 : ram_0_20; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10683 = 3'h5 == state ? _GEN_9652 : ram_0_21; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10684 = 3'h5 == state ? _GEN_9653 : ram_0_22; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10685 = 3'h5 == state ? _GEN_9654 : ram_0_23; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10686 = 3'h5 == state ? _GEN_9655 : ram_0_24; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10687 = 3'h5 == state ? _GEN_9656 : ram_0_25; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10688 = 3'h5 == state ? _GEN_9657 : ram_0_26; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10689 = 3'h5 == state ? _GEN_9658 : ram_0_27; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10690 = 3'h5 == state ? _GEN_9659 : ram_0_28; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10691 = 3'h5 == state ? _GEN_9660 : ram_0_29; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10692 = 3'h5 == state ? _GEN_9661 : ram_0_30; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10693 = 3'h5 == state ? _GEN_9662 : ram_0_31; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10694 = 3'h5 == state ? _GEN_9663 : ram_0_32; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10695 = 3'h5 == state ? _GEN_9664 : ram_0_33; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10696 = 3'h5 == state ? _GEN_9665 : ram_0_34; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10697 = 3'h5 == state ? _GEN_9666 : ram_0_35; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10698 = 3'h5 == state ? _GEN_9667 : ram_0_36; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10699 = 3'h5 == state ? _GEN_9668 : ram_0_37; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10700 = 3'h5 == state ? _GEN_9669 : ram_0_38; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10701 = 3'h5 == state ? _GEN_9670 : ram_0_39; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10702 = 3'h5 == state ? _GEN_9671 : ram_0_40; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10703 = 3'h5 == state ? _GEN_9672 : ram_0_41; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10704 = 3'h5 == state ? _GEN_9673 : ram_0_42; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10705 = 3'h5 == state ? _GEN_9674 : ram_0_43; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10706 = 3'h5 == state ? _GEN_9675 : ram_0_44; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10707 = 3'h5 == state ? _GEN_9676 : ram_0_45; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10708 = 3'h5 == state ? _GEN_9677 : ram_0_46; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10709 = 3'h5 == state ? _GEN_9678 : ram_0_47; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10710 = 3'h5 == state ? _GEN_9679 : ram_0_48; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10711 = 3'h5 == state ? _GEN_9680 : ram_0_49; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10712 = 3'h5 == state ? _GEN_9681 : ram_0_50; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10713 = 3'h5 == state ? _GEN_9682 : ram_0_51; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10714 = 3'h5 == state ? _GEN_9683 : ram_0_52; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10715 = 3'h5 == state ? _GEN_9684 : ram_0_53; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10716 = 3'h5 == state ? _GEN_9685 : ram_0_54; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10717 = 3'h5 == state ? _GEN_9686 : ram_0_55; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10718 = 3'h5 == state ? _GEN_9687 : ram_0_56; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10719 = 3'h5 == state ? _GEN_9688 : ram_0_57; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10720 = 3'h5 == state ? _GEN_9689 : ram_0_58; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10721 = 3'h5 == state ? _GEN_9690 : ram_0_59; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10722 = 3'h5 == state ? _GEN_9691 : ram_0_60; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10723 = 3'h5 == state ? _GEN_9692 : ram_0_61; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10724 = 3'h5 == state ? _GEN_9693 : ram_0_62; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10725 = 3'h5 == state ? _GEN_9694 : ram_0_63; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10726 = 3'h5 == state ? _GEN_9695 : ram_0_64; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10727 = 3'h5 == state ? _GEN_9696 : ram_0_65; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10728 = 3'h5 == state ? _GEN_9697 : ram_0_66; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10729 = 3'h5 == state ? _GEN_9698 : ram_0_67; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10730 = 3'h5 == state ? _GEN_9699 : ram_0_68; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10731 = 3'h5 == state ? _GEN_9700 : ram_0_69; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10732 = 3'h5 == state ? _GEN_9701 : ram_0_70; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10733 = 3'h5 == state ? _GEN_9702 : ram_0_71; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10734 = 3'h5 == state ? _GEN_9703 : ram_0_72; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10735 = 3'h5 == state ? _GEN_9704 : ram_0_73; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10736 = 3'h5 == state ? _GEN_9705 : ram_0_74; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10737 = 3'h5 == state ? _GEN_9706 : ram_0_75; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10738 = 3'h5 == state ? _GEN_9707 : ram_0_76; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10739 = 3'h5 == state ? _GEN_9708 : ram_0_77; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10740 = 3'h5 == state ? _GEN_9709 : ram_0_78; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10741 = 3'h5 == state ? _GEN_9710 : ram_0_79; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10742 = 3'h5 == state ? _GEN_9711 : ram_0_80; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10743 = 3'h5 == state ? _GEN_9712 : ram_0_81; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10744 = 3'h5 == state ? _GEN_9713 : ram_0_82; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10745 = 3'h5 == state ? _GEN_9714 : ram_0_83; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10746 = 3'h5 == state ? _GEN_9715 : ram_0_84; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10747 = 3'h5 == state ? _GEN_9716 : ram_0_85; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10748 = 3'h5 == state ? _GEN_9717 : ram_0_86; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10749 = 3'h5 == state ? _GEN_9718 : ram_0_87; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10750 = 3'h5 == state ? _GEN_9719 : ram_0_88; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10751 = 3'h5 == state ? _GEN_9720 : ram_0_89; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10752 = 3'h5 == state ? _GEN_9721 : ram_0_90; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10753 = 3'h5 == state ? _GEN_9722 : ram_0_91; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10754 = 3'h5 == state ? _GEN_9723 : ram_0_92; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10755 = 3'h5 == state ? _GEN_9724 : ram_0_93; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10756 = 3'h5 == state ? _GEN_9725 : ram_0_94; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10757 = 3'h5 == state ? _GEN_9726 : ram_0_95; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10758 = 3'h5 == state ? _GEN_9727 : ram_0_96; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10759 = 3'h5 == state ? _GEN_9728 : ram_0_97; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10760 = 3'h5 == state ? _GEN_9729 : ram_0_98; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10761 = 3'h5 == state ? _GEN_9730 : ram_0_99; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10762 = 3'h5 == state ? _GEN_9731 : ram_0_100; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10763 = 3'h5 == state ? _GEN_9732 : ram_0_101; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10764 = 3'h5 == state ? _GEN_9733 : ram_0_102; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10765 = 3'h5 == state ? _GEN_9734 : ram_0_103; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10766 = 3'h5 == state ? _GEN_9735 : ram_0_104; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10767 = 3'h5 == state ? _GEN_9736 : ram_0_105; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10768 = 3'h5 == state ? _GEN_9737 : ram_0_106; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10769 = 3'h5 == state ? _GEN_9738 : ram_0_107; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10770 = 3'h5 == state ? _GEN_9739 : ram_0_108; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10771 = 3'h5 == state ? _GEN_9740 : ram_0_109; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10772 = 3'h5 == state ? _GEN_9741 : ram_0_110; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10773 = 3'h5 == state ? _GEN_9742 : ram_0_111; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10774 = 3'h5 == state ? _GEN_9743 : ram_0_112; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10775 = 3'h5 == state ? _GEN_9744 : ram_0_113; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10776 = 3'h5 == state ? _GEN_9745 : ram_0_114; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10777 = 3'h5 == state ? _GEN_9746 : ram_0_115; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10778 = 3'h5 == state ? _GEN_9747 : ram_0_116; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10779 = 3'h5 == state ? _GEN_9748 : ram_0_117; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10780 = 3'h5 == state ? _GEN_9749 : ram_0_118; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10781 = 3'h5 == state ? _GEN_9750 : ram_0_119; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10782 = 3'h5 == state ? _GEN_9751 : ram_0_120; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10783 = 3'h5 == state ? _GEN_9752 : ram_0_121; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10784 = 3'h5 == state ? _GEN_9753 : ram_0_122; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10785 = 3'h5 == state ? _GEN_9754 : ram_0_123; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10786 = 3'h5 == state ? _GEN_9755 : ram_0_124; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10787 = 3'h5 == state ? _GEN_9756 : ram_0_125; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10788 = 3'h5 == state ? _GEN_9757 : ram_0_126; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_10789 = 3'h5 == state ? _GEN_9758 : ram_0_127; // @[d_cache.scala 81:18 18:24]
  wire [31:0] _GEN_10790 = 3'h5 == state ? _GEN_9759 : tag_0_0; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10791 = 3'h5 == state ? _GEN_9760 : tag_0_1; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10792 = 3'h5 == state ? _GEN_9761 : tag_0_2; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10793 = 3'h5 == state ? _GEN_9762 : tag_0_3; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10794 = 3'h5 == state ? _GEN_9763 : tag_0_4; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10795 = 3'h5 == state ? _GEN_9764 : tag_0_5; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10796 = 3'h5 == state ? _GEN_9765 : tag_0_6; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10797 = 3'h5 == state ? _GEN_9766 : tag_0_7; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10798 = 3'h5 == state ? _GEN_9767 : tag_0_8; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10799 = 3'h5 == state ? _GEN_9768 : tag_0_9; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10800 = 3'h5 == state ? _GEN_9769 : tag_0_10; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10801 = 3'h5 == state ? _GEN_9770 : tag_0_11; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10802 = 3'h5 == state ? _GEN_9771 : tag_0_12; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10803 = 3'h5 == state ? _GEN_9772 : tag_0_13; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10804 = 3'h5 == state ? _GEN_9773 : tag_0_14; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10805 = 3'h5 == state ? _GEN_9774 : tag_0_15; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10806 = 3'h5 == state ? _GEN_9775 : tag_0_16; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10807 = 3'h5 == state ? _GEN_9776 : tag_0_17; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10808 = 3'h5 == state ? _GEN_9777 : tag_0_18; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10809 = 3'h5 == state ? _GEN_9778 : tag_0_19; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10810 = 3'h5 == state ? _GEN_9779 : tag_0_20; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10811 = 3'h5 == state ? _GEN_9780 : tag_0_21; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10812 = 3'h5 == state ? _GEN_9781 : tag_0_22; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10813 = 3'h5 == state ? _GEN_9782 : tag_0_23; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10814 = 3'h5 == state ? _GEN_9783 : tag_0_24; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10815 = 3'h5 == state ? _GEN_9784 : tag_0_25; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10816 = 3'h5 == state ? _GEN_9785 : tag_0_26; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10817 = 3'h5 == state ? _GEN_9786 : tag_0_27; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10818 = 3'h5 == state ? _GEN_9787 : tag_0_28; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10819 = 3'h5 == state ? _GEN_9788 : tag_0_29; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10820 = 3'h5 == state ? _GEN_9789 : tag_0_30; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10821 = 3'h5 == state ? _GEN_9790 : tag_0_31; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10822 = 3'h5 == state ? _GEN_9791 : tag_0_32; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10823 = 3'h5 == state ? _GEN_9792 : tag_0_33; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10824 = 3'h5 == state ? _GEN_9793 : tag_0_34; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10825 = 3'h5 == state ? _GEN_9794 : tag_0_35; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10826 = 3'h5 == state ? _GEN_9795 : tag_0_36; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10827 = 3'h5 == state ? _GEN_9796 : tag_0_37; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10828 = 3'h5 == state ? _GEN_9797 : tag_0_38; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10829 = 3'h5 == state ? _GEN_9798 : tag_0_39; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10830 = 3'h5 == state ? _GEN_9799 : tag_0_40; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10831 = 3'h5 == state ? _GEN_9800 : tag_0_41; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10832 = 3'h5 == state ? _GEN_9801 : tag_0_42; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10833 = 3'h5 == state ? _GEN_9802 : tag_0_43; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10834 = 3'h5 == state ? _GEN_9803 : tag_0_44; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10835 = 3'h5 == state ? _GEN_9804 : tag_0_45; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10836 = 3'h5 == state ? _GEN_9805 : tag_0_46; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10837 = 3'h5 == state ? _GEN_9806 : tag_0_47; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10838 = 3'h5 == state ? _GEN_9807 : tag_0_48; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10839 = 3'h5 == state ? _GEN_9808 : tag_0_49; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10840 = 3'h5 == state ? _GEN_9809 : tag_0_50; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10841 = 3'h5 == state ? _GEN_9810 : tag_0_51; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10842 = 3'h5 == state ? _GEN_9811 : tag_0_52; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10843 = 3'h5 == state ? _GEN_9812 : tag_0_53; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10844 = 3'h5 == state ? _GEN_9813 : tag_0_54; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10845 = 3'h5 == state ? _GEN_9814 : tag_0_55; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10846 = 3'h5 == state ? _GEN_9815 : tag_0_56; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10847 = 3'h5 == state ? _GEN_9816 : tag_0_57; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10848 = 3'h5 == state ? _GEN_9817 : tag_0_58; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10849 = 3'h5 == state ? _GEN_9818 : tag_0_59; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10850 = 3'h5 == state ? _GEN_9819 : tag_0_60; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10851 = 3'h5 == state ? _GEN_9820 : tag_0_61; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10852 = 3'h5 == state ? _GEN_9821 : tag_0_62; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10853 = 3'h5 == state ? _GEN_9822 : tag_0_63; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10854 = 3'h5 == state ? _GEN_9823 : tag_0_64; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10855 = 3'h5 == state ? _GEN_9824 : tag_0_65; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10856 = 3'h5 == state ? _GEN_9825 : tag_0_66; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10857 = 3'h5 == state ? _GEN_9826 : tag_0_67; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10858 = 3'h5 == state ? _GEN_9827 : tag_0_68; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10859 = 3'h5 == state ? _GEN_9828 : tag_0_69; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10860 = 3'h5 == state ? _GEN_9829 : tag_0_70; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10861 = 3'h5 == state ? _GEN_9830 : tag_0_71; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10862 = 3'h5 == state ? _GEN_9831 : tag_0_72; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10863 = 3'h5 == state ? _GEN_9832 : tag_0_73; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10864 = 3'h5 == state ? _GEN_9833 : tag_0_74; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10865 = 3'h5 == state ? _GEN_9834 : tag_0_75; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10866 = 3'h5 == state ? _GEN_9835 : tag_0_76; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10867 = 3'h5 == state ? _GEN_9836 : tag_0_77; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10868 = 3'h5 == state ? _GEN_9837 : tag_0_78; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10869 = 3'h5 == state ? _GEN_9838 : tag_0_79; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10870 = 3'h5 == state ? _GEN_9839 : tag_0_80; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10871 = 3'h5 == state ? _GEN_9840 : tag_0_81; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10872 = 3'h5 == state ? _GEN_9841 : tag_0_82; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10873 = 3'h5 == state ? _GEN_9842 : tag_0_83; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10874 = 3'h5 == state ? _GEN_9843 : tag_0_84; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10875 = 3'h5 == state ? _GEN_9844 : tag_0_85; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10876 = 3'h5 == state ? _GEN_9845 : tag_0_86; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10877 = 3'h5 == state ? _GEN_9846 : tag_0_87; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10878 = 3'h5 == state ? _GEN_9847 : tag_0_88; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10879 = 3'h5 == state ? _GEN_9848 : tag_0_89; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10880 = 3'h5 == state ? _GEN_9849 : tag_0_90; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10881 = 3'h5 == state ? _GEN_9850 : tag_0_91; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10882 = 3'h5 == state ? _GEN_9851 : tag_0_92; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10883 = 3'h5 == state ? _GEN_9852 : tag_0_93; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10884 = 3'h5 == state ? _GEN_9853 : tag_0_94; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10885 = 3'h5 == state ? _GEN_9854 : tag_0_95; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10886 = 3'h5 == state ? _GEN_9855 : tag_0_96; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10887 = 3'h5 == state ? _GEN_9856 : tag_0_97; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10888 = 3'h5 == state ? _GEN_9857 : tag_0_98; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10889 = 3'h5 == state ? _GEN_9858 : tag_0_99; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10890 = 3'h5 == state ? _GEN_9859 : tag_0_100; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10891 = 3'h5 == state ? _GEN_9860 : tag_0_101; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10892 = 3'h5 == state ? _GEN_9861 : tag_0_102; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10893 = 3'h5 == state ? _GEN_9862 : tag_0_103; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10894 = 3'h5 == state ? _GEN_9863 : tag_0_104; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10895 = 3'h5 == state ? _GEN_9864 : tag_0_105; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10896 = 3'h5 == state ? _GEN_9865 : tag_0_106; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10897 = 3'h5 == state ? _GEN_9866 : tag_0_107; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10898 = 3'h5 == state ? _GEN_9867 : tag_0_108; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10899 = 3'h5 == state ? _GEN_9868 : tag_0_109; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10900 = 3'h5 == state ? _GEN_9869 : tag_0_110; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10901 = 3'h5 == state ? _GEN_9870 : tag_0_111; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10902 = 3'h5 == state ? _GEN_9871 : tag_0_112; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10903 = 3'h5 == state ? _GEN_9872 : tag_0_113; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10904 = 3'h5 == state ? _GEN_9873 : tag_0_114; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10905 = 3'h5 == state ? _GEN_9874 : tag_0_115; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10906 = 3'h5 == state ? _GEN_9875 : tag_0_116; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10907 = 3'h5 == state ? _GEN_9876 : tag_0_117; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10908 = 3'h5 == state ? _GEN_9877 : tag_0_118; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10909 = 3'h5 == state ? _GEN_9878 : tag_0_119; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10910 = 3'h5 == state ? _GEN_9879 : tag_0_120; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10911 = 3'h5 == state ? _GEN_9880 : tag_0_121; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10912 = 3'h5 == state ? _GEN_9881 : tag_0_122; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10913 = 3'h5 == state ? _GEN_9882 : tag_0_123; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10914 = 3'h5 == state ? _GEN_9883 : tag_0_124; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10915 = 3'h5 == state ? _GEN_9884 : tag_0_125; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10916 = 3'h5 == state ? _GEN_9885 : tag_0_126; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_10917 = 3'h5 == state ? _GEN_9886 : tag_0_127; // @[d_cache.scala 81:18 22:24]
  wire  _GEN_10918 = 3'h5 == state ? _GEN_9887 : valid_0_0; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10919 = 3'h5 == state ? _GEN_9888 : valid_0_1; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10920 = 3'h5 == state ? _GEN_9889 : valid_0_2; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10921 = 3'h5 == state ? _GEN_9890 : valid_0_3; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10922 = 3'h5 == state ? _GEN_9891 : valid_0_4; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10923 = 3'h5 == state ? _GEN_9892 : valid_0_5; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10924 = 3'h5 == state ? _GEN_9893 : valid_0_6; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10925 = 3'h5 == state ? _GEN_9894 : valid_0_7; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10926 = 3'h5 == state ? _GEN_9895 : valid_0_8; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10927 = 3'h5 == state ? _GEN_9896 : valid_0_9; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10928 = 3'h5 == state ? _GEN_9897 : valid_0_10; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10929 = 3'h5 == state ? _GEN_9898 : valid_0_11; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10930 = 3'h5 == state ? _GEN_9899 : valid_0_12; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10931 = 3'h5 == state ? _GEN_9900 : valid_0_13; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10932 = 3'h5 == state ? _GEN_9901 : valid_0_14; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10933 = 3'h5 == state ? _GEN_9902 : valid_0_15; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10934 = 3'h5 == state ? _GEN_9903 : valid_0_16; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10935 = 3'h5 == state ? _GEN_9904 : valid_0_17; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10936 = 3'h5 == state ? _GEN_9905 : valid_0_18; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10937 = 3'h5 == state ? _GEN_9906 : valid_0_19; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10938 = 3'h5 == state ? _GEN_9907 : valid_0_20; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10939 = 3'h5 == state ? _GEN_9908 : valid_0_21; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10940 = 3'h5 == state ? _GEN_9909 : valid_0_22; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10941 = 3'h5 == state ? _GEN_9910 : valid_0_23; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10942 = 3'h5 == state ? _GEN_9911 : valid_0_24; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10943 = 3'h5 == state ? _GEN_9912 : valid_0_25; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10944 = 3'h5 == state ? _GEN_9913 : valid_0_26; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10945 = 3'h5 == state ? _GEN_9914 : valid_0_27; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10946 = 3'h5 == state ? _GEN_9915 : valid_0_28; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10947 = 3'h5 == state ? _GEN_9916 : valid_0_29; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10948 = 3'h5 == state ? _GEN_9917 : valid_0_30; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10949 = 3'h5 == state ? _GEN_9918 : valid_0_31; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10950 = 3'h5 == state ? _GEN_9919 : valid_0_32; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10951 = 3'h5 == state ? _GEN_9920 : valid_0_33; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10952 = 3'h5 == state ? _GEN_9921 : valid_0_34; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10953 = 3'h5 == state ? _GEN_9922 : valid_0_35; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10954 = 3'h5 == state ? _GEN_9923 : valid_0_36; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10955 = 3'h5 == state ? _GEN_9924 : valid_0_37; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10956 = 3'h5 == state ? _GEN_9925 : valid_0_38; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10957 = 3'h5 == state ? _GEN_9926 : valid_0_39; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10958 = 3'h5 == state ? _GEN_9927 : valid_0_40; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10959 = 3'h5 == state ? _GEN_9928 : valid_0_41; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10960 = 3'h5 == state ? _GEN_9929 : valid_0_42; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10961 = 3'h5 == state ? _GEN_9930 : valid_0_43; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10962 = 3'h5 == state ? _GEN_9931 : valid_0_44; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10963 = 3'h5 == state ? _GEN_9932 : valid_0_45; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10964 = 3'h5 == state ? _GEN_9933 : valid_0_46; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10965 = 3'h5 == state ? _GEN_9934 : valid_0_47; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10966 = 3'h5 == state ? _GEN_9935 : valid_0_48; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10967 = 3'h5 == state ? _GEN_9936 : valid_0_49; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10968 = 3'h5 == state ? _GEN_9937 : valid_0_50; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10969 = 3'h5 == state ? _GEN_9938 : valid_0_51; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10970 = 3'h5 == state ? _GEN_9939 : valid_0_52; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10971 = 3'h5 == state ? _GEN_9940 : valid_0_53; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10972 = 3'h5 == state ? _GEN_9941 : valid_0_54; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10973 = 3'h5 == state ? _GEN_9942 : valid_0_55; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10974 = 3'h5 == state ? _GEN_9943 : valid_0_56; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10975 = 3'h5 == state ? _GEN_9944 : valid_0_57; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10976 = 3'h5 == state ? _GEN_9945 : valid_0_58; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10977 = 3'h5 == state ? _GEN_9946 : valid_0_59; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10978 = 3'h5 == state ? _GEN_9947 : valid_0_60; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10979 = 3'h5 == state ? _GEN_9948 : valid_0_61; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10980 = 3'h5 == state ? _GEN_9949 : valid_0_62; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10981 = 3'h5 == state ? _GEN_9950 : valid_0_63; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10982 = 3'h5 == state ? _GEN_9951 : valid_0_64; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10983 = 3'h5 == state ? _GEN_9952 : valid_0_65; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10984 = 3'h5 == state ? _GEN_9953 : valid_0_66; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10985 = 3'h5 == state ? _GEN_9954 : valid_0_67; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10986 = 3'h5 == state ? _GEN_9955 : valid_0_68; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10987 = 3'h5 == state ? _GEN_9956 : valid_0_69; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10988 = 3'h5 == state ? _GEN_9957 : valid_0_70; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10989 = 3'h5 == state ? _GEN_9958 : valid_0_71; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10990 = 3'h5 == state ? _GEN_9959 : valid_0_72; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10991 = 3'h5 == state ? _GEN_9960 : valid_0_73; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10992 = 3'h5 == state ? _GEN_9961 : valid_0_74; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10993 = 3'h5 == state ? _GEN_9962 : valid_0_75; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10994 = 3'h5 == state ? _GEN_9963 : valid_0_76; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10995 = 3'h5 == state ? _GEN_9964 : valid_0_77; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10996 = 3'h5 == state ? _GEN_9965 : valid_0_78; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10997 = 3'h5 == state ? _GEN_9966 : valid_0_79; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10998 = 3'h5 == state ? _GEN_9967 : valid_0_80; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_10999 = 3'h5 == state ? _GEN_9968 : valid_0_81; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11000 = 3'h5 == state ? _GEN_9969 : valid_0_82; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11001 = 3'h5 == state ? _GEN_9970 : valid_0_83; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11002 = 3'h5 == state ? _GEN_9971 : valid_0_84; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11003 = 3'h5 == state ? _GEN_9972 : valid_0_85; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11004 = 3'h5 == state ? _GEN_9973 : valid_0_86; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11005 = 3'h5 == state ? _GEN_9974 : valid_0_87; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11006 = 3'h5 == state ? _GEN_9975 : valid_0_88; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11007 = 3'h5 == state ? _GEN_9976 : valid_0_89; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11008 = 3'h5 == state ? _GEN_9977 : valid_0_90; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11009 = 3'h5 == state ? _GEN_9978 : valid_0_91; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11010 = 3'h5 == state ? _GEN_9979 : valid_0_92; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11011 = 3'h5 == state ? _GEN_9980 : valid_0_93; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11012 = 3'h5 == state ? _GEN_9981 : valid_0_94; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11013 = 3'h5 == state ? _GEN_9982 : valid_0_95; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11014 = 3'h5 == state ? _GEN_9983 : valid_0_96; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11015 = 3'h5 == state ? _GEN_9984 : valid_0_97; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11016 = 3'h5 == state ? _GEN_9985 : valid_0_98; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11017 = 3'h5 == state ? _GEN_9986 : valid_0_99; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11018 = 3'h5 == state ? _GEN_9987 : valid_0_100; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11019 = 3'h5 == state ? _GEN_9988 : valid_0_101; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11020 = 3'h5 == state ? _GEN_9989 : valid_0_102; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11021 = 3'h5 == state ? _GEN_9990 : valid_0_103; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11022 = 3'h5 == state ? _GEN_9991 : valid_0_104; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11023 = 3'h5 == state ? _GEN_9992 : valid_0_105; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11024 = 3'h5 == state ? _GEN_9993 : valid_0_106; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11025 = 3'h5 == state ? _GEN_9994 : valid_0_107; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11026 = 3'h5 == state ? _GEN_9995 : valid_0_108; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11027 = 3'h5 == state ? _GEN_9996 : valid_0_109; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11028 = 3'h5 == state ? _GEN_9997 : valid_0_110; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11029 = 3'h5 == state ? _GEN_9998 : valid_0_111; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11030 = 3'h5 == state ? _GEN_9999 : valid_0_112; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11031 = 3'h5 == state ? _GEN_10000 : valid_0_113; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11032 = 3'h5 == state ? _GEN_10001 : valid_0_114; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11033 = 3'h5 == state ? _GEN_10002 : valid_0_115; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11034 = 3'h5 == state ? _GEN_10003 : valid_0_116; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11035 = 3'h5 == state ? _GEN_10004 : valid_0_117; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11036 = 3'h5 == state ? _GEN_10005 : valid_0_118; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11037 = 3'h5 == state ? _GEN_10006 : valid_0_119; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11038 = 3'h5 == state ? _GEN_10007 : valid_0_120; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11039 = 3'h5 == state ? _GEN_10008 : valid_0_121; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11040 = 3'h5 == state ? _GEN_10009 : valid_0_122; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11041 = 3'h5 == state ? _GEN_10010 : valid_0_123; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11042 = 3'h5 == state ? _GEN_10011 : valid_0_124; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11043 = 3'h5 == state ? _GEN_10012 : valid_0_125; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11044 = 3'h5 == state ? _GEN_10013 : valid_0_126; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11045 = 3'h5 == state ? _GEN_10014 : valid_0_127; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11046 = 3'h5 == state ? _GEN_10015 : quene; // @[d_cache.scala 81:18 37:24]
  wire [63:0] _GEN_11047 = 3'h5 == state ? _GEN_10016 : ram_1_0; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11048 = 3'h5 == state ? _GEN_10017 : ram_1_1; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11049 = 3'h5 == state ? _GEN_10018 : ram_1_2; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11050 = 3'h5 == state ? _GEN_10019 : ram_1_3; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11051 = 3'h5 == state ? _GEN_10020 : ram_1_4; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11052 = 3'h5 == state ? _GEN_10021 : ram_1_5; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11053 = 3'h5 == state ? _GEN_10022 : ram_1_6; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11054 = 3'h5 == state ? _GEN_10023 : ram_1_7; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11055 = 3'h5 == state ? _GEN_10024 : ram_1_8; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11056 = 3'h5 == state ? _GEN_10025 : ram_1_9; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11057 = 3'h5 == state ? _GEN_10026 : ram_1_10; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11058 = 3'h5 == state ? _GEN_10027 : ram_1_11; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11059 = 3'h5 == state ? _GEN_10028 : ram_1_12; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11060 = 3'h5 == state ? _GEN_10029 : ram_1_13; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11061 = 3'h5 == state ? _GEN_10030 : ram_1_14; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11062 = 3'h5 == state ? _GEN_10031 : ram_1_15; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11063 = 3'h5 == state ? _GEN_10032 : ram_1_16; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11064 = 3'h5 == state ? _GEN_10033 : ram_1_17; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11065 = 3'h5 == state ? _GEN_10034 : ram_1_18; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11066 = 3'h5 == state ? _GEN_10035 : ram_1_19; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11067 = 3'h5 == state ? _GEN_10036 : ram_1_20; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11068 = 3'h5 == state ? _GEN_10037 : ram_1_21; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11069 = 3'h5 == state ? _GEN_10038 : ram_1_22; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11070 = 3'h5 == state ? _GEN_10039 : ram_1_23; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11071 = 3'h5 == state ? _GEN_10040 : ram_1_24; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11072 = 3'h5 == state ? _GEN_10041 : ram_1_25; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11073 = 3'h5 == state ? _GEN_10042 : ram_1_26; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11074 = 3'h5 == state ? _GEN_10043 : ram_1_27; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11075 = 3'h5 == state ? _GEN_10044 : ram_1_28; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11076 = 3'h5 == state ? _GEN_10045 : ram_1_29; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11077 = 3'h5 == state ? _GEN_10046 : ram_1_30; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11078 = 3'h5 == state ? _GEN_10047 : ram_1_31; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11079 = 3'h5 == state ? _GEN_10048 : ram_1_32; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11080 = 3'h5 == state ? _GEN_10049 : ram_1_33; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11081 = 3'h5 == state ? _GEN_10050 : ram_1_34; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11082 = 3'h5 == state ? _GEN_10051 : ram_1_35; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11083 = 3'h5 == state ? _GEN_10052 : ram_1_36; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11084 = 3'h5 == state ? _GEN_10053 : ram_1_37; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11085 = 3'h5 == state ? _GEN_10054 : ram_1_38; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11086 = 3'h5 == state ? _GEN_10055 : ram_1_39; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11087 = 3'h5 == state ? _GEN_10056 : ram_1_40; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11088 = 3'h5 == state ? _GEN_10057 : ram_1_41; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11089 = 3'h5 == state ? _GEN_10058 : ram_1_42; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11090 = 3'h5 == state ? _GEN_10059 : ram_1_43; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11091 = 3'h5 == state ? _GEN_10060 : ram_1_44; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11092 = 3'h5 == state ? _GEN_10061 : ram_1_45; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11093 = 3'h5 == state ? _GEN_10062 : ram_1_46; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11094 = 3'h5 == state ? _GEN_10063 : ram_1_47; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11095 = 3'h5 == state ? _GEN_10064 : ram_1_48; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11096 = 3'h5 == state ? _GEN_10065 : ram_1_49; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11097 = 3'h5 == state ? _GEN_10066 : ram_1_50; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11098 = 3'h5 == state ? _GEN_10067 : ram_1_51; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11099 = 3'h5 == state ? _GEN_10068 : ram_1_52; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11100 = 3'h5 == state ? _GEN_10069 : ram_1_53; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11101 = 3'h5 == state ? _GEN_10070 : ram_1_54; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11102 = 3'h5 == state ? _GEN_10071 : ram_1_55; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11103 = 3'h5 == state ? _GEN_10072 : ram_1_56; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11104 = 3'h5 == state ? _GEN_10073 : ram_1_57; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11105 = 3'h5 == state ? _GEN_10074 : ram_1_58; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11106 = 3'h5 == state ? _GEN_10075 : ram_1_59; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11107 = 3'h5 == state ? _GEN_10076 : ram_1_60; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11108 = 3'h5 == state ? _GEN_10077 : ram_1_61; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11109 = 3'h5 == state ? _GEN_10078 : ram_1_62; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11110 = 3'h5 == state ? _GEN_10079 : ram_1_63; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11111 = 3'h5 == state ? _GEN_10080 : ram_1_64; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11112 = 3'h5 == state ? _GEN_10081 : ram_1_65; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11113 = 3'h5 == state ? _GEN_10082 : ram_1_66; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11114 = 3'h5 == state ? _GEN_10083 : ram_1_67; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11115 = 3'h5 == state ? _GEN_10084 : ram_1_68; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11116 = 3'h5 == state ? _GEN_10085 : ram_1_69; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11117 = 3'h5 == state ? _GEN_10086 : ram_1_70; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11118 = 3'h5 == state ? _GEN_10087 : ram_1_71; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11119 = 3'h5 == state ? _GEN_10088 : ram_1_72; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11120 = 3'h5 == state ? _GEN_10089 : ram_1_73; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11121 = 3'h5 == state ? _GEN_10090 : ram_1_74; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11122 = 3'h5 == state ? _GEN_10091 : ram_1_75; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11123 = 3'h5 == state ? _GEN_10092 : ram_1_76; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11124 = 3'h5 == state ? _GEN_10093 : ram_1_77; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11125 = 3'h5 == state ? _GEN_10094 : ram_1_78; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11126 = 3'h5 == state ? _GEN_10095 : ram_1_79; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11127 = 3'h5 == state ? _GEN_10096 : ram_1_80; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11128 = 3'h5 == state ? _GEN_10097 : ram_1_81; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11129 = 3'h5 == state ? _GEN_10098 : ram_1_82; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11130 = 3'h5 == state ? _GEN_10099 : ram_1_83; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11131 = 3'h5 == state ? _GEN_10100 : ram_1_84; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11132 = 3'h5 == state ? _GEN_10101 : ram_1_85; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11133 = 3'h5 == state ? _GEN_10102 : ram_1_86; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11134 = 3'h5 == state ? _GEN_10103 : ram_1_87; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11135 = 3'h5 == state ? _GEN_10104 : ram_1_88; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11136 = 3'h5 == state ? _GEN_10105 : ram_1_89; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11137 = 3'h5 == state ? _GEN_10106 : ram_1_90; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11138 = 3'h5 == state ? _GEN_10107 : ram_1_91; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11139 = 3'h5 == state ? _GEN_10108 : ram_1_92; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11140 = 3'h5 == state ? _GEN_10109 : ram_1_93; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11141 = 3'h5 == state ? _GEN_10110 : ram_1_94; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11142 = 3'h5 == state ? _GEN_10111 : ram_1_95; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11143 = 3'h5 == state ? _GEN_10112 : ram_1_96; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11144 = 3'h5 == state ? _GEN_10113 : ram_1_97; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11145 = 3'h5 == state ? _GEN_10114 : ram_1_98; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11146 = 3'h5 == state ? _GEN_10115 : ram_1_99; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11147 = 3'h5 == state ? _GEN_10116 : ram_1_100; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11148 = 3'h5 == state ? _GEN_10117 : ram_1_101; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11149 = 3'h5 == state ? _GEN_10118 : ram_1_102; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11150 = 3'h5 == state ? _GEN_10119 : ram_1_103; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11151 = 3'h5 == state ? _GEN_10120 : ram_1_104; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11152 = 3'h5 == state ? _GEN_10121 : ram_1_105; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11153 = 3'h5 == state ? _GEN_10122 : ram_1_106; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11154 = 3'h5 == state ? _GEN_10123 : ram_1_107; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11155 = 3'h5 == state ? _GEN_10124 : ram_1_108; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11156 = 3'h5 == state ? _GEN_10125 : ram_1_109; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11157 = 3'h5 == state ? _GEN_10126 : ram_1_110; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11158 = 3'h5 == state ? _GEN_10127 : ram_1_111; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11159 = 3'h5 == state ? _GEN_10128 : ram_1_112; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11160 = 3'h5 == state ? _GEN_10129 : ram_1_113; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11161 = 3'h5 == state ? _GEN_10130 : ram_1_114; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11162 = 3'h5 == state ? _GEN_10131 : ram_1_115; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11163 = 3'h5 == state ? _GEN_10132 : ram_1_116; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11164 = 3'h5 == state ? _GEN_10133 : ram_1_117; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11165 = 3'h5 == state ? _GEN_10134 : ram_1_118; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11166 = 3'h5 == state ? _GEN_10135 : ram_1_119; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11167 = 3'h5 == state ? _GEN_10136 : ram_1_120; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11168 = 3'h5 == state ? _GEN_10137 : ram_1_121; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11169 = 3'h5 == state ? _GEN_10138 : ram_1_122; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11170 = 3'h5 == state ? _GEN_10139 : ram_1_123; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11171 = 3'h5 == state ? _GEN_10140 : ram_1_124; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11172 = 3'h5 == state ? _GEN_10141 : ram_1_125; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11173 = 3'h5 == state ? _GEN_10142 : ram_1_126; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_11174 = 3'h5 == state ? _GEN_10143 : ram_1_127; // @[d_cache.scala 81:18 19:24]
  wire [31:0] _GEN_11175 = 3'h5 == state ? _GEN_10144 : tag_1_0; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11176 = 3'h5 == state ? _GEN_10145 : tag_1_1; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11177 = 3'h5 == state ? _GEN_10146 : tag_1_2; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11178 = 3'h5 == state ? _GEN_10147 : tag_1_3; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11179 = 3'h5 == state ? _GEN_10148 : tag_1_4; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11180 = 3'h5 == state ? _GEN_10149 : tag_1_5; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11181 = 3'h5 == state ? _GEN_10150 : tag_1_6; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11182 = 3'h5 == state ? _GEN_10151 : tag_1_7; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11183 = 3'h5 == state ? _GEN_10152 : tag_1_8; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11184 = 3'h5 == state ? _GEN_10153 : tag_1_9; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11185 = 3'h5 == state ? _GEN_10154 : tag_1_10; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11186 = 3'h5 == state ? _GEN_10155 : tag_1_11; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11187 = 3'h5 == state ? _GEN_10156 : tag_1_12; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11188 = 3'h5 == state ? _GEN_10157 : tag_1_13; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11189 = 3'h5 == state ? _GEN_10158 : tag_1_14; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11190 = 3'h5 == state ? _GEN_10159 : tag_1_15; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11191 = 3'h5 == state ? _GEN_10160 : tag_1_16; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11192 = 3'h5 == state ? _GEN_10161 : tag_1_17; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11193 = 3'h5 == state ? _GEN_10162 : tag_1_18; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11194 = 3'h5 == state ? _GEN_10163 : tag_1_19; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11195 = 3'h5 == state ? _GEN_10164 : tag_1_20; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11196 = 3'h5 == state ? _GEN_10165 : tag_1_21; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11197 = 3'h5 == state ? _GEN_10166 : tag_1_22; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11198 = 3'h5 == state ? _GEN_10167 : tag_1_23; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11199 = 3'h5 == state ? _GEN_10168 : tag_1_24; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11200 = 3'h5 == state ? _GEN_10169 : tag_1_25; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11201 = 3'h5 == state ? _GEN_10170 : tag_1_26; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11202 = 3'h5 == state ? _GEN_10171 : tag_1_27; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11203 = 3'h5 == state ? _GEN_10172 : tag_1_28; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11204 = 3'h5 == state ? _GEN_10173 : tag_1_29; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11205 = 3'h5 == state ? _GEN_10174 : tag_1_30; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11206 = 3'h5 == state ? _GEN_10175 : tag_1_31; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11207 = 3'h5 == state ? _GEN_10176 : tag_1_32; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11208 = 3'h5 == state ? _GEN_10177 : tag_1_33; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11209 = 3'h5 == state ? _GEN_10178 : tag_1_34; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11210 = 3'h5 == state ? _GEN_10179 : tag_1_35; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11211 = 3'h5 == state ? _GEN_10180 : tag_1_36; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11212 = 3'h5 == state ? _GEN_10181 : tag_1_37; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11213 = 3'h5 == state ? _GEN_10182 : tag_1_38; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11214 = 3'h5 == state ? _GEN_10183 : tag_1_39; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11215 = 3'h5 == state ? _GEN_10184 : tag_1_40; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11216 = 3'h5 == state ? _GEN_10185 : tag_1_41; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11217 = 3'h5 == state ? _GEN_10186 : tag_1_42; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11218 = 3'h5 == state ? _GEN_10187 : tag_1_43; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11219 = 3'h5 == state ? _GEN_10188 : tag_1_44; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11220 = 3'h5 == state ? _GEN_10189 : tag_1_45; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11221 = 3'h5 == state ? _GEN_10190 : tag_1_46; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11222 = 3'h5 == state ? _GEN_10191 : tag_1_47; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11223 = 3'h5 == state ? _GEN_10192 : tag_1_48; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11224 = 3'h5 == state ? _GEN_10193 : tag_1_49; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11225 = 3'h5 == state ? _GEN_10194 : tag_1_50; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11226 = 3'h5 == state ? _GEN_10195 : tag_1_51; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11227 = 3'h5 == state ? _GEN_10196 : tag_1_52; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11228 = 3'h5 == state ? _GEN_10197 : tag_1_53; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11229 = 3'h5 == state ? _GEN_10198 : tag_1_54; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11230 = 3'h5 == state ? _GEN_10199 : tag_1_55; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11231 = 3'h5 == state ? _GEN_10200 : tag_1_56; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11232 = 3'h5 == state ? _GEN_10201 : tag_1_57; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11233 = 3'h5 == state ? _GEN_10202 : tag_1_58; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11234 = 3'h5 == state ? _GEN_10203 : tag_1_59; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11235 = 3'h5 == state ? _GEN_10204 : tag_1_60; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11236 = 3'h5 == state ? _GEN_10205 : tag_1_61; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11237 = 3'h5 == state ? _GEN_10206 : tag_1_62; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11238 = 3'h5 == state ? _GEN_10207 : tag_1_63; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11239 = 3'h5 == state ? _GEN_10208 : tag_1_64; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11240 = 3'h5 == state ? _GEN_10209 : tag_1_65; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11241 = 3'h5 == state ? _GEN_10210 : tag_1_66; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11242 = 3'h5 == state ? _GEN_10211 : tag_1_67; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11243 = 3'h5 == state ? _GEN_10212 : tag_1_68; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11244 = 3'h5 == state ? _GEN_10213 : tag_1_69; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11245 = 3'h5 == state ? _GEN_10214 : tag_1_70; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11246 = 3'h5 == state ? _GEN_10215 : tag_1_71; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11247 = 3'h5 == state ? _GEN_10216 : tag_1_72; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11248 = 3'h5 == state ? _GEN_10217 : tag_1_73; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11249 = 3'h5 == state ? _GEN_10218 : tag_1_74; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11250 = 3'h5 == state ? _GEN_10219 : tag_1_75; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11251 = 3'h5 == state ? _GEN_10220 : tag_1_76; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11252 = 3'h5 == state ? _GEN_10221 : tag_1_77; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11253 = 3'h5 == state ? _GEN_10222 : tag_1_78; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11254 = 3'h5 == state ? _GEN_10223 : tag_1_79; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11255 = 3'h5 == state ? _GEN_10224 : tag_1_80; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11256 = 3'h5 == state ? _GEN_10225 : tag_1_81; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11257 = 3'h5 == state ? _GEN_10226 : tag_1_82; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11258 = 3'h5 == state ? _GEN_10227 : tag_1_83; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11259 = 3'h5 == state ? _GEN_10228 : tag_1_84; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11260 = 3'h5 == state ? _GEN_10229 : tag_1_85; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11261 = 3'h5 == state ? _GEN_10230 : tag_1_86; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11262 = 3'h5 == state ? _GEN_10231 : tag_1_87; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11263 = 3'h5 == state ? _GEN_10232 : tag_1_88; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11264 = 3'h5 == state ? _GEN_10233 : tag_1_89; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11265 = 3'h5 == state ? _GEN_10234 : tag_1_90; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11266 = 3'h5 == state ? _GEN_10235 : tag_1_91; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11267 = 3'h5 == state ? _GEN_10236 : tag_1_92; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11268 = 3'h5 == state ? _GEN_10237 : tag_1_93; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11269 = 3'h5 == state ? _GEN_10238 : tag_1_94; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11270 = 3'h5 == state ? _GEN_10239 : tag_1_95; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11271 = 3'h5 == state ? _GEN_10240 : tag_1_96; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11272 = 3'h5 == state ? _GEN_10241 : tag_1_97; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11273 = 3'h5 == state ? _GEN_10242 : tag_1_98; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11274 = 3'h5 == state ? _GEN_10243 : tag_1_99; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11275 = 3'h5 == state ? _GEN_10244 : tag_1_100; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11276 = 3'h5 == state ? _GEN_10245 : tag_1_101; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11277 = 3'h5 == state ? _GEN_10246 : tag_1_102; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11278 = 3'h5 == state ? _GEN_10247 : tag_1_103; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11279 = 3'h5 == state ? _GEN_10248 : tag_1_104; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11280 = 3'h5 == state ? _GEN_10249 : tag_1_105; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11281 = 3'h5 == state ? _GEN_10250 : tag_1_106; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11282 = 3'h5 == state ? _GEN_10251 : tag_1_107; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11283 = 3'h5 == state ? _GEN_10252 : tag_1_108; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11284 = 3'h5 == state ? _GEN_10253 : tag_1_109; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11285 = 3'h5 == state ? _GEN_10254 : tag_1_110; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11286 = 3'h5 == state ? _GEN_10255 : tag_1_111; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11287 = 3'h5 == state ? _GEN_10256 : tag_1_112; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11288 = 3'h5 == state ? _GEN_10257 : tag_1_113; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11289 = 3'h5 == state ? _GEN_10258 : tag_1_114; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11290 = 3'h5 == state ? _GEN_10259 : tag_1_115; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11291 = 3'h5 == state ? _GEN_10260 : tag_1_116; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11292 = 3'h5 == state ? _GEN_10261 : tag_1_117; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11293 = 3'h5 == state ? _GEN_10262 : tag_1_118; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11294 = 3'h5 == state ? _GEN_10263 : tag_1_119; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11295 = 3'h5 == state ? _GEN_10264 : tag_1_120; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11296 = 3'h5 == state ? _GEN_10265 : tag_1_121; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11297 = 3'h5 == state ? _GEN_10266 : tag_1_122; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11298 = 3'h5 == state ? _GEN_10267 : tag_1_123; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11299 = 3'h5 == state ? _GEN_10268 : tag_1_124; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11300 = 3'h5 == state ? _GEN_10269 : tag_1_125; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11301 = 3'h5 == state ? _GEN_10270 : tag_1_126; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_11302 = 3'h5 == state ? _GEN_10271 : tag_1_127; // @[d_cache.scala 81:18 23:24]
  wire  _GEN_11303 = 3'h5 == state ? _GEN_10272 : valid_1_0; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11304 = 3'h5 == state ? _GEN_10273 : valid_1_1; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11305 = 3'h5 == state ? _GEN_10274 : valid_1_2; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11306 = 3'h5 == state ? _GEN_10275 : valid_1_3; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11307 = 3'h5 == state ? _GEN_10276 : valid_1_4; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11308 = 3'h5 == state ? _GEN_10277 : valid_1_5; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11309 = 3'h5 == state ? _GEN_10278 : valid_1_6; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11310 = 3'h5 == state ? _GEN_10279 : valid_1_7; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11311 = 3'h5 == state ? _GEN_10280 : valid_1_8; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11312 = 3'h5 == state ? _GEN_10281 : valid_1_9; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11313 = 3'h5 == state ? _GEN_10282 : valid_1_10; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11314 = 3'h5 == state ? _GEN_10283 : valid_1_11; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11315 = 3'h5 == state ? _GEN_10284 : valid_1_12; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11316 = 3'h5 == state ? _GEN_10285 : valid_1_13; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11317 = 3'h5 == state ? _GEN_10286 : valid_1_14; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11318 = 3'h5 == state ? _GEN_10287 : valid_1_15; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11319 = 3'h5 == state ? _GEN_10288 : valid_1_16; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11320 = 3'h5 == state ? _GEN_10289 : valid_1_17; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11321 = 3'h5 == state ? _GEN_10290 : valid_1_18; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11322 = 3'h5 == state ? _GEN_10291 : valid_1_19; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11323 = 3'h5 == state ? _GEN_10292 : valid_1_20; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11324 = 3'h5 == state ? _GEN_10293 : valid_1_21; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11325 = 3'h5 == state ? _GEN_10294 : valid_1_22; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11326 = 3'h5 == state ? _GEN_10295 : valid_1_23; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11327 = 3'h5 == state ? _GEN_10296 : valid_1_24; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11328 = 3'h5 == state ? _GEN_10297 : valid_1_25; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11329 = 3'h5 == state ? _GEN_10298 : valid_1_26; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11330 = 3'h5 == state ? _GEN_10299 : valid_1_27; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11331 = 3'h5 == state ? _GEN_10300 : valid_1_28; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11332 = 3'h5 == state ? _GEN_10301 : valid_1_29; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11333 = 3'h5 == state ? _GEN_10302 : valid_1_30; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11334 = 3'h5 == state ? _GEN_10303 : valid_1_31; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11335 = 3'h5 == state ? _GEN_10304 : valid_1_32; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11336 = 3'h5 == state ? _GEN_10305 : valid_1_33; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11337 = 3'h5 == state ? _GEN_10306 : valid_1_34; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11338 = 3'h5 == state ? _GEN_10307 : valid_1_35; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11339 = 3'h5 == state ? _GEN_10308 : valid_1_36; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11340 = 3'h5 == state ? _GEN_10309 : valid_1_37; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11341 = 3'h5 == state ? _GEN_10310 : valid_1_38; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11342 = 3'h5 == state ? _GEN_10311 : valid_1_39; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11343 = 3'h5 == state ? _GEN_10312 : valid_1_40; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11344 = 3'h5 == state ? _GEN_10313 : valid_1_41; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11345 = 3'h5 == state ? _GEN_10314 : valid_1_42; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11346 = 3'h5 == state ? _GEN_10315 : valid_1_43; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11347 = 3'h5 == state ? _GEN_10316 : valid_1_44; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11348 = 3'h5 == state ? _GEN_10317 : valid_1_45; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11349 = 3'h5 == state ? _GEN_10318 : valid_1_46; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11350 = 3'h5 == state ? _GEN_10319 : valid_1_47; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11351 = 3'h5 == state ? _GEN_10320 : valid_1_48; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11352 = 3'h5 == state ? _GEN_10321 : valid_1_49; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11353 = 3'h5 == state ? _GEN_10322 : valid_1_50; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11354 = 3'h5 == state ? _GEN_10323 : valid_1_51; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11355 = 3'h5 == state ? _GEN_10324 : valid_1_52; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11356 = 3'h5 == state ? _GEN_10325 : valid_1_53; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11357 = 3'h5 == state ? _GEN_10326 : valid_1_54; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11358 = 3'h5 == state ? _GEN_10327 : valid_1_55; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11359 = 3'h5 == state ? _GEN_10328 : valid_1_56; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11360 = 3'h5 == state ? _GEN_10329 : valid_1_57; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11361 = 3'h5 == state ? _GEN_10330 : valid_1_58; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11362 = 3'h5 == state ? _GEN_10331 : valid_1_59; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11363 = 3'h5 == state ? _GEN_10332 : valid_1_60; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11364 = 3'h5 == state ? _GEN_10333 : valid_1_61; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11365 = 3'h5 == state ? _GEN_10334 : valid_1_62; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11366 = 3'h5 == state ? _GEN_10335 : valid_1_63; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11367 = 3'h5 == state ? _GEN_10336 : valid_1_64; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11368 = 3'h5 == state ? _GEN_10337 : valid_1_65; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11369 = 3'h5 == state ? _GEN_10338 : valid_1_66; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11370 = 3'h5 == state ? _GEN_10339 : valid_1_67; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11371 = 3'h5 == state ? _GEN_10340 : valid_1_68; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11372 = 3'h5 == state ? _GEN_10341 : valid_1_69; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11373 = 3'h5 == state ? _GEN_10342 : valid_1_70; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11374 = 3'h5 == state ? _GEN_10343 : valid_1_71; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11375 = 3'h5 == state ? _GEN_10344 : valid_1_72; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11376 = 3'h5 == state ? _GEN_10345 : valid_1_73; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11377 = 3'h5 == state ? _GEN_10346 : valid_1_74; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11378 = 3'h5 == state ? _GEN_10347 : valid_1_75; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11379 = 3'h5 == state ? _GEN_10348 : valid_1_76; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11380 = 3'h5 == state ? _GEN_10349 : valid_1_77; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11381 = 3'h5 == state ? _GEN_10350 : valid_1_78; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11382 = 3'h5 == state ? _GEN_10351 : valid_1_79; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11383 = 3'h5 == state ? _GEN_10352 : valid_1_80; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11384 = 3'h5 == state ? _GEN_10353 : valid_1_81; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11385 = 3'h5 == state ? _GEN_10354 : valid_1_82; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11386 = 3'h5 == state ? _GEN_10355 : valid_1_83; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11387 = 3'h5 == state ? _GEN_10356 : valid_1_84; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11388 = 3'h5 == state ? _GEN_10357 : valid_1_85; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11389 = 3'h5 == state ? _GEN_10358 : valid_1_86; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11390 = 3'h5 == state ? _GEN_10359 : valid_1_87; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11391 = 3'h5 == state ? _GEN_10360 : valid_1_88; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11392 = 3'h5 == state ? _GEN_10361 : valid_1_89; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11393 = 3'h5 == state ? _GEN_10362 : valid_1_90; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11394 = 3'h5 == state ? _GEN_10363 : valid_1_91; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11395 = 3'h5 == state ? _GEN_10364 : valid_1_92; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11396 = 3'h5 == state ? _GEN_10365 : valid_1_93; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11397 = 3'h5 == state ? _GEN_10366 : valid_1_94; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11398 = 3'h5 == state ? _GEN_10367 : valid_1_95; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11399 = 3'h5 == state ? _GEN_10368 : valid_1_96; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11400 = 3'h5 == state ? _GEN_10369 : valid_1_97; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11401 = 3'h5 == state ? _GEN_10370 : valid_1_98; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11402 = 3'h5 == state ? _GEN_10371 : valid_1_99; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11403 = 3'h5 == state ? _GEN_10372 : valid_1_100; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11404 = 3'h5 == state ? _GEN_10373 : valid_1_101; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11405 = 3'h5 == state ? _GEN_10374 : valid_1_102; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11406 = 3'h5 == state ? _GEN_10375 : valid_1_103; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11407 = 3'h5 == state ? _GEN_10376 : valid_1_104; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11408 = 3'h5 == state ? _GEN_10377 : valid_1_105; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11409 = 3'h5 == state ? _GEN_10378 : valid_1_106; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11410 = 3'h5 == state ? _GEN_10379 : valid_1_107; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11411 = 3'h5 == state ? _GEN_10380 : valid_1_108; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11412 = 3'h5 == state ? _GEN_10381 : valid_1_109; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11413 = 3'h5 == state ? _GEN_10382 : valid_1_110; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11414 = 3'h5 == state ? _GEN_10383 : valid_1_111; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11415 = 3'h5 == state ? _GEN_10384 : valid_1_112; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11416 = 3'h5 == state ? _GEN_10385 : valid_1_113; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11417 = 3'h5 == state ? _GEN_10386 : valid_1_114; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11418 = 3'h5 == state ? _GEN_10387 : valid_1_115; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11419 = 3'h5 == state ? _GEN_10388 : valid_1_116; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11420 = 3'h5 == state ? _GEN_10389 : valid_1_117; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11421 = 3'h5 == state ? _GEN_10390 : valid_1_118; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11422 = 3'h5 == state ? _GEN_10391 : valid_1_119; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11423 = 3'h5 == state ? _GEN_10392 : valid_1_120; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11424 = 3'h5 == state ? _GEN_10393 : valid_1_121; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11425 = 3'h5 == state ? _GEN_10394 : valid_1_122; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11426 = 3'h5 == state ? _GEN_10395 : valid_1_123; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11427 = 3'h5 == state ? _GEN_10396 : valid_1_124; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11428 = 3'h5 == state ? _GEN_10397 : valid_1_125; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11429 = 3'h5 == state ? _GEN_10398 : valid_1_126; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_11430 = 3'h5 == state ? _GEN_10399 : valid_1_127; // @[d_cache.scala 81:18 25:26]
  wire [63:0] _GEN_11431 = 3'h5 == state ? _GEN_10400 : write_back_data; // @[d_cache.scala 81:18 31:34]
  wire [41:0] _GEN_11432 = 3'h5 == state ? _GEN_10401 : {{10'd0}, write_back_addr}; // @[d_cache.scala 81:18 32:34]
  wire  _GEN_11433 = 3'h5 == state ? _GEN_10402 : dirty_0_0; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11434 = 3'h5 == state ? _GEN_10403 : dirty_0_1; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11435 = 3'h5 == state ? _GEN_10404 : dirty_0_2; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11436 = 3'h5 == state ? _GEN_10405 : dirty_0_3; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11437 = 3'h5 == state ? _GEN_10406 : dirty_0_4; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11438 = 3'h5 == state ? _GEN_10407 : dirty_0_5; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11439 = 3'h5 == state ? _GEN_10408 : dirty_0_6; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11440 = 3'h5 == state ? _GEN_10409 : dirty_0_7; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11441 = 3'h5 == state ? _GEN_10410 : dirty_0_8; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11442 = 3'h5 == state ? _GEN_10411 : dirty_0_9; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11443 = 3'h5 == state ? _GEN_10412 : dirty_0_10; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11444 = 3'h5 == state ? _GEN_10413 : dirty_0_11; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11445 = 3'h5 == state ? _GEN_10414 : dirty_0_12; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11446 = 3'h5 == state ? _GEN_10415 : dirty_0_13; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11447 = 3'h5 == state ? _GEN_10416 : dirty_0_14; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11448 = 3'h5 == state ? _GEN_10417 : dirty_0_15; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11449 = 3'h5 == state ? _GEN_10418 : dirty_0_16; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11450 = 3'h5 == state ? _GEN_10419 : dirty_0_17; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11451 = 3'h5 == state ? _GEN_10420 : dirty_0_18; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11452 = 3'h5 == state ? _GEN_10421 : dirty_0_19; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11453 = 3'h5 == state ? _GEN_10422 : dirty_0_20; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11454 = 3'h5 == state ? _GEN_10423 : dirty_0_21; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11455 = 3'h5 == state ? _GEN_10424 : dirty_0_22; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11456 = 3'h5 == state ? _GEN_10425 : dirty_0_23; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11457 = 3'h5 == state ? _GEN_10426 : dirty_0_24; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11458 = 3'h5 == state ? _GEN_10427 : dirty_0_25; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11459 = 3'h5 == state ? _GEN_10428 : dirty_0_26; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11460 = 3'h5 == state ? _GEN_10429 : dirty_0_27; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11461 = 3'h5 == state ? _GEN_10430 : dirty_0_28; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11462 = 3'h5 == state ? _GEN_10431 : dirty_0_29; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11463 = 3'h5 == state ? _GEN_10432 : dirty_0_30; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11464 = 3'h5 == state ? _GEN_10433 : dirty_0_31; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11465 = 3'h5 == state ? _GEN_10434 : dirty_0_32; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11466 = 3'h5 == state ? _GEN_10435 : dirty_0_33; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11467 = 3'h5 == state ? _GEN_10436 : dirty_0_34; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11468 = 3'h5 == state ? _GEN_10437 : dirty_0_35; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11469 = 3'h5 == state ? _GEN_10438 : dirty_0_36; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11470 = 3'h5 == state ? _GEN_10439 : dirty_0_37; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11471 = 3'h5 == state ? _GEN_10440 : dirty_0_38; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11472 = 3'h5 == state ? _GEN_10441 : dirty_0_39; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11473 = 3'h5 == state ? _GEN_10442 : dirty_0_40; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11474 = 3'h5 == state ? _GEN_10443 : dirty_0_41; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11475 = 3'h5 == state ? _GEN_10444 : dirty_0_42; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11476 = 3'h5 == state ? _GEN_10445 : dirty_0_43; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11477 = 3'h5 == state ? _GEN_10446 : dirty_0_44; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11478 = 3'h5 == state ? _GEN_10447 : dirty_0_45; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11479 = 3'h5 == state ? _GEN_10448 : dirty_0_46; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11480 = 3'h5 == state ? _GEN_10449 : dirty_0_47; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11481 = 3'h5 == state ? _GEN_10450 : dirty_0_48; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11482 = 3'h5 == state ? _GEN_10451 : dirty_0_49; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11483 = 3'h5 == state ? _GEN_10452 : dirty_0_50; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11484 = 3'h5 == state ? _GEN_10453 : dirty_0_51; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11485 = 3'h5 == state ? _GEN_10454 : dirty_0_52; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11486 = 3'h5 == state ? _GEN_10455 : dirty_0_53; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11487 = 3'h5 == state ? _GEN_10456 : dirty_0_54; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11488 = 3'h5 == state ? _GEN_10457 : dirty_0_55; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11489 = 3'h5 == state ? _GEN_10458 : dirty_0_56; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11490 = 3'h5 == state ? _GEN_10459 : dirty_0_57; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11491 = 3'h5 == state ? _GEN_10460 : dirty_0_58; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11492 = 3'h5 == state ? _GEN_10461 : dirty_0_59; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11493 = 3'h5 == state ? _GEN_10462 : dirty_0_60; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11494 = 3'h5 == state ? _GEN_10463 : dirty_0_61; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11495 = 3'h5 == state ? _GEN_10464 : dirty_0_62; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11496 = 3'h5 == state ? _GEN_10465 : dirty_0_63; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11497 = 3'h5 == state ? _GEN_10466 : dirty_0_64; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11498 = 3'h5 == state ? _GEN_10467 : dirty_0_65; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11499 = 3'h5 == state ? _GEN_10468 : dirty_0_66; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11500 = 3'h5 == state ? _GEN_10469 : dirty_0_67; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11501 = 3'h5 == state ? _GEN_10470 : dirty_0_68; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11502 = 3'h5 == state ? _GEN_10471 : dirty_0_69; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11503 = 3'h5 == state ? _GEN_10472 : dirty_0_70; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11504 = 3'h5 == state ? _GEN_10473 : dirty_0_71; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11505 = 3'h5 == state ? _GEN_10474 : dirty_0_72; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11506 = 3'h5 == state ? _GEN_10475 : dirty_0_73; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11507 = 3'h5 == state ? _GEN_10476 : dirty_0_74; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11508 = 3'h5 == state ? _GEN_10477 : dirty_0_75; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11509 = 3'h5 == state ? _GEN_10478 : dirty_0_76; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11510 = 3'h5 == state ? _GEN_10479 : dirty_0_77; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11511 = 3'h5 == state ? _GEN_10480 : dirty_0_78; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11512 = 3'h5 == state ? _GEN_10481 : dirty_0_79; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11513 = 3'h5 == state ? _GEN_10482 : dirty_0_80; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11514 = 3'h5 == state ? _GEN_10483 : dirty_0_81; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11515 = 3'h5 == state ? _GEN_10484 : dirty_0_82; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11516 = 3'h5 == state ? _GEN_10485 : dirty_0_83; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11517 = 3'h5 == state ? _GEN_10486 : dirty_0_84; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11518 = 3'h5 == state ? _GEN_10487 : dirty_0_85; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11519 = 3'h5 == state ? _GEN_10488 : dirty_0_86; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11520 = 3'h5 == state ? _GEN_10489 : dirty_0_87; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11521 = 3'h5 == state ? _GEN_10490 : dirty_0_88; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11522 = 3'h5 == state ? _GEN_10491 : dirty_0_89; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11523 = 3'h5 == state ? _GEN_10492 : dirty_0_90; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11524 = 3'h5 == state ? _GEN_10493 : dirty_0_91; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11525 = 3'h5 == state ? _GEN_10494 : dirty_0_92; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11526 = 3'h5 == state ? _GEN_10495 : dirty_0_93; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11527 = 3'h5 == state ? _GEN_10496 : dirty_0_94; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11528 = 3'h5 == state ? _GEN_10497 : dirty_0_95; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11529 = 3'h5 == state ? _GEN_10498 : dirty_0_96; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11530 = 3'h5 == state ? _GEN_10499 : dirty_0_97; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11531 = 3'h5 == state ? _GEN_10500 : dirty_0_98; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11532 = 3'h5 == state ? _GEN_10501 : dirty_0_99; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11533 = 3'h5 == state ? _GEN_10502 : dirty_0_100; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11534 = 3'h5 == state ? _GEN_10503 : dirty_0_101; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11535 = 3'h5 == state ? _GEN_10504 : dirty_0_102; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11536 = 3'h5 == state ? _GEN_10505 : dirty_0_103; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11537 = 3'h5 == state ? _GEN_10506 : dirty_0_104; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11538 = 3'h5 == state ? _GEN_10507 : dirty_0_105; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11539 = 3'h5 == state ? _GEN_10508 : dirty_0_106; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11540 = 3'h5 == state ? _GEN_10509 : dirty_0_107; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11541 = 3'h5 == state ? _GEN_10510 : dirty_0_108; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11542 = 3'h5 == state ? _GEN_10511 : dirty_0_109; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11543 = 3'h5 == state ? _GEN_10512 : dirty_0_110; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11544 = 3'h5 == state ? _GEN_10513 : dirty_0_111; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11545 = 3'h5 == state ? _GEN_10514 : dirty_0_112; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11546 = 3'h5 == state ? _GEN_10515 : dirty_0_113; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11547 = 3'h5 == state ? _GEN_10516 : dirty_0_114; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11548 = 3'h5 == state ? _GEN_10517 : dirty_0_115; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11549 = 3'h5 == state ? _GEN_10518 : dirty_0_116; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11550 = 3'h5 == state ? _GEN_10519 : dirty_0_117; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11551 = 3'h5 == state ? _GEN_10520 : dirty_0_118; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11552 = 3'h5 == state ? _GEN_10521 : dirty_0_119; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11553 = 3'h5 == state ? _GEN_10522 : dirty_0_120; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11554 = 3'h5 == state ? _GEN_10523 : dirty_0_121; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11555 = 3'h5 == state ? _GEN_10524 : dirty_0_122; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11556 = 3'h5 == state ? _GEN_10525 : dirty_0_123; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11557 = 3'h5 == state ? _GEN_10526 : dirty_0_124; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11558 = 3'h5 == state ? _GEN_10527 : dirty_0_125; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11559 = 3'h5 == state ? _GEN_10528 : dirty_0_126; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11560 = 3'h5 == state ? _GEN_10529 : dirty_0_127; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_11561 = 3'h5 == state ? _GEN_10530 : dirty_1_0; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11562 = 3'h5 == state ? _GEN_10531 : dirty_1_1; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11563 = 3'h5 == state ? _GEN_10532 : dirty_1_2; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11564 = 3'h5 == state ? _GEN_10533 : dirty_1_3; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11565 = 3'h5 == state ? _GEN_10534 : dirty_1_4; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11566 = 3'h5 == state ? _GEN_10535 : dirty_1_5; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11567 = 3'h5 == state ? _GEN_10536 : dirty_1_6; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11568 = 3'h5 == state ? _GEN_10537 : dirty_1_7; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11569 = 3'h5 == state ? _GEN_10538 : dirty_1_8; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11570 = 3'h5 == state ? _GEN_10539 : dirty_1_9; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11571 = 3'h5 == state ? _GEN_10540 : dirty_1_10; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11572 = 3'h5 == state ? _GEN_10541 : dirty_1_11; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11573 = 3'h5 == state ? _GEN_10542 : dirty_1_12; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11574 = 3'h5 == state ? _GEN_10543 : dirty_1_13; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11575 = 3'h5 == state ? _GEN_10544 : dirty_1_14; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11576 = 3'h5 == state ? _GEN_10545 : dirty_1_15; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11577 = 3'h5 == state ? _GEN_10546 : dirty_1_16; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11578 = 3'h5 == state ? _GEN_10547 : dirty_1_17; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11579 = 3'h5 == state ? _GEN_10548 : dirty_1_18; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11580 = 3'h5 == state ? _GEN_10549 : dirty_1_19; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11581 = 3'h5 == state ? _GEN_10550 : dirty_1_20; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11582 = 3'h5 == state ? _GEN_10551 : dirty_1_21; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11583 = 3'h5 == state ? _GEN_10552 : dirty_1_22; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11584 = 3'h5 == state ? _GEN_10553 : dirty_1_23; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11585 = 3'h5 == state ? _GEN_10554 : dirty_1_24; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11586 = 3'h5 == state ? _GEN_10555 : dirty_1_25; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11587 = 3'h5 == state ? _GEN_10556 : dirty_1_26; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11588 = 3'h5 == state ? _GEN_10557 : dirty_1_27; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11589 = 3'h5 == state ? _GEN_10558 : dirty_1_28; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11590 = 3'h5 == state ? _GEN_10559 : dirty_1_29; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11591 = 3'h5 == state ? _GEN_10560 : dirty_1_30; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11592 = 3'h5 == state ? _GEN_10561 : dirty_1_31; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11593 = 3'h5 == state ? _GEN_10562 : dirty_1_32; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11594 = 3'h5 == state ? _GEN_10563 : dirty_1_33; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11595 = 3'h5 == state ? _GEN_10564 : dirty_1_34; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11596 = 3'h5 == state ? _GEN_10565 : dirty_1_35; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11597 = 3'h5 == state ? _GEN_10566 : dirty_1_36; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11598 = 3'h5 == state ? _GEN_10567 : dirty_1_37; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11599 = 3'h5 == state ? _GEN_10568 : dirty_1_38; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11600 = 3'h5 == state ? _GEN_10569 : dirty_1_39; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11601 = 3'h5 == state ? _GEN_10570 : dirty_1_40; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11602 = 3'h5 == state ? _GEN_10571 : dirty_1_41; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11603 = 3'h5 == state ? _GEN_10572 : dirty_1_42; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11604 = 3'h5 == state ? _GEN_10573 : dirty_1_43; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11605 = 3'h5 == state ? _GEN_10574 : dirty_1_44; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11606 = 3'h5 == state ? _GEN_10575 : dirty_1_45; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11607 = 3'h5 == state ? _GEN_10576 : dirty_1_46; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11608 = 3'h5 == state ? _GEN_10577 : dirty_1_47; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11609 = 3'h5 == state ? _GEN_10578 : dirty_1_48; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11610 = 3'h5 == state ? _GEN_10579 : dirty_1_49; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11611 = 3'h5 == state ? _GEN_10580 : dirty_1_50; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11612 = 3'h5 == state ? _GEN_10581 : dirty_1_51; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11613 = 3'h5 == state ? _GEN_10582 : dirty_1_52; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11614 = 3'h5 == state ? _GEN_10583 : dirty_1_53; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11615 = 3'h5 == state ? _GEN_10584 : dirty_1_54; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11616 = 3'h5 == state ? _GEN_10585 : dirty_1_55; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11617 = 3'h5 == state ? _GEN_10586 : dirty_1_56; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11618 = 3'h5 == state ? _GEN_10587 : dirty_1_57; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11619 = 3'h5 == state ? _GEN_10588 : dirty_1_58; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11620 = 3'h5 == state ? _GEN_10589 : dirty_1_59; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11621 = 3'h5 == state ? _GEN_10590 : dirty_1_60; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11622 = 3'h5 == state ? _GEN_10591 : dirty_1_61; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11623 = 3'h5 == state ? _GEN_10592 : dirty_1_62; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11624 = 3'h5 == state ? _GEN_10593 : dirty_1_63; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11625 = 3'h5 == state ? _GEN_10594 : dirty_1_64; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11626 = 3'h5 == state ? _GEN_10595 : dirty_1_65; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11627 = 3'h5 == state ? _GEN_10596 : dirty_1_66; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11628 = 3'h5 == state ? _GEN_10597 : dirty_1_67; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11629 = 3'h5 == state ? _GEN_10598 : dirty_1_68; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11630 = 3'h5 == state ? _GEN_10599 : dirty_1_69; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11631 = 3'h5 == state ? _GEN_10600 : dirty_1_70; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11632 = 3'h5 == state ? _GEN_10601 : dirty_1_71; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11633 = 3'h5 == state ? _GEN_10602 : dirty_1_72; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11634 = 3'h5 == state ? _GEN_10603 : dirty_1_73; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11635 = 3'h5 == state ? _GEN_10604 : dirty_1_74; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11636 = 3'h5 == state ? _GEN_10605 : dirty_1_75; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11637 = 3'h5 == state ? _GEN_10606 : dirty_1_76; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11638 = 3'h5 == state ? _GEN_10607 : dirty_1_77; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11639 = 3'h5 == state ? _GEN_10608 : dirty_1_78; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11640 = 3'h5 == state ? _GEN_10609 : dirty_1_79; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11641 = 3'h5 == state ? _GEN_10610 : dirty_1_80; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11642 = 3'h5 == state ? _GEN_10611 : dirty_1_81; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11643 = 3'h5 == state ? _GEN_10612 : dirty_1_82; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11644 = 3'h5 == state ? _GEN_10613 : dirty_1_83; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11645 = 3'h5 == state ? _GEN_10614 : dirty_1_84; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11646 = 3'h5 == state ? _GEN_10615 : dirty_1_85; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11647 = 3'h5 == state ? _GEN_10616 : dirty_1_86; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11648 = 3'h5 == state ? _GEN_10617 : dirty_1_87; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11649 = 3'h5 == state ? _GEN_10618 : dirty_1_88; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11650 = 3'h5 == state ? _GEN_10619 : dirty_1_89; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11651 = 3'h5 == state ? _GEN_10620 : dirty_1_90; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11652 = 3'h5 == state ? _GEN_10621 : dirty_1_91; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11653 = 3'h5 == state ? _GEN_10622 : dirty_1_92; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11654 = 3'h5 == state ? _GEN_10623 : dirty_1_93; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11655 = 3'h5 == state ? _GEN_10624 : dirty_1_94; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11656 = 3'h5 == state ? _GEN_10625 : dirty_1_95; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11657 = 3'h5 == state ? _GEN_10626 : dirty_1_96; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11658 = 3'h5 == state ? _GEN_10627 : dirty_1_97; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11659 = 3'h5 == state ? _GEN_10628 : dirty_1_98; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11660 = 3'h5 == state ? _GEN_10629 : dirty_1_99; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11661 = 3'h5 == state ? _GEN_10630 : dirty_1_100; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11662 = 3'h5 == state ? _GEN_10631 : dirty_1_101; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11663 = 3'h5 == state ? _GEN_10632 : dirty_1_102; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11664 = 3'h5 == state ? _GEN_10633 : dirty_1_103; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11665 = 3'h5 == state ? _GEN_10634 : dirty_1_104; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11666 = 3'h5 == state ? _GEN_10635 : dirty_1_105; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11667 = 3'h5 == state ? _GEN_10636 : dirty_1_106; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11668 = 3'h5 == state ? _GEN_10637 : dirty_1_107; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11669 = 3'h5 == state ? _GEN_10638 : dirty_1_108; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11670 = 3'h5 == state ? _GEN_10639 : dirty_1_109; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11671 = 3'h5 == state ? _GEN_10640 : dirty_1_110; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11672 = 3'h5 == state ? _GEN_10641 : dirty_1_111; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11673 = 3'h5 == state ? _GEN_10642 : dirty_1_112; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11674 = 3'h5 == state ? _GEN_10643 : dirty_1_113; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11675 = 3'h5 == state ? _GEN_10644 : dirty_1_114; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11676 = 3'h5 == state ? _GEN_10645 : dirty_1_115; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11677 = 3'h5 == state ? _GEN_10646 : dirty_1_116; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11678 = 3'h5 == state ? _GEN_10647 : dirty_1_117; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11679 = 3'h5 == state ? _GEN_10648 : dirty_1_118; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11680 = 3'h5 == state ? _GEN_10649 : dirty_1_119; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11681 = 3'h5 == state ? _GEN_10650 : dirty_1_120; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11682 = 3'h5 == state ? _GEN_10651 : dirty_1_121; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11683 = 3'h5 == state ? _GEN_10652 : dirty_1_122; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11684 = 3'h5 == state ? _GEN_10653 : dirty_1_123; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11685 = 3'h5 == state ? _GEN_10654 : dirty_1_124; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11686 = 3'h5 == state ? _GEN_10655 : dirty_1_125; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11687 = 3'h5 == state ? _GEN_10656 : dirty_1_126; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_11688 = 3'h5 == state ? _GEN_10657 : dirty_1_127; // @[d_cache.scala 81:18 27:26]
  wire [2:0] _GEN_11689 = 3'h4 == state ? _GEN_3213 : _GEN_10661; // @[d_cache.scala 81:18]
  wire [63:0] _GEN_11690 = 3'h4 == state ? ram_0_0 : _GEN_10662; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11691 = 3'h4 == state ? ram_0_1 : _GEN_10663; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11692 = 3'h4 == state ? ram_0_2 : _GEN_10664; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11693 = 3'h4 == state ? ram_0_3 : _GEN_10665; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11694 = 3'h4 == state ? ram_0_4 : _GEN_10666; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11695 = 3'h4 == state ? ram_0_5 : _GEN_10667; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11696 = 3'h4 == state ? ram_0_6 : _GEN_10668; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11697 = 3'h4 == state ? ram_0_7 : _GEN_10669; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11698 = 3'h4 == state ? ram_0_8 : _GEN_10670; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11699 = 3'h4 == state ? ram_0_9 : _GEN_10671; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11700 = 3'h4 == state ? ram_0_10 : _GEN_10672; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11701 = 3'h4 == state ? ram_0_11 : _GEN_10673; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11702 = 3'h4 == state ? ram_0_12 : _GEN_10674; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11703 = 3'h4 == state ? ram_0_13 : _GEN_10675; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11704 = 3'h4 == state ? ram_0_14 : _GEN_10676; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11705 = 3'h4 == state ? ram_0_15 : _GEN_10677; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11706 = 3'h4 == state ? ram_0_16 : _GEN_10678; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11707 = 3'h4 == state ? ram_0_17 : _GEN_10679; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11708 = 3'h4 == state ? ram_0_18 : _GEN_10680; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11709 = 3'h4 == state ? ram_0_19 : _GEN_10681; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11710 = 3'h4 == state ? ram_0_20 : _GEN_10682; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11711 = 3'h4 == state ? ram_0_21 : _GEN_10683; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11712 = 3'h4 == state ? ram_0_22 : _GEN_10684; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11713 = 3'h4 == state ? ram_0_23 : _GEN_10685; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11714 = 3'h4 == state ? ram_0_24 : _GEN_10686; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11715 = 3'h4 == state ? ram_0_25 : _GEN_10687; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11716 = 3'h4 == state ? ram_0_26 : _GEN_10688; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11717 = 3'h4 == state ? ram_0_27 : _GEN_10689; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11718 = 3'h4 == state ? ram_0_28 : _GEN_10690; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11719 = 3'h4 == state ? ram_0_29 : _GEN_10691; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11720 = 3'h4 == state ? ram_0_30 : _GEN_10692; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11721 = 3'h4 == state ? ram_0_31 : _GEN_10693; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11722 = 3'h4 == state ? ram_0_32 : _GEN_10694; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11723 = 3'h4 == state ? ram_0_33 : _GEN_10695; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11724 = 3'h4 == state ? ram_0_34 : _GEN_10696; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11725 = 3'h4 == state ? ram_0_35 : _GEN_10697; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11726 = 3'h4 == state ? ram_0_36 : _GEN_10698; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11727 = 3'h4 == state ? ram_0_37 : _GEN_10699; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11728 = 3'h4 == state ? ram_0_38 : _GEN_10700; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11729 = 3'h4 == state ? ram_0_39 : _GEN_10701; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11730 = 3'h4 == state ? ram_0_40 : _GEN_10702; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11731 = 3'h4 == state ? ram_0_41 : _GEN_10703; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11732 = 3'h4 == state ? ram_0_42 : _GEN_10704; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11733 = 3'h4 == state ? ram_0_43 : _GEN_10705; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11734 = 3'h4 == state ? ram_0_44 : _GEN_10706; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11735 = 3'h4 == state ? ram_0_45 : _GEN_10707; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11736 = 3'h4 == state ? ram_0_46 : _GEN_10708; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11737 = 3'h4 == state ? ram_0_47 : _GEN_10709; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11738 = 3'h4 == state ? ram_0_48 : _GEN_10710; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11739 = 3'h4 == state ? ram_0_49 : _GEN_10711; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11740 = 3'h4 == state ? ram_0_50 : _GEN_10712; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11741 = 3'h4 == state ? ram_0_51 : _GEN_10713; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11742 = 3'h4 == state ? ram_0_52 : _GEN_10714; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11743 = 3'h4 == state ? ram_0_53 : _GEN_10715; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11744 = 3'h4 == state ? ram_0_54 : _GEN_10716; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11745 = 3'h4 == state ? ram_0_55 : _GEN_10717; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11746 = 3'h4 == state ? ram_0_56 : _GEN_10718; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11747 = 3'h4 == state ? ram_0_57 : _GEN_10719; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11748 = 3'h4 == state ? ram_0_58 : _GEN_10720; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11749 = 3'h4 == state ? ram_0_59 : _GEN_10721; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11750 = 3'h4 == state ? ram_0_60 : _GEN_10722; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11751 = 3'h4 == state ? ram_0_61 : _GEN_10723; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11752 = 3'h4 == state ? ram_0_62 : _GEN_10724; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11753 = 3'h4 == state ? ram_0_63 : _GEN_10725; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11754 = 3'h4 == state ? ram_0_64 : _GEN_10726; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11755 = 3'h4 == state ? ram_0_65 : _GEN_10727; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11756 = 3'h4 == state ? ram_0_66 : _GEN_10728; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11757 = 3'h4 == state ? ram_0_67 : _GEN_10729; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11758 = 3'h4 == state ? ram_0_68 : _GEN_10730; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11759 = 3'h4 == state ? ram_0_69 : _GEN_10731; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11760 = 3'h4 == state ? ram_0_70 : _GEN_10732; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11761 = 3'h4 == state ? ram_0_71 : _GEN_10733; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11762 = 3'h4 == state ? ram_0_72 : _GEN_10734; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11763 = 3'h4 == state ? ram_0_73 : _GEN_10735; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11764 = 3'h4 == state ? ram_0_74 : _GEN_10736; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11765 = 3'h4 == state ? ram_0_75 : _GEN_10737; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11766 = 3'h4 == state ? ram_0_76 : _GEN_10738; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11767 = 3'h4 == state ? ram_0_77 : _GEN_10739; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11768 = 3'h4 == state ? ram_0_78 : _GEN_10740; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11769 = 3'h4 == state ? ram_0_79 : _GEN_10741; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11770 = 3'h4 == state ? ram_0_80 : _GEN_10742; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11771 = 3'h4 == state ? ram_0_81 : _GEN_10743; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11772 = 3'h4 == state ? ram_0_82 : _GEN_10744; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11773 = 3'h4 == state ? ram_0_83 : _GEN_10745; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11774 = 3'h4 == state ? ram_0_84 : _GEN_10746; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11775 = 3'h4 == state ? ram_0_85 : _GEN_10747; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11776 = 3'h4 == state ? ram_0_86 : _GEN_10748; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11777 = 3'h4 == state ? ram_0_87 : _GEN_10749; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11778 = 3'h4 == state ? ram_0_88 : _GEN_10750; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11779 = 3'h4 == state ? ram_0_89 : _GEN_10751; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11780 = 3'h4 == state ? ram_0_90 : _GEN_10752; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11781 = 3'h4 == state ? ram_0_91 : _GEN_10753; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11782 = 3'h4 == state ? ram_0_92 : _GEN_10754; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11783 = 3'h4 == state ? ram_0_93 : _GEN_10755; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11784 = 3'h4 == state ? ram_0_94 : _GEN_10756; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11785 = 3'h4 == state ? ram_0_95 : _GEN_10757; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11786 = 3'h4 == state ? ram_0_96 : _GEN_10758; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11787 = 3'h4 == state ? ram_0_97 : _GEN_10759; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11788 = 3'h4 == state ? ram_0_98 : _GEN_10760; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11789 = 3'h4 == state ? ram_0_99 : _GEN_10761; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11790 = 3'h4 == state ? ram_0_100 : _GEN_10762; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11791 = 3'h4 == state ? ram_0_101 : _GEN_10763; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11792 = 3'h4 == state ? ram_0_102 : _GEN_10764; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11793 = 3'h4 == state ? ram_0_103 : _GEN_10765; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11794 = 3'h4 == state ? ram_0_104 : _GEN_10766; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11795 = 3'h4 == state ? ram_0_105 : _GEN_10767; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11796 = 3'h4 == state ? ram_0_106 : _GEN_10768; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11797 = 3'h4 == state ? ram_0_107 : _GEN_10769; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11798 = 3'h4 == state ? ram_0_108 : _GEN_10770; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11799 = 3'h4 == state ? ram_0_109 : _GEN_10771; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11800 = 3'h4 == state ? ram_0_110 : _GEN_10772; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11801 = 3'h4 == state ? ram_0_111 : _GEN_10773; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11802 = 3'h4 == state ? ram_0_112 : _GEN_10774; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11803 = 3'h4 == state ? ram_0_113 : _GEN_10775; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11804 = 3'h4 == state ? ram_0_114 : _GEN_10776; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11805 = 3'h4 == state ? ram_0_115 : _GEN_10777; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11806 = 3'h4 == state ? ram_0_116 : _GEN_10778; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11807 = 3'h4 == state ? ram_0_117 : _GEN_10779; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11808 = 3'h4 == state ? ram_0_118 : _GEN_10780; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11809 = 3'h4 == state ? ram_0_119 : _GEN_10781; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11810 = 3'h4 == state ? ram_0_120 : _GEN_10782; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11811 = 3'h4 == state ? ram_0_121 : _GEN_10783; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11812 = 3'h4 == state ? ram_0_122 : _GEN_10784; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11813 = 3'h4 == state ? ram_0_123 : _GEN_10785; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11814 = 3'h4 == state ? ram_0_124 : _GEN_10786; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11815 = 3'h4 == state ? ram_0_125 : _GEN_10787; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11816 = 3'h4 == state ? ram_0_126 : _GEN_10788; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_11817 = 3'h4 == state ? ram_0_127 : _GEN_10789; // @[d_cache.scala 81:18 18:24]
  wire [31:0] _GEN_11818 = 3'h4 == state ? tag_0_0 : _GEN_10790; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11819 = 3'h4 == state ? tag_0_1 : _GEN_10791; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11820 = 3'h4 == state ? tag_0_2 : _GEN_10792; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11821 = 3'h4 == state ? tag_0_3 : _GEN_10793; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11822 = 3'h4 == state ? tag_0_4 : _GEN_10794; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11823 = 3'h4 == state ? tag_0_5 : _GEN_10795; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11824 = 3'h4 == state ? tag_0_6 : _GEN_10796; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11825 = 3'h4 == state ? tag_0_7 : _GEN_10797; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11826 = 3'h4 == state ? tag_0_8 : _GEN_10798; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11827 = 3'h4 == state ? tag_0_9 : _GEN_10799; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11828 = 3'h4 == state ? tag_0_10 : _GEN_10800; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11829 = 3'h4 == state ? tag_0_11 : _GEN_10801; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11830 = 3'h4 == state ? tag_0_12 : _GEN_10802; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11831 = 3'h4 == state ? tag_0_13 : _GEN_10803; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11832 = 3'h4 == state ? tag_0_14 : _GEN_10804; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11833 = 3'h4 == state ? tag_0_15 : _GEN_10805; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11834 = 3'h4 == state ? tag_0_16 : _GEN_10806; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11835 = 3'h4 == state ? tag_0_17 : _GEN_10807; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11836 = 3'h4 == state ? tag_0_18 : _GEN_10808; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11837 = 3'h4 == state ? tag_0_19 : _GEN_10809; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11838 = 3'h4 == state ? tag_0_20 : _GEN_10810; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11839 = 3'h4 == state ? tag_0_21 : _GEN_10811; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11840 = 3'h4 == state ? tag_0_22 : _GEN_10812; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11841 = 3'h4 == state ? tag_0_23 : _GEN_10813; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11842 = 3'h4 == state ? tag_0_24 : _GEN_10814; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11843 = 3'h4 == state ? tag_0_25 : _GEN_10815; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11844 = 3'h4 == state ? tag_0_26 : _GEN_10816; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11845 = 3'h4 == state ? tag_0_27 : _GEN_10817; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11846 = 3'h4 == state ? tag_0_28 : _GEN_10818; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11847 = 3'h4 == state ? tag_0_29 : _GEN_10819; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11848 = 3'h4 == state ? tag_0_30 : _GEN_10820; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11849 = 3'h4 == state ? tag_0_31 : _GEN_10821; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11850 = 3'h4 == state ? tag_0_32 : _GEN_10822; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11851 = 3'h4 == state ? tag_0_33 : _GEN_10823; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11852 = 3'h4 == state ? tag_0_34 : _GEN_10824; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11853 = 3'h4 == state ? tag_0_35 : _GEN_10825; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11854 = 3'h4 == state ? tag_0_36 : _GEN_10826; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11855 = 3'h4 == state ? tag_0_37 : _GEN_10827; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11856 = 3'h4 == state ? tag_0_38 : _GEN_10828; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11857 = 3'h4 == state ? tag_0_39 : _GEN_10829; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11858 = 3'h4 == state ? tag_0_40 : _GEN_10830; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11859 = 3'h4 == state ? tag_0_41 : _GEN_10831; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11860 = 3'h4 == state ? tag_0_42 : _GEN_10832; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11861 = 3'h4 == state ? tag_0_43 : _GEN_10833; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11862 = 3'h4 == state ? tag_0_44 : _GEN_10834; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11863 = 3'h4 == state ? tag_0_45 : _GEN_10835; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11864 = 3'h4 == state ? tag_0_46 : _GEN_10836; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11865 = 3'h4 == state ? tag_0_47 : _GEN_10837; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11866 = 3'h4 == state ? tag_0_48 : _GEN_10838; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11867 = 3'h4 == state ? tag_0_49 : _GEN_10839; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11868 = 3'h4 == state ? tag_0_50 : _GEN_10840; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11869 = 3'h4 == state ? tag_0_51 : _GEN_10841; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11870 = 3'h4 == state ? tag_0_52 : _GEN_10842; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11871 = 3'h4 == state ? tag_0_53 : _GEN_10843; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11872 = 3'h4 == state ? tag_0_54 : _GEN_10844; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11873 = 3'h4 == state ? tag_0_55 : _GEN_10845; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11874 = 3'h4 == state ? tag_0_56 : _GEN_10846; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11875 = 3'h4 == state ? tag_0_57 : _GEN_10847; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11876 = 3'h4 == state ? tag_0_58 : _GEN_10848; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11877 = 3'h4 == state ? tag_0_59 : _GEN_10849; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11878 = 3'h4 == state ? tag_0_60 : _GEN_10850; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11879 = 3'h4 == state ? tag_0_61 : _GEN_10851; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11880 = 3'h4 == state ? tag_0_62 : _GEN_10852; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11881 = 3'h4 == state ? tag_0_63 : _GEN_10853; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11882 = 3'h4 == state ? tag_0_64 : _GEN_10854; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11883 = 3'h4 == state ? tag_0_65 : _GEN_10855; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11884 = 3'h4 == state ? tag_0_66 : _GEN_10856; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11885 = 3'h4 == state ? tag_0_67 : _GEN_10857; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11886 = 3'h4 == state ? tag_0_68 : _GEN_10858; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11887 = 3'h4 == state ? tag_0_69 : _GEN_10859; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11888 = 3'h4 == state ? tag_0_70 : _GEN_10860; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11889 = 3'h4 == state ? tag_0_71 : _GEN_10861; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11890 = 3'h4 == state ? tag_0_72 : _GEN_10862; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11891 = 3'h4 == state ? tag_0_73 : _GEN_10863; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11892 = 3'h4 == state ? tag_0_74 : _GEN_10864; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11893 = 3'h4 == state ? tag_0_75 : _GEN_10865; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11894 = 3'h4 == state ? tag_0_76 : _GEN_10866; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11895 = 3'h4 == state ? tag_0_77 : _GEN_10867; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11896 = 3'h4 == state ? tag_0_78 : _GEN_10868; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11897 = 3'h4 == state ? tag_0_79 : _GEN_10869; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11898 = 3'h4 == state ? tag_0_80 : _GEN_10870; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11899 = 3'h4 == state ? tag_0_81 : _GEN_10871; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11900 = 3'h4 == state ? tag_0_82 : _GEN_10872; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11901 = 3'h4 == state ? tag_0_83 : _GEN_10873; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11902 = 3'h4 == state ? tag_0_84 : _GEN_10874; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11903 = 3'h4 == state ? tag_0_85 : _GEN_10875; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11904 = 3'h4 == state ? tag_0_86 : _GEN_10876; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11905 = 3'h4 == state ? tag_0_87 : _GEN_10877; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11906 = 3'h4 == state ? tag_0_88 : _GEN_10878; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11907 = 3'h4 == state ? tag_0_89 : _GEN_10879; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11908 = 3'h4 == state ? tag_0_90 : _GEN_10880; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11909 = 3'h4 == state ? tag_0_91 : _GEN_10881; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11910 = 3'h4 == state ? tag_0_92 : _GEN_10882; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11911 = 3'h4 == state ? tag_0_93 : _GEN_10883; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11912 = 3'h4 == state ? tag_0_94 : _GEN_10884; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11913 = 3'h4 == state ? tag_0_95 : _GEN_10885; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11914 = 3'h4 == state ? tag_0_96 : _GEN_10886; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11915 = 3'h4 == state ? tag_0_97 : _GEN_10887; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11916 = 3'h4 == state ? tag_0_98 : _GEN_10888; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11917 = 3'h4 == state ? tag_0_99 : _GEN_10889; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11918 = 3'h4 == state ? tag_0_100 : _GEN_10890; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11919 = 3'h4 == state ? tag_0_101 : _GEN_10891; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11920 = 3'h4 == state ? tag_0_102 : _GEN_10892; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11921 = 3'h4 == state ? tag_0_103 : _GEN_10893; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11922 = 3'h4 == state ? tag_0_104 : _GEN_10894; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11923 = 3'h4 == state ? tag_0_105 : _GEN_10895; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11924 = 3'h4 == state ? tag_0_106 : _GEN_10896; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11925 = 3'h4 == state ? tag_0_107 : _GEN_10897; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11926 = 3'h4 == state ? tag_0_108 : _GEN_10898; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11927 = 3'h4 == state ? tag_0_109 : _GEN_10899; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11928 = 3'h4 == state ? tag_0_110 : _GEN_10900; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11929 = 3'h4 == state ? tag_0_111 : _GEN_10901; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11930 = 3'h4 == state ? tag_0_112 : _GEN_10902; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11931 = 3'h4 == state ? tag_0_113 : _GEN_10903; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11932 = 3'h4 == state ? tag_0_114 : _GEN_10904; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11933 = 3'h4 == state ? tag_0_115 : _GEN_10905; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11934 = 3'h4 == state ? tag_0_116 : _GEN_10906; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11935 = 3'h4 == state ? tag_0_117 : _GEN_10907; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11936 = 3'h4 == state ? tag_0_118 : _GEN_10908; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11937 = 3'h4 == state ? tag_0_119 : _GEN_10909; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11938 = 3'h4 == state ? tag_0_120 : _GEN_10910; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11939 = 3'h4 == state ? tag_0_121 : _GEN_10911; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11940 = 3'h4 == state ? tag_0_122 : _GEN_10912; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11941 = 3'h4 == state ? tag_0_123 : _GEN_10913; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11942 = 3'h4 == state ? tag_0_124 : _GEN_10914; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11943 = 3'h4 == state ? tag_0_125 : _GEN_10915; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11944 = 3'h4 == state ? tag_0_126 : _GEN_10916; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_11945 = 3'h4 == state ? tag_0_127 : _GEN_10917; // @[d_cache.scala 81:18 22:24]
  wire  _GEN_11946 = 3'h4 == state ? valid_0_0 : _GEN_10918; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11947 = 3'h4 == state ? valid_0_1 : _GEN_10919; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11948 = 3'h4 == state ? valid_0_2 : _GEN_10920; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11949 = 3'h4 == state ? valid_0_3 : _GEN_10921; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11950 = 3'h4 == state ? valid_0_4 : _GEN_10922; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11951 = 3'h4 == state ? valid_0_5 : _GEN_10923; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11952 = 3'h4 == state ? valid_0_6 : _GEN_10924; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11953 = 3'h4 == state ? valid_0_7 : _GEN_10925; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11954 = 3'h4 == state ? valid_0_8 : _GEN_10926; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11955 = 3'h4 == state ? valid_0_9 : _GEN_10927; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11956 = 3'h4 == state ? valid_0_10 : _GEN_10928; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11957 = 3'h4 == state ? valid_0_11 : _GEN_10929; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11958 = 3'h4 == state ? valid_0_12 : _GEN_10930; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11959 = 3'h4 == state ? valid_0_13 : _GEN_10931; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11960 = 3'h4 == state ? valid_0_14 : _GEN_10932; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11961 = 3'h4 == state ? valid_0_15 : _GEN_10933; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11962 = 3'h4 == state ? valid_0_16 : _GEN_10934; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11963 = 3'h4 == state ? valid_0_17 : _GEN_10935; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11964 = 3'h4 == state ? valid_0_18 : _GEN_10936; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11965 = 3'h4 == state ? valid_0_19 : _GEN_10937; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11966 = 3'h4 == state ? valid_0_20 : _GEN_10938; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11967 = 3'h4 == state ? valid_0_21 : _GEN_10939; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11968 = 3'h4 == state ? valid_0_22 : _GEN_10940; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11969 = 3'h4 == state ? valid_0_23 : _GEN_10941; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11970 = 3'h4 == state ? valid_0_24 : _GEN_10942; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11971 = 3'h4 == state ? valid_0_25 : _GEN_10943; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11972 = 3'h4 == state ? valid_0_26 : _GEN_10944; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11973 = 3'h4 == state ? valid_0_27 : _GEN_10945; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11974 = 3'h4 == state ? valid_0_28 : _GEN_10946; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11975 = 3'h4 == state ? valid_0_29 : _GEN_10947; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11976 = 3'h4 == state ? valid_0_30 : _GEN_10948; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11977 = 3'h4 == state ? valid_0_31 : _GEN_10949; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11978 = 3'h4 == state ? valid_0_32 : _GEN_10950; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11979 = 3'h4 == state ? valid_0_33 : _GEN_10951; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11980 = 3'h4 == state ? valid_0_34 : _GEN_10952; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11981 = 3'h4 == state ? valid_0_35 : _GEN_10953; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11982 = 3'h4 == state ? valid_0_36 : _GEN_10954; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11983 = 3'h4 == state ? valid_0_37 : _GEN_10955; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11984 = 3'h4 == state ? valid_0_38 : _GEN_10956; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11985 = 3'h4 == state ? valid_0_39 : _GEN_10957; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11986 = 3'h4 == state ? valid_0_40 : _GEN_10958; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11987 = 3'h4 == state ? valid_0_41 : _GEN_10959; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11988 = 3'h4 == state ? valid_0_42 : _GEN_10960; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11989 = 3'h4 == state ? valid_0_43 : _GEN_10961; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11990 = 3'h4 == state ? valid_0_44 : _GEN_10962; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11991 = 3'h4 == state ? valid_0_45 : _GEN_10963; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11992 = 3'h4 == state ? valid_0_46 : _GEN_10964; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11993 = 3'h4 == state ? valid_0_47 : _GEN_10965; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11994 = 3'h4 == state ? valid_0_48 : _GEN_10966; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11995 = 3'h4 == state ? valid_0_49 : _GEN_10967; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11996 = 3'h4 == state ? valid_0_50 : _GEN_10968; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11997 = 3'h4 == state ? valid_0_51 : _GEN_10969; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11998 = 3'h4 == state ? valid_0_52 : _GEN_10970; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_11999 = 3'h4 == state ? valid_0_53 : _GEN_10971; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12000 = 3'h4 == state ? valid_0_54 : _GEN_10972; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12001 = 3'h4 == state ? valid_0_55 : _GEN_10973; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12002 = 3'h4 == state ? valid_0_56 : _GEN_10974; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12003 = 3'h4 == state ? valid_0_57 : _GEN_10975; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12004 = 3'h4 == state ? valid_0_58 : _GEN_10976; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12005 = 3'h4 == state ? valid_0_59 : _GEN_10977; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12006 = 3'h4 == state ? valid_0_60 : _GEN_10978; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12007 = 3'h4 == state ? valid_0_61 : _GEN_10979; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12008 = 3'h4 == state ? valid_0_62 : _GEN_10980; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12009 = 3'h4 == state ? valid_0_63 : _GEN_10981; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12010 = 3'h4 == state ? valid_0_64 : _GEN_10982; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12011 = 3'h4 == state ? valid_0_65 : _GEN_10983; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12012 = 3'h4 == state ? valid_0_66 : _GEN_10984; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12013 = 3'h4 == state ? valid_0_67 : _GEN_10985; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12014 = 3'h4 == state ? valid_0_68 : _GEN_10986; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12015 = 3'h4 == state ? valid_0_69 : _GEN_10987; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12016 = 3'h4 == state ? valid_0_70 : _GEN_10988; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12017 = 3'h4 == state ? valid_0_71 : _GEN_10989; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12018 = 3'h4 == state ? valid_0_72 : _GEN_10990; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12019 = 3'h4 == state ? valid_0_73 : _GEN_10991; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12020 = 3'h4 == state ? valid_0_74 : _GEN_10992; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12021 = 3'h4 == state ? valid_0_75 : _GEN_10993; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12022 = 3'h4 == state ? valid_0_76 : _GEN_10994; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12023 = 3'h4 == state ? valid_0_77 : _GEN_10995; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12024 = 3'h4 == state ? valid_0_78 : _GEN_10996; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12025 = 3'h4 == state ? valid_0_79 : _GEN_10997; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12026 = 3'h4 == state ? valid_0_80 : _GEN_10998; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12027 = 3'h4 == state ? valid_0_81 : _GEN_10999; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12028 = 3'h4 == state ? valid_0_82 : _GEN_11000; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12029 = 3'h4 == state ? valid_0_83 : _GEN_11001; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12030 = 3'h4 == state ? valid_0_84 : _GEN_11002; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12031 = 3'h4 == state ? valid_0_85 : _GEN_11003; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12032 = 3'h4 == state ? valid_0_86 : _GEN_11004; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12033 = 3'h4 == state ? valid_0_87 : _GEN_11005; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12034 = 3'h4 == state ? valid_0_88 : _GEN_11006; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12035 = 3'h4 == state ? valid_0_89 : _GEN_11007; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12036 = 3'h4 == state ? valid_0_90 : _GEN_11008; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12037 = 3'h4 == state ? valid_0_91 : _GEN_11009; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12038 = 3'h4 == state ? valid_0_92 : _GEN_11010; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12039 = 3'h4 == state ? valid_0_93 : _GEN_11011; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12040 = 3'h4 == state ? valid_0_94 : _GEN_11012; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12041 = 3'h4 == state ? valid_0_95 : _GEN_11013; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12042 = 3'h4 == state ? valid_0_96 : _GEN_11014; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12043 = 3'h4 == state ? valid_0_97 : _GEN_11015; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12044 = 3'h4 == state ? valid_0_98 : _GEN_11016; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12045 = 3'h4 == state ? valid_0_99 : _GEN_11017; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12046 = 3'h4 == state ? valid_0_100 : _GEN_11018; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12047 = 3'h4 == state ? valid_0_101 : _GEN_11019; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12048 = 3'h4 == state ? valid_0_102 : _GEN_11020; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12049 = 3'h4 == state ? valid_0_103 : _GEN_11021; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12050 = 3'h4 == state ? valid_0_104 : _GEN_11022; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12051 = 3'h4 == state ? valid_0_105 : _GEN_11023; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12052 = 3'h4 == state ? valid_0_106 : _GEN_11024; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12053 = 3'h4 == state ? valid_0_107 : _GEN_11025; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12054 = 3'h4 == state ? valid_0_108 : _GEN_11026; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12055 = 3'h4 == state ? valid_0_109 : _GEN_11027; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12056 = 3'h4 == state ? valid_0_110 : _GEN_11028; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12057 = 3'h4 == state ? valid_0_111 : _GEN_11029; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12058 = 3'h4 == state ? valid_0_112 : _GEN_11030; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12059 = 3'h4 == state ? valid_0_113 : _GEN_11031; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12060 = 3'h4 == state ? valid_0_114 : _GEN_11032; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12061 = 3'h4 == state ? valid_0_115 : _GEN_11033; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12062 = 3'h4 == state ? valid_0_116 : _GEN_11034; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12063 = 3'h4 == state ? valid_0_117 : _GEN_11035; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12064 = 3'h4 == state ? valid_0_118 : _GEN_11036; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12065 = 3'h4 == state ? valid_0_119 : _GEN_11037; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12066 = 3'h4 == state ? valid_0_120 : _GEN_11038; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12067 = 3'h4 == state ? valid_0_121 : _GEN_11039; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12068 = 3'h4 == state ? valid_0_122 : _GEN_11040; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12069 = 3'h4 == state ? valid_0_123 : _GEN_11041; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12070 = 3'h4 == state ? valid_0_124 : _GEN_11042; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12071 = 3'h4 == state ? valid_0_125 : _GEN_11043; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12072 = 3'h4 == state ? valid_0_126 : _GEN_11044; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12073 = 3'h4 == state ? valid_0_127 : _GEN_11045; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12074 = 3'h4 == state ? quene : _GEN_11046; // @[d_cache.scala 81:18 37:24]
  wire [63:0] _GEN_12075 = 3'h4 == state ? ram_1_0 : _GEN_11047; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12076 = 3'h4 == state ? ram_1_1 : _GEN_11048; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12077 = 3'h4 == state ? ram_1_2 : _GEN_11049; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12078 = 3'h4 == state ? ram_1_3 : _GEN_11050; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12079 = 3'h4 == state ? ram_1_4 : _GEN_11051; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12080 = 3'h4 == state ? ram_1_5 : _GEN_11052; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12081 = 3'h4 == state ? ram_1_6 : _GEN_11053; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12082 = 3'h4 == state ? ram_1_7 : _GEN_11054; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12083 = 3'h4 == state ? ram_1_8 : _GEN_11055; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12084 = 3'h4 == state ? ram_1_9 : _GEN_11056; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12085 = 3'h4 == state ? ram_1_10 : _GEN_11057; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12086 = 3'h4 == state ? ram_1_11 : _GEN_11058; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12087 = 3'h4 == state ? ram_1_12 : _GEN_11059; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12088 = 3'h4 == state ? ram_1_13 : _GEN_11060; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12089 = 3'h4 == state ? ram_1_14 : _GEN_11061; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12090 = 3'h4 == state ? ram_1_15 : _GEN_11062; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12091 = 3'h4 == state ? ram_1_16 : _GEN_11063; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12092 = 3'h4 == state ? ram_1_17 : _GEN_11064; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12093 = 3'h4 == state ? ram_1_18 : _GEN_11065; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12094 = 3'h4 == state ? ram_1_19 : _GEN_11066; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12095 = 3'h4 == state ? ram_1_20 : _GEN_11067; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12096 = 3'h4 == state ? ram_1_21 : _GEN_11068; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12097 = 3'h4 == state ? ram_1_22 : _GEN_11069; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12098 = 3'h4 == state ? ram_1_23 : _GEN_11070; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12099 = 3'h4 == state ? ram_1_24 : _GEN_11071; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12100 = 3'h4 == state ? ram_1_25 : _GEN_11072; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12101 = 3'h4 == state ? ram_1_26 : _GEN_11073; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12102 = 3'h4 == state ? ram_1_27 : _GEN_11074; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12103 = 3'h4 == state ? ram_1_28 : _GEN_11075; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12104 = 3'h4 == state ? ram_1_29 : _GEN_11076; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12105 = 3'h4 == state ? ram_1_30 : _GEN_11077; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12106 = 3'h4 == state ? ram_1_31 : _GEN_11078; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12107 = 3'h4 == state ? ram_1_32 : _GEN_11079; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12108 = 3'h4 == state ? ram_1_33 : _GEN_11080; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12109 = 3'h4 == state ? ram_1_34 : _GEN_11081; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12110 = 3'h4 == state ? ram_1_35 : _GEN_11082; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12111 = 3'h4 == state ? ram_1_36 : _GEN_11083; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12112 = 3'h4 == state ? ram_1_37 : _GEN_11084; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12113 = 3'h4 == state ? ram_1_38 : _GEN_11085; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12114 = 3'h4 == state ? ram_1_39 : _GEN_11086; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12115 = 3'h4 == state ? ram_1_40 : _GEN_11087; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12116 = 3'h4 == state ? ram_1_41 : _GEN_11088; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12117 = 3'h4 == state ? ram_1_42 : _GEN_11089; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12118 = 3'h4 == state ? ram_1_43 : _GEN_11090; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12119 = 3'h4 == state ? ram_1_44 : _GEN_11091; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12120 = 3'h4 == state ? ram_1_45 : _GEN_11092; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12121 = 3'h4 == state ? ram_1_46 : _GEN_11093; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12122 = 3'h4 == state ? ram_1_47 : _GEN_11094; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12123 = 3'h4 == state ? ram_1_48 : _GEN_11095; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12124 = 3'h4 == state ? ram_1_49 : _GEN_11096; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12125 = 3'h4 == state ? ram_1_50 : _GEN_11097; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12126 = 3'h4 == state ? ram_1_51 : _GEN_11098; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12127 = 3'h4 == state ? ram_1_52 : _GEN_11099; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12128 = 3'h4 == state ? ram_1_53 : _GEN_11100; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12129 = 3'h4 == state ? ram_1_54 : _GEN_11101; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12130 = 3'h4 == state ? ram_1_55 : _GEN_11102; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12131 = 3'h4 == state ? ram_1_56 : _GEN_11103; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12132 = 3'h4 == state ? ram_1_57 : _GEN_11104; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12133 = 3'h4 == state ? ram_1_58 : _GEN_11105; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12134 = 3'h4 == state ? ram_1_59 : _GEN_11106; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12135 = 3'h4 == state ? ram_1_60 : _GEN_11107; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12136 = 3'h4 == state ? ram_1_61 : _GEN_11108; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12137 = 3'h4 == state ? ram_1_62 : _GEN_11109; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12138 = 3'h4 == state ? ram_1_63 : _GEN_11110; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12139 = 3'h4 == state ? ram_1_64 : _GEN_11111; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12140 = 3'h4 == state ? ram_1_65 : _GEN_11112; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12141 = 3'h4 == state ? ram_1_66 : _GEN_11113; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12142 = 3'h4 == state ? ram_1_67 : _GEN_11114; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12143 = 3'h4 == state ? ram_1_68 : _GEN_11115; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12144 = 3'h4 == state ? ram_1_69 : _GEN_11116; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12145 = 3'h4 == state ? ram_1_70 : _GEN_11117; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12146 = 3'h4 == state ? ram_1_71 : _GEN_11118; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12147 = 3'h4 == state ? ram_1_72 : _GEN_11119; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12148 = 3'h4 == state ? ram_1_73 : _GEN_11120; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12149 = 3'h4 == state ? ram_1_74 : _GEN_11121; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12150 = 3'h4 == state ? ram_1_75 : _GEN_11122; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12151 = 3'h4 == state ? ram_1_76 : _GEN_11123; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12152 = 3'h4 == state ? ram_1_77 : _GEN_11124; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12153 = 3'h4 == state ? ram_1_78 : _GEN_11125; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12154 = 3'h4 == state ? ram_1_79 : _GEN_11126; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12155 = 3'h4 == state ? ram_1_80 : _GEN_11127; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12156 = 3'h4 == state ? ram_1_81 : _GEN_11128; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12157 = 3'h4 == state ? ram_1_82 : _GEN_11129; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12158 = 3'h4 == state ? ram_1_83 : _GEN_11130; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12159 = 3'h4 == state ? ram_1_84 : _GEN_11131; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12160 = 3'h4 == state ? ram_1_85 : _GEN_11132; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12161 = 3'h4 == state ? ram_1_86 : _GEN_11133; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12162 = 3'h4 == state ? ram_1_87 : _GEN_11134; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12163 = 3'h4 == state ? ram_1_88 : _GEN_11135; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12164 = 3'h4 == state ? ram_1_89 : _GEN_11136; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12165 = 3'h4 == state ? ram_1_90 : _GEN_11137; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12166 = 3'h4 == state ? ram_1_91 : _GEN_11138; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12167 = 3'h4 == state ? ram_1_92 : _GEN_11139; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12168 = 3'h4 == state ? ram_1_93 : _GEN_11140; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12169 = 3'h4 == state ? ram_1_94 : _GEN_11141; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12170 = 3'h4 == state ? ram_1_95 : _GEN_11142; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12171 = 3'h4 == state ? ram_1_96 : _GEN_11143; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12172 = 3'h4 == state ? ram_1_97 : _GEN_11144; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12173 = 3'h4 == state ? ram_1_98 : _GEN_11145; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12174 = 3'h4 == state ? ram_1_99 : _GEN_11146; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12175 = 3'h4 == state ? ram_1_100 : _GEN_11147; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12176 = 3'h4 == state ? ram_1_101 : _GEN_11148; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12177 = 3'h4 == state ? ram_1_102 : _GEN_11149; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12178 = 3'h4 == state ? ram_1_103 : _GEN_11150; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12179 = 3'h4 == state ? ram_1_104 : _GEN_11151; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12180 = 3'h4 == state ? ram_1_105 : _GEN_11152; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12181 = 3'h4 == state ? ram_1_106 : _GEN_11153; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12182 = 3'h4 == state ? ram_1_107 : _GEN_11154; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12183 = 3'h4 == state ? ram_1_108 : _GEN_11155; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12184 = 3'h4 == state ? ram_1_109 : _GEN_11156; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12185 = 3'h4 == state ? ram_1_110 : _GEN_11157; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12186 = 3'h4 == state ? ram_1_111 : _GEN_11158; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12187 = 3'h4 == state ? ram_1_112 : _GEN_11159; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12188 = 3'h4 == state ? ram_1_113 : _GEN_11160; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12189 = 3'h4 == state ? ram_1_114 : _GEN_11161; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12190 = 3'h4 == state ? ram_1_115 : _GEN_11162; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12191 = 3'h4 == state ? ram_1_116 : _GEN_11163; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12192 = 3'h4 == state ? ram_1_117 : _GEN_11164; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12193 = 3'h4 == state ? ram_1_118 : _GEN_11165; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12194 = 3'h4 == state ? ram_1_119 : _GEN_11166; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12195 = 3'h4 == state ? ram_1_120 : _GEN_11167; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12196 = 3'h4 == state ? ram_1_121 : _GEN_11168; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12197 = 3'h4 == state ? ram_1_122 : _GEN_11169; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12198 = 3'h4 == state ? ram_1_123 : _GEN_11170; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12199 = 3'h4 == state ? ram_1_124 : _GEN_11171; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12200 = 3'h4 == state ? ram_1_125 : _GEN_11172; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12201 = 3'h4 == state ? ram_1_126 : _GEN_11173; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_12202 = 3'h4 == state ? ram_1_127 : _GEN_11174; // @[d_cache.scala 81:18 19:24]
  wire [31:0] _GEN_12203 = 3'h4 == state ? tag_1_0 : _GEN_11175; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12204 = 3'h4 == state ? tag_1_1 : _GEN_11176; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12205 = 3'h4 == state ? tag_1_2 : _GEN_11177; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12206 = 3'h4 == state ? tag_1_3 : _GEN_11178; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12207 = 3'h4 == state ? tag_1_4 : _GEN_11179; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12208 = 3'h4 == state ? tag_1_5 : _GEN_11180; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12209 = 3'h4 == state ? tag_1_6 : _GEN_11181; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12210 = 3'h4 == state ? tag_1_7 : _GEN_11182; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12211 = 3'h4 == state ? tag_1_8 : _GEN_11183; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12212 = 3'h4 == state ? tag_1_9 : _GEN_11184; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12213 = 3'h4 == state ? tag_1_10 : _GEN_11185; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12214 = 3'h4 == state ? tag_1_11 : _GEN_11186; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12215 = 3'h4 == state ? tag_1_12 : _GEN_11187; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12216 = 3'h4 == state ? tag_1_13 : _GEN_11188; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12217 = 3'h4 == state ? tag_1_14 : _GEN_11189; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12218 = 3'h4 == state ? tag_1_15 : _GEN_11190; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12219 = 3'h4 == state ? tag_1_16 : _GEN_11191; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12220 = 3'h4 == state ? tag_1_17 : _GEN_11192; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12221 = 3'h4 == state ? tag_1_18 : _GEN_11193; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12222 = 3'h4 == state ? tag_1_19 : _GEN_11194; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12223 = 3'h4 == state ? tag_1_20 : _GEN_11195; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12224 = 3'h4 == state ? tag_1_21 : _GEN_11196; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12225 = 3'h4 == state ? tag_1_22 : _GEN_11197; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12226 = 3'h4 == state ? tag_1_23 : _GEN_11198; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12227 = 3'h4 == state ? tag_1_24 : _GEN_11199; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12228 = 3'h4 == state ? tag_1_25 : _GEN_11200; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12229 = 3'h4 == state ? tag_1_26 : _GEN_11201; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12230 = 3'h4 == state ? tag_1_27 : _GEN_11202; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12231 = 3'h4 == state ? tag_1_28 : _GEN_11203; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12232 = 3'h4 == state ? tag_1_29 : _GEN_11204; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12233 = 3'h4 == state ? tag_1_30 : _GEN_11205; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12234 = 3'h4 == state ? tag_1_31 : _GEN_11206; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12235 = 3'h4 == state ? tag_1_32 : _GEN_11207; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12236 = 3'h4 == state ? tag_1_33 : _GEN_11208; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12237 = 3'h4 == state ? tag_1_34 : _GEN_11209; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12238 = 3'h4 == state ? tag_1_35 : _GEN_11210; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12239 = 3'h4 == state ? tag_1_36 : _GEN_11211; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12240 = 3'h4 == state ? tag_1_37 : _GEN_11212; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12241 = 3'h4 == state ? tag_1_38 : _GEN_11213; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12242 = 3'h4 == state ? tag_1_39 : _GEN_11214; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12243 = 3'h4 == state ? tag_1_40 : _GEN_11215; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12244 = 3'h4 == state ? tag_1_41 : _GEN_11216; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12245 = 3'h4 == state ? tag_1_42 : _GEN_11217; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12246 = 3'h4 == state ? tag_1_43 : _GEN_11218; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12247 = 3'h4 == state ? tag_1_44 : _GEN_11219; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12248 = 3'h4 == state ? tag_1_45 : _GEN_11220; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12249 = 3'h4 == state ? tag_1_46 : _GEN_11221; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12250 = 3'h4 == state ? tag_1_47 : _GEN_11222; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12251 = 3'h4 == state ? tag_1_48 : _GEN_11223; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12252 = 3'h4 == state ? tag_1_49 : _GEN_11224; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12253 = 3'h4 == state ? tag_1_50 : _GEN_11225; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12254 = 3'h4 == state ? tag_1_51 : _GEN_11226; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12255 = 3'h4 == state ? tag_1_52 : _GEN_11227; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12256 = 3'h4 == state ? tag_1_53 : _GEN_11228; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12257 = 3'h4 == state ? tag_1_54 : _GEN_11229; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12258 = 3'h4 == state ? tag_1_55 : _GEN_11230; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12259 = 3'h4 == state ? tag_1_56 : _GEN_11231; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12260 = 3'h4 == state ? tag_1_57 : _GEN_11232; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12261 = 3'h4 == state ? tag_1_58 : _GEN_11233; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12262 = 3'h4 == state ? tag_1_59 : _GEN_11234; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12263 = 3'h4 == state ? tag_1_60 : _GEN_11235; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12264 = 3'h4 == state ? tag_1_61 : _GEN_11236; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12265 = 3'h4 == state ? tag_1_62 : _GEN_11237; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12266 = 3'h4 == state ? tag_1_63 : _GEN_11238; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12267 = 3'h4 == state ? tag_1_64 : _GEN_11239; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12268 = 3'h4 == state ? tag_1_65 : _GEN_11240; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12269 = 3'h4 == state ? tag_1_66 : _GEN_11241; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12270 = 3'h4 == state ? tag_1_67 : _GEN_11242; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12271 = 3'h4 == state ? tag_1_68 : _GEN_11243; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12272 = 3'h4 == state ? tag_1_69 : _GEN_11244; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12273 = 3'h4 == state ? tag_1_70 : _GEN_11245; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12274 = 3'h4 == state ? tag_1_71 : _GEN_11246; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12275 = 3'h4 == state ? tag_1_72 : _GEN_11247; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12276 = 3'h4 == state ? tag_1_73 : _GEN_11248; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12277 = 3'h4 == state ? tag_1_74 : _GEN_11249; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12278 = 3'h4 == state ? tag_1_75 : _GEN_11250; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12279 = 3'h4 == state ? tag_1_76 : _GEN_11251; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12280 = 3'h4 == state ? tag_1_77 : _GEN_11252; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12281 = 3'h4 == state ? tag_1_78 : _GEN_11253; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12282 = 3'h4 == state ? tag_1_79 : _GEN_11254; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12283 = 3'h4 == state ? tag_1_80 : _GEN_11255; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12284 = 3'h4 == state ? tag_1_81 : _GEN_11256; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12285 = 3'h4 == state ? tag_1_82 : _GEN_11257; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12286 = 3'h4 == state ? tag_1_83 : _GEN_11258; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12287 = 3'h4 == state ? tag_1_84 : _GEN_11259; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12288 = 3'h4 == state ? tag_1_85 : _GEN_11260; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12289 = 3'h4 == state ? tag_1_86 : _GEN_11261; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12290 = 3'h4 == state ? tag_1_87 : _GEN_11262; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12291 = 3'h4 == state ? tag_1_88 : _GEN_11263; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12292 = 3'h4 == state ? tag_1_89 : _GEN_11264; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12293 = 3'h4 == state ? tag_1_90 : _GEN_11265; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12294 = 3'h4 == state ? tag_1_91 : _GEN_11266; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12295 = 3'h4 == state ? tag_1_92 : _GEN_11267; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12296 = 3'h4 == state ? tag_1_93 : _GEN_11268; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12297 = 3'h4 == state ? tag_1_94 : _GEN_11269; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12298 = 3'h4 == state ? tag_1_95 : _GEN_11270; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12299 = 3'h4 == state ? tag_1_96 : _GEN_11271; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12300 = 3'h4 == state ? tag_1_97 : _GEN_11272; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12301 = 3'h4 == state ? tag_1_98 : _GEN_11273; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12302 = 3'h4 == state ? tag_1_99 : _GEN_11274; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12303 = 3'h4 == state ? tag_1_100 : _GEN_11275; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12304 = 3'h4 == state ? tag_1_101 : _GEN_11276; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12305 = 3'h4 == state ? tag_1_102 : _GEN_11277; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12306 = 3'h4 == state ? tag_1_103 : _GEN_11278; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12307 = 3'h4 == state ? tag_1_104 : _GEN_11279; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12308 = 3'h4 == state ? tag_1_105 : _GEN_11280; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12309 = 3'h4 == state ? tag_1_106 : _GEN_11281; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12310 = 3'h4 == state ? tag_1_107 : _GEN_11282; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12311 = 3'h4 == state ? tag_1_108 : _GEN_11283; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12312 = 3'h4 == state ? tag_1_109 : _GEN_11284; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12313 = 3'h4 == state ? tag_1_110 : _GEN_11285; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12314 = 3'h4 == state ? tag_1_111 : _GEN_11286; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12315 = 3'h4 == state ? tag_1_112 : _GEN_11287; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12316 = 3'h4 == state ? tag_1_113 : _GEN_11288; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12317 = 3'h4 == state ? tag_1_114 : _GEN_11289; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12318 = 3'h4 == state ? tag_1_115 : _GEN_11290; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12319 = 3'h4 == state ? tag_1_116 : _GEN_11291; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12320 = 3'h4 == state ? tag_1_117 : _GEN_11292; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12321 = 3'h4 == state ? tag_1_118 : _GEN_11293; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12322 = 3'h4 == state ? tag_1_119 : _GEN_11294; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12323 = 3'h4 == state ? tag_1_120 : _GEN_11295; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12324 = 3'h4 == state ? tag_1_121 : _GEN_11296; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12325 = 3'h4 == state ? tag_1_122 : _GEN_11297; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12326 = 3'h4 == state ? tag_1_123 : _GEN_11298; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12327 = 3'h4 == state ? tag_1_124 : _GEN_11299; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12328 = 3'h4 == state ? tag_1_125 : _GEN_11300; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12329 = 3'h4 == state ? tag_1_126 : _GEN_11301; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_12330 = 3'h4 == state ? tag_1_127 : _GEN_11302; // @[d_cache.scala 81:18 23:24]
  wire  _GEN_12331 = 3'h4 == state ? valid_1_0 : _GEN_11303; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12332 = 3'h4 == state ? valid_1_1 : _GEN_11304; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12333 = 3'h4 == state ? valid_1_2 : _GEN_11305; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12334 = 3'h4 == state ? valid_1_3 : _GEN_11306; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12335 = 3'h4 == state ? valid_1_4 : _GEN_11307; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12336 = 3'h4 == state ? valid_1_5 : _GEN_11308; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12337 = 3'h4 == state ? valid_1_6 : _GEN_11309; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12338 = 3'h4 == state ? valid_1_7 : _GEN_11310; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12339 = 3'h4 == state ? valid_1_8 : _GEN_11311; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12340 = 3'h4 == state ? valid_1_9 : _GEN_11312; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12341 = 3'h4 == state ? valid_1_10 : _GEN_11313; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12342 = 3'h4 == state ? valid_1_11 : _GEN_11314; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12343 = 3'h4 == state ? valid_1_12 : _GEN_11315; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12344 = 3'h4 == state ? valid_1_13 : _GEN_11316; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12345 = 3'h4 == state ? valid_1_14 : _GEN_11317; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12346 = 3'h4 == state ? valid_1_15 : _GEN_11318; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12347 = 3'h4 == state ? valid_1_16 : _GEN_11319; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12348 = 3'h4 == state ? valid_1_17 : _GEN_11320; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12349 = 3'h4 == state ? valid_1_18 : _GEN_11321; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12350 = 3'h4 == state ? valid_1_19 : _GEN_11322; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12351 = 3'h4 == state ? valid_1_20 : _GEN_11323; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12352 = 3'h4 == state ? valid_1_21 : _GEN_11324; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12353 = 3'h4 == state ? valid_1_22 : _GEN_11325; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12354 = 3'h4 == state ? valid_1_23 : _GEN_11326; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12355 = 3'h4 == state ? valid_1_24 : _GEN_11327; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12356 = 3'h4 == state ? valid_1_25 : _GEN_11328; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12357 = 3'h4 == state ? valid_1_26 : _GEN_11329; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12358 = 3'h4 == state ? valid_1_27 : _GEN_11330; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12359 = 3'h4 == state ? valid_1_28 : _GEN_11331; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12360 = 3'h4 == state ? valid_1_29 : _GEN_11332; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12361 = 3'h4 == state ? valid_1_30 : _GEN_11333; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12362 = 3'h4 == state ? valid_1_31 : _GEN_11334; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12363 = 3'h4 == state ? valid_1_32 : _GEN_11335; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12364 = 3'h4 == state ? valid_1_33 : _GEN_11336; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12365 = 3'h4 == state ? valid_1_34 : _GEN_11337; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12366 = 3'h4 == state ? valid_1_35 : _GEN_11338; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12367 = 3'h4 == state ? valid_1_36 : _GEN_11339; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12368 = 3'h4 == state ? valid_1_37 : _GEN_11340; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12369 = 3'h4 == state ? valid_1_38 : _GEN_11341; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12370 = 3'h4 == state ? valid_1_39 : _GEN_11342; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12371 = 3'h4 == state ? valid_1_40 : _GEN_11343; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12372 = 3'h4 == state ? valid_1_41 : _GEN_11344; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12373 = 3'h4 == state ? valid_1_42 : _GEN_11345; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12374 = 3'h4 == state ? valid_1_43 : _GEN_11346; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12375 = 3'h4 == state ? valid_1_44 : _GEN_11347; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12376 = 3'h4 == state ? valid_1_45 : _GEN_11348; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12377 = 3'h4 == state ? valid_1_46 : _GEN_11349; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12378 = 3'h4 == state ? valid_1_47 : _GEN_11350; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12379 = 3'h4 == state ? valid_1_48 : _GEN_11351; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12380 = 3'h4 == state ? valid_1_49 : _GEN_11352; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12381 = 3'h4 == state ? valid_1_50 : _GEN_11353; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12382 = 3'h4 == state ? valid_1_51 : _GEN_11354; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12383 = 3'h4 == state ? valid_1_52 : _GEN_11355; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12384 = 3'h4 == state ? valid_1_53 : _GEN_11356; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12385 = 3'h4 == state ? valid_1_54 : _GEN_11357; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12386 = 3'h4 == state ? valid_1_55 : _GEN_11358; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12387 = 3'h4 == state ? valid_1_56 : _GEN_11359; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12388 = 3'h4 == state ? valid_1_57 : _GEN_11360; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12389 = 3'h4 == state ? valid_1_58 : _GEN_11361; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12390 = 3'h4 == state ? valid_1_59 : _GEN_11362; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12391 = 3'h4 == state ? valid_1_60 : _GEN_11363; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12392 = 3'h4 == state ? valid_1_61 : _GEN_11364; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12393 = 3'h4 == state ? valid_1_62 : _GEN_11365; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12394 = 3'h4 == state ? valid_1_63 : _GEN_11366; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12395 = 3'h4 == state ? valid_1_64 : _GEN_11367; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12396 = 3'h4 == state ? valid_1_65 : _GEN_11368; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12397 = 3'h4 == state ? valid_1_66 : _GEN_11369; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12398 = 3'h4 == state ? valid_1_67 : _GEN_11370; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12399 = 3'h4 == state ? valid_1_68 : _GEN_11371; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12400 = 3'h4 == state ? valid_1_69 : _GEN_11372; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12401 = 3'h4 == state ? valid_1_70 : _GEN_11373; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12402 = 3'h4 == state ? valid_1_71 : _GEN_11374; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12403 = 3'h4 == state ? valid_1_72 : _GEN_11375; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12404 = 3'h4 == state ? valid_1_73 : _GEN_11376; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12405 = 3'h4 == state ? valid_1_74 : _GEN_11377; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12406 = 3'h4 == state ? valid_1_75 : _GEN_11378; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12407 = 3'h4 == state ? valid_1_76 : _GEN_11379; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12408 = 3'h4 == state ? valid_1_77 : _GEN_11380; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12409 = 3'h4 == state ? valid_1_78 : _GEN_11381; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12410 = 3'h4 == state ? valid_1_79 : _GEN_11382; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12411 = 3'h4 == state ? valid_1_80 : _GEN_11383; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12412 = 3'h4 == state ? valid_1_81 : _GEN_11384; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12413 = 3'h4 == state ? valid_1_82 : _GEN_11385; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12414 = 3'h4 == state ? valid_1_83 : _GEN_11386; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12415 = 3'h4 == state ? valid_1_84 : _GEN_11387; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12416 = 3'h4 == state ? valid_1_85 : _GEN_11388; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12417 = 3'h4 == state ? valid_1_86 : _GEN_11389; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12418 = 3'h4 == state ? valid_1_87 : _GEN_11390; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12419 = 3'h4 == state ? valid_1_88 : _GEN_11391; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12420 = 3'h4 == state ? valid_1_89 : _GEN_11392; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12421 = 3'h4 == state ? valid_1_90 : _GEN_11393; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12422 = 3'h4 == state ? valid_1_91 : _GEN_11394; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12423 = 3'h4 == state ? valid_1_92 : _GEN_11395; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12424 = 3'h4 == state ? valid_1_93 : _GEN_11396; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12425 = 3'h4 == state ? valid_1_94 : _GEN_11397; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12426 = 3'h4 == state ? valid_1_95 : _GEN_11398; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12427 = 3'h4 == state ? valid_1_96 : _GEN_11399; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12428 = 3'h4 == state ? valid_1_97 : _GEN_11400; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12429 = 3'h4 == state ? valid_1_98 : _GEN_11401; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12430 = 3'h4 == state ? valid_1_99 : _GEN_11402; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12431 = 3'h4 == state ? valid_1_100 : _GEN_11403; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12432 = 3'h4 == state ? valid_1_101 : _GEN_11404; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12433 = 3'h4 == state ? valid_1_102 : _GEN_11405; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12434 = 3'h4 == state ? valid_1_103 : _GEN_11406; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12435 = 3'h4 == state ? valid_1_104 : _GEN_11407; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12436 = 3'h4 == state ? valid_1_105 : _GEN_11408; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12437 = 3'h4 == state ? valid_1_106 : _GEN_11409; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12438 = 3'h4 == state ? valid_1_107 : _GEN_11410; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12439 = 3'h4 == state ? valid_1_108 : _GEN_11411; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12440 = 3'h4 == state ? valid_1_109 : _GEN_11412; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12441 = 3'h4 == state ? valid_1_110 : _GEN_11413; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12442 = 3'h4 == state ? valid_1_111 : _GEN_11414; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12443 = 3'h4 == state ? valid_1_112 : _GEN_11415; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12444 = 3'h4 == state ? valid_1_113 : _GEN_11416; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12445 = 3'h4 == state ? valid_1_114 : _GEN_11417; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12446 = 3'h4 == state ? valid_1_115 : _GEN_11418; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12447 = 3'h4 == state ? valid_1_116 : _GEN_11419; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12448 = 3'h4 == state ? valid_1_117 : _GEN_11420; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12449 = 3'h4 == state ? valid_1_118 : _GEN_11421; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12450 = 3'h4 == state ? valid_1_119 : _GEN_11422; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12451 = 3'h4 == state ? valid_1_120 : _GEN_11423; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12452 = 3'h4 == state ? valid_1_121 : _GEN_11424; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12453 = 3'h4 == state ? valid_1_122 : _GEN_11425; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12454 = 3'h4 == state ? valid_1_123 : _GEN_11426; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12455 = 3'h4 == state ? valid_1_124 : _GEN_11427; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12456 = 3'h4 == state ? valid_1_125 : _GEN_11428; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12457 = 3'h4 == state ? valid_1_126 : _GEN_11429; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_12458 = 3'h4 == state ? valid_1_127 : _GEN_11430; // @[d_cache.scala 81:18 25:26]
  wire [63:0] _GEN_12459 = 3'h4 == state ? write_back_data : _GEN_11431; // @[d_cache.scala 81:18 31:34]
  wire [41:0] _GEN_12460 = 3'h4 == state ? {{10'd0}, write_back_addr} : _GEN_11432; // @[d_cache.scala 81:18 32:34]
  wire  _GEN_12461 = 3'h4 == state ? dirty_0_0 : _GEN_11433; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12462 = 3'h4 == state ? dirty_0_1 : _GEN_11434; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12463 = 3'h4 == state ? dirty_0_2 : _GEN_11435; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12464 = 3'h4 == state ? dirty_0_3 : _GEN_11436; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12465 = 3'h4 == state ? dirty_0_4 : _GEN_11437; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12466 = 3'h4 == state ? dirty_0_5 : _GEN_11438; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12467 = 3'h4 == state ? dirty_0_6 : _GEN_11439; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12468 = 3'h4 == state ? dirty_0_7 : _GEN_11440; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12469 = 3'h4 == state ? dirty_0_8 : _GEN_11441; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12470 = 3'h4 == state ? dirty_0_9 : _GEN_11442; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12471 = 3'h4 == state ? dirty_0_10 : _GEN_11443; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12472 = 3'h4 == state ? dirty_0_11 : _GEN_11444; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12473 = 3'h4 == state ? dirty_0_12 : _GEN_11445; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12474 = 3'h4 == state ? dirty_0_13 : _GEN_11446; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12475 = 3'h4 == state ? dirty_0_14 : _GEN_11447; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12476 = 3'h4 == state ? dirty_0_15 : _GEN_11448; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12477 = 3'h4 == state ? dirty_0_16 : _GEN_11449; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12478 = 3'h4 == state ? dirty_0_17 : _GEN_11450; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12479 = 3'h4 == state ? dirty_0_18 : _GEN_11451; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12480 = 3'h4 == state ? dirty_0_19 : _GEN_11452; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12481 = 3'h4 == state ? dirty_0_20 : _GEN_11453; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12482 = 3'h4 == state ? dirty_0_21 : _GEN_11454; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12483 = 3'h4 == state ? dirty_0_22 : _GEN_11455; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12484 = 3'h4 == state ? dirty_0_23 : _GEN_11456; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12485 = 3'h4 == state ? dirty_0_24 : _GEN_11457; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12486 = 3'h4 == state ? dirty_0_25 : _GEN_11458; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12487 = 3'h4 == state ? dirty_0_26 : _GEN_11459; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12488 = 3'h4 == state ? dirty_0_27 : _GEN_11460; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12489 = 3'h4 == state ? dirty_0_28 : _GEN_11461; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12490 = 3'h4 == state ? dirty_0_29 : _GEN_11462; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12491 = 3'h4 == state ? dirty_0_30 : _GEN_11463; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12492 = 3'h4 == state ? dirty_0_31 : _GEN_11464; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12493 = 3'h4 == state ? dirty_0_32 : _GEN_11465; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12494 = 3'h4 == state ? dirty_0_33 : _GEN_11466; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12495 = 3'h4 == state ? dirty_0_34 : _GEN_11467; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12496 = 3'h4 == state ? dirty_0_35 : _GEN_11468; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12497 = 3'h4 == state ? dirty_0_36 : _GEN_11469; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12498 = 3'h4 == state ? dirty_0_37 : _GEN_11470; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12499 = 3'h4 == state ? dirty_0_38 : _GEN_11471; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12500 = 3'h4 == state ? dirty_0_39 : _GEN_11472; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12501 = 3'h4 == state ? dirty_0_40 : _GEN_11473; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12502 = 3'h4 == state ? dirty_0_41 : _GEN_11474; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12503 = 3'h4 == state ? dirty_0_42 : _GEN_11475; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12504 = 3'h4 == state ? dirty_0_43 : _GEN_11476; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12505 = 3'h4 == state ? dirty_0_44 : _GEN_11477; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12506 = 3'h4 == state ? dirty_0_45 : _GEN_11478; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12507 = 3'h4 == state ? dirty_0_46 : _GEN_11479; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12508 = 3'h4 == state ? dirty_0_47 : _GEN_11480; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12509 = 3'h4 == state ? dirty_0_48 : _GEN_11481; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12510 = 3'h4 == state ? dirty_0_49 : _GEN_11482; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12511 = 3'h4 == state ? dirty_0_50 : _GEN_11483; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12512 = 3'h4 == state ? dirty_0_51 : _GEN_11484; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12513 = 3'h4 == state ? dirty_0_52 : _GEN_11485; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12514 = 3'h4 == state ? dirty_0_53 : _GEN_11486; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12515 = 3'h4 == state ? dirty_0_54 : _GEN_11487; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12516 = 3'h4 == state ? dirty_0_55 : _GEN_11488; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12517 = 3'h4 == state ? dirty_0_56 : _GEN_11489; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12518 = 3'h4 == state ? dirty_0_57 : _GEN_11490; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12519 = 3'h4 == state ? dirty_0_58 : _GEN_11491; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12520 = 3'h4 == state ? dirty_0_59 : _GEN_11492; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12521 = 3'h4 == state ? dirty_0_60 : _GEN_11493; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12522 = 3'h4 == state ? dirty_0_61 : _GEN_11494; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12523 = 3'h4 == state ? dirty_0_62 : _GEN_11495; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12524 = 3'h4 == state ? dirty_0_63 : _GEN_11496; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12525 = 3'h4 == state ? dirty_0_64 : _GEN_11497; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12526 = 3'h4 == state ? dirty_0_65 : _GEN_11498; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12527 = 3'h4 == state ? dirty_0_66 : _GEN_11499; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12528 = 3'h4 == state ? dirty_0_67 : _GEN_11500; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12529 = 3'h4 == state ? dirty_0_68 : _GEN_11501; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12530 = 3'h4 == state ? dirty_0_69 : _GEN_11502; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12531 = 3'h4 == state ? dirty_0_70 : _GEN_11503; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12532 = 3'h4 == state ? dirty_0_71 : _GEN_11504; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12533 = 3'h4 == state ? dirty_0_72 : _GEN_11505; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12534 = 3'h4 == state ? dirty_0_73 : _GEN_11506; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12535 = 3'h4 == state ? dirty_0_74 : _GEN_11507; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12536 = 3'h4 == state ? dirty_0_75 : _GEN_11508; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12537 = 3'h4 == state ? dirty_0_76 : _GEN_11509; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12538 = 3'h4 == state ? dirty_0_77 : _GEN_11510; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12539 = 3'h4 == state ? dirty_0_78 : _GEN_11511; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12540 = 3'h4 == state ? dirty_0_79 : _GEN_11512; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12541 = 3'h4 == state ? dirty_0_80 : _GEN_11513; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12542 = 3'h4 == state ? dirty_0_81 : _GEN_11514; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12543 = 3'h4 == state ? dirty_0_82 : _GEN_11515; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12544 = 3'h4 == state ? dirty_0_83 : _GEN_11516; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12545 = 3'h4 == state ? dirty_0_84 : _GEN_11517; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12546 = 3'h4 == state ? dirty_0_85 : _GEN_11518; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12547 = 3'h4 == state ? dirty_0_86 : _GEN_11519; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12548 = 3'h4 == state ? dirty_0_87 : _GEN_11520; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12549 = 3'h4 == state ? dirty_0_88 : _GEN_11521; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12550 = 3'h4 == state ? dirty_0_89 : _GEN_11522; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12551 = 3'h4 == state ? dirty_0_90 : _GEN_11523; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12552 = 3'h4 == state ? dirty_0_91 : _GEN_11524; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12553 = 3'h4 == state ? dirty_0_92 : _GEN_11525; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12554 = 3'h4 == state ? dirty_0_93 : _GEN_11526; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12555 = 3'h4 == state ? dirty_0_94 : _GEN_11527; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12556 = 3'h4 == state ? dirty_0_95 : _GEN_11528; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12557 = 3'h4 == state ? dirty_0_96 : _GEN_11529; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12558 = 3'h4 == state ? dirty_0_97 : _GEN_11530; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12559 = 3'h4 == state ? dirty_0_98 : _GEN_11531; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12560 = 3'h4 == state ? dirty_0_99 : _GEN_11532; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12561 = 3'h4 == state ? dirty_0_100 : _GEN_11533; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12562 = 3'h4 == state ? dirty_0_101 : _GEN_11534; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12563 = 3'h4 == state ? dirty_0_102 : _GEN_11535; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12564 = 3'h4 == state ? dirty_0_103 : _GEN_11536; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12565 = 3'h4 == state ? dirty_0_104 : _GEN_11537; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12566 = 3'h4 == state ? dirty_0_105 : _GEN_11538; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12567 = 3'h4 == state ? dirty_0_106 : _GEN_11539; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12568 = 3'h4 == state ? dirty_0_107 : _GEN_11540; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12569 = 3'h4 == state ? dirty_0_108 : _GEN_11541; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12570 = 3'h4 == state ? dirty_0_109 : _GEN_11542; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12571 = 3'h4 == state ? dirty_0_110 : _GEN_11543; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12572 = 3'h4 == state ? dirty_0_111 : _GEN_11544; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12573 = 3'h4 == state ? dirty_0_112 : _GEN_11545; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12574 = 3'h4 == state ? dirty_0_113 : _GEN_11546; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12575 = 3'h4 == state ? dirty_0_114 : _GEN_11547; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12576 = 3'h4 == state ? dirty_0_115 : _GEN_11548; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12577 = 3'h4 == state ? dirty_0_116 : _GEN_11549; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12578 = 3'h4 == state ? dirty_0_117 : _GEN_11550; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12579 = 3'h4 == state ? dirty_0_118 : _GEN_11551; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12580 = 3'h4 == state ? dirty_0_119 : _GEN_11552; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12581 = 3'h4 == state ? dirty_0_120 : _GEN_11553; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12582 = 3'h4 == state ? dirty_0_121 : _GEN_11554; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12583 = 3'h4 == state ? dirty_0_122 : _GEN_11555; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12584 = 3'h4 == state ? dirty_0_123 : _GEN_11556; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12585 = 3'h4 == state ? dirty_0_124 : _GEN_11557; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12586 = 3'h4 == state ? dirty_0_125 : _GEN_11558; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12587 = 3'h4 == state ? dirty_0_126 : _GEN_11559; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12588 = 3'h4 == state ? dirty_0_127 : _GEN_11560; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_12589 = 3'h4 == state ? dirty_1_0 : _GEN_11561; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12590 = 3'h4 == state ? dirty_1_1 : _GEN_11562; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12591 = 3'h4 == state ? dirty_1_2 : _GEN_11563; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12592 = 3'h4 == state ? dirty_1_3 : _GEN_11564; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12593 = 3'h4 == state ? dirty_1_4 : _GEN_11565; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12594 = 3'h4 == state ? dirty_1_5 : _GEN_11566; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12595 = 3'h4 == state ? dirty_1_6 : _GEN_11567; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12596 = 3'h4 == state ? dirty_1_7 : _GEN_11568; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12597 = 3'h4 == state ? dirty_1_8 : _GEN_11569; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12598 = 3'h4 == state ? dirty_1_9 : _GEN_11570; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12599 = 3'h4 == state ? dirty_1_10 : _GEN_11571; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12600 = 3'h4 == state ? dirty_1_11 : _GEN_11572; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12601 = 3'h4 == state ? dirty_1_12 : _GEN_11573; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12602 = 3'h4 == state ? dirty_1_13 : _GEN_11574; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12603 = 3'h4 == state ? dirty_1_14 : _GEN_11575; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12604 = 3'h4 == state ? dirty_1_15 : _GEN_11576; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12605 = 3'h4 == state ? dirty_1_16 : _GEN_11577; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12606 = 3'h4 == state ? dirty_1_17 : _GEN_11578; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12607 = 3'h4 == state ? dirty_1_18 : _GEN_11579; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12608 = 3'h4 == state ? dirty_1_19 : _GEN_11580; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12609 = 3'h4 == state ? dirty_1_20 : _GEN_11581; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12610 = 3'h4 == state ? dirty_1_21 : _GEN_11582; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12611 = 3'h4 == state ? dirty_1_22 : _GEN_11583; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12612 = 3'h4 == state ? dirty_1_23 : _GEN_11584; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12613 = 3'h4 == state ? dirty_1_24 : _GEN_11585; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12614 = 3'h4 == state ? dirty_1_25 : _GEN_11586; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12615 = 3'h4 == state ? dirty_1_26 : _GEN_11587; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12616 = 3'h4 == state ? dirty_1_27 : _GEN_11588; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12617 = 3'h4 == state ? dirty_1_28 : _GEN_11589; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12618 = 3'h4 == state ? dirty_1_29 : _GEN_11590; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12619 = 3'h4 == state ? dirty_1_30 : _GEN_11591; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12620 = 3'h4 == state ? dirty_1_31 : _GEN_11592; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12621 = 3'h4 == state ? dirty_1_32 : _GEN_11593; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12622 = 3'h4 == state ? dirty_1_33 : _GEN_11594; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12623 = 3'h4 == state ? dirty_1_34 : _GEN_11595; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12624 = 3'h4 == state ? dirty_1_35 : _GEN_11596; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12625 = 3'h4 == state ? dirty_1_36 : _GEN_11597; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12626 = 3'h4 == state ? dirty_1_37 : _GEN_11598; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12627 = 3'h4 == state ? dirty_1_38 : _GEN_11599; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12628 = 3'h4 == state ? dirty_1_39 : _GEN_11600; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12629 = 3'h4 == state ? dirty_1_40 : _GEN_11601; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12630 = 3'h4 == state ? dirty_1_41 : _GEN_11602; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12631 = 3'h4 == state ? dirty_1_42 : _GEN_11603; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12632 = 3'h4 == state ? dirty_1_43 : _GEN_11604; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12633 = 3'h4 == state ? dirty_1_44 : _GEN_11605; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12634 = 3'h4 == state ? dirty_1_45 : _GEN_11606; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12635 = 3'h4 == state ? dirty_1_46 : _GEN_11607; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12636 = 3'h4 == state ? dirty_1_47 : _GEN_11608; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12637 = 3'h4 == state ? dirty_1_48 : _GEN_11609; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12638 = 3'h4 == state ? dirty_1_49 : _GEN_11610; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12639 = 3'h4 == state ? dirty_1_50 : _GEN_11611; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12640 = 3'h4 == state ? dirty_1_51 : _GEN_11612; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12641 = 3'h4 == state ? dirty_1_52 : _GEN_11613; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12642 = 3'h4 == state ? dirty_1_53 : _GEN_11614; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12643 = 3'h4 == state ? dirty_1_54 : _GEN_11615; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12644 = 3'h4 == state ? dirty_1_55 : _GEN_11616; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12645 = 3'h4 == state ? dirty_1_56 : _GEN_11617; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12646 = 3'h4 == state ? dirty_1_57 : _GEN_11618; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12647 = 3'h4 == state ? dirty_1_58 : _GEN_11619; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12648 = 3'h4 == state ? dirty_1_59 : _GEN_11620; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12649 = 3'h4 == state ? dirty_1_60 : _GEN_11621; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12650 = 3'h4 == state ? dirty_1_61 : _GEN_11622; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12651 = 3'h4 == state ? dirty_1_62 : _GEN_11623; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12652 = 3'h4 == state ? dirty_1_63 : _GEN_11624; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12653 = 3'h4 == state ? dirty_1_64 : _GEN_11625; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12654 = 3'h4 == state ? dirty_1_65 : _GEN_11626; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12655 = 3'h4 == state ? dirty_1_66 : _GEN_11627; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12656 = 3'h4 == state ? dirty_1_67 : _GEN_11628; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12657 = 3'h4 == state ? dirty_1_68 : _GEN_11629; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12658 = 3'h4 == state ? dirty_1_69 : _GEN_11630; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12659 = 3'h4 == state ? dirty_1_70 : _GEN_11631; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12660 = 3'h4 == state ? dirty_1_71 : _GEN_11632; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12661 = 3'h4 == state ? dirty_1_72 : _GEN_11633; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12662 = 3'h4 == state ? dirty_1_73 : _GEN_11634; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12663 = 3'h4 == state ? dirty_1_74 : _GEN_11635; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12664 = 3'h4 == state ? dirty_1_75 : _GEN_11636; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12665 = 3'h4 == state ? dirty_1_76 : _GEN_11637; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12666 = 3'h4 == state ? dirty_1_77 : _GEN_11638; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12667 = 3'h4 == state ? dirty_1_78 : _GEN_11639; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12668 = 3'h4 == state ? dirty_1_79 : _GEN_11640; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12669 = 3'h4 == state ? dirty_1_80 : _GEN_11641; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12670 = 3'h4 == state ? dirty_1_81 : _GEN_11642; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12671 = 3'h4 == state ? dirty_1_82 : _GEN_11643; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12672 = 3'h4 == state ? dirty_1_83 : _GEN_11644; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12673 = 3'h4 == state ? dirty_1_84 : _GEN_11645; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12674 = 3'h4 == state ? dirty_1_85 : _GEN_11646; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12675 = 3'h4 == state ? dirty_1_86 : _GEN_11647; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12676 = 3'h4 == state ? dirty_1_87 : _GEN_11648; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12677 = 3'h4 == state ? dirty_1_88 : _GEN_11649; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12678 = 3'h4 == state ? dirty_1_89 : _GEN_11650; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12679 = 3'h4 == state ? dirty_1_90 : _GEN_11651; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12680 = 3'h4 == state ? dirty_1_91 : _GEN_11652; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12681 = 3'h4 == state ? dirty_1_92 : _GEN_11653; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12682 = 3'h4 == state ? dirty_1_93 : _GEN_11654; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12683 = 3'h4 == state ? dirty_1_94 : _GEN_11655; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12684 = 3'h4 == state ? dirty_1_95 : _GEN_11656; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12685 = 3'h4 == state ? dirty_1_96 : _GEN_11657; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12686 = 3'h4 == state ? dirty_1_97 : _GEN_11658; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12687 = 3'h4 == state ? dirty_1_98 : _GEN_11659; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12688 = 3'h4 == state ? dirty_1_99 : _GEN_11660; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12689 = 3'h4 == state ? dirty_1_100 : _GEN_11661; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12690 = 3'h4 == state ? dirty_1_101 : _GEN_11662; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12691 = 3'h4 == state ? dirty_1_102 : _GEN_11663; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12692 = 3'h4 == state ? dirty_1_103 : _GEN_11664; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12693 = 3'h4 == state ? dirty_1_104 : _GEN_11665; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12694 = 3'h4 == state ? dirty_1_105 : _GEN_11666; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12695 = 3'h4 == state ? dirty_1_106 : _GEN_11667; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12696 = 3'h4 == state ? dirty_1_107 : _GEN_11668; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12697 = 3'h4 == state ? dirty_1_108 : _GEN_11669; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12698 = 3'h4 == state ? dirty_1_109 : _GEN_11670; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12699 = 3'h4 == state ? dirty_1_110 : _GEN_11671; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12700 = 3'h4 == state ? dirty_1_111 : _GEN_11672; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12701 = 3'h4 == state ? dirty_1_112 : _GEN_11673; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12702 = 3'h4 == state ? dirty_1_113 : _GEN_11674; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12703 = 3'h4 == state ? dirty_1_114 : _GEN_11675; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12704 = 3'h4 == state ? dirty_1_115 : _GEN_11676; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12705 = 3'h4 == state ? dirty_1_116 : _GEN_11677; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12706 = 3'h4 == state ? dirty_1_117 : _GEN_11678; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12707 = 3'h4 == state ? dirty_1_118 : _GEN_11679; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12708 = 3'h4 == state ? dirty_1_119 : _GEN_11680; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12709 = 3'h4 == state ? dirty_1_120 : _GEN_11681; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12710 = 3'h4 == state ? dirty_1_121 : _GEN_11682; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12711 = 3'h4 == state ? dirty_1_122 : _GEN_11683; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12712 = 3'h4 == state ? dirty_1_123 : _GEN_11684; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12713 = 3'h4 == state ? dirty_1_124 : _GEN_11685; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12714 = 3'h4 == state ? dirty_1_125 : _GEN_11686; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12715 = 3'h4 == state ? dirty_1_126 : _GEN_11687; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_12716 = 3'h4 == state ? dirty_1_127 : _GEN_11688; // @[d_cache.scala 81:18 27:26]
  wire [2:0] _GEN_12717 = 3'h3 == state ? _GEN_3211 : _GEN_11689; // @[d_cache.scala 81:18]
  wire [63:0] _GEN_12718 = 3'h3 == state ? _GEN_3212 : receive_data; // @[d_cache.scala 81:18 36:31]
  wire [63:0] _GEN_12719 = 3'h3 == state ? ram_0_0 : _GEN_11690; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12720 = 3'h3 == state ? ram_0_1 : _GEN_11691; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12721 = 3'h3 == state ? ram_0_2 : _GEN_11692; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12722 = 3'h3 == state ? ram_0_3 : _GEN_11693; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12723 = 3'h3 == state ? ram_0_4 : _GEN_11694; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12724 = 3'h3 == state ? ram_0_5 : _GEN_11695; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12725 = 3'h3 == state ? ram_0_6 : _GEN_11696; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12726 = 3'h3 == state ? ram_0_7 : _GEN_11697; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12727 = 3'h3 == state ? ram_0_8 : _GEN_11698; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12728 = 3'h3 == state ? ram_0_9 : _GEN_11699; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12729 = 3'h3 == state ? ram_0_10 : _GEN_11700; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12730 = 3'h3 == state ? ram_0_11 : _GEN_11701; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12731 = 3'h3 == state ? ram_0_12 : _GEN_11702; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12732 = 3'h3 == state ? ram_0_13 : _GEN_11703; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12733 = 3'h3 == state ? ram_0_14 : _GEN_11704; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12734 = 3'h3 == state ? ram_0_15 : _GEN_11705; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12735 = 3'h3 == state ? ram_0_16 : _GEN_11706; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12736 = 3'h3 == state ? ram_0_17 : _GEN_11707; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12737 = 3'h3 == state ? ram_0_18 : _GEN_11708; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12738 = 3'h3 == state ? ram_0_19 : _GEN_11709; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12739 = 3'h3 == state ? ram_0_20 : _GEN_11710; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12740 = 3'h3 == state ? ram_0_21 : _GEN_11711; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12741 = 3'h3 == state ? ram_0_22 : _GEN_11712; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12742 = 3'h3 == state ? ram_0_23 : _GEN_11713; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12743 = 3'h3 == state ? ram_0_24 : _GEN_11714; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12744 = 3'h3 == state ? ram_0_25 : _GEN_11715; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12745 = 3'h3 == state ? ram_0_26 : _GEN_11716; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12746 = 3'h3 == state ? ram_0_27 : _GEN_11717; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12747 = 3'h3 == state ? ram_0_28 : _GEN_11718; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12748 = 3'h3 == state ? ram_0_29 : _GEN_11719; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12749 = 3'h3 == state ? ram_0_30 : _GEN_11720; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12750 = 3'h3 == state ? ram_0_31 : _GEN_11721; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12751 = 3'h3 == state ? ram_0_32 : _GEN_11722; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12752 = 3'h3 == state ? ram_0_33 : _GEN_11723; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12753 = 3'h3 == state ? ram_0_34 : _GEN_11724; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12754 = 3'h3 == state ? ram_0_35 : _GEN_11725; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12755 = 3'h3 == state ? ram_0_36 : _GEN_11726; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12756 = 3'h3 == state ? ram_0_37 : _GEN_11727; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12757 = 3'h3 == state ? ram_0_38 : _GEN_11728; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12758 = 3'h3 == state ? ram_0_39 : _GEN_11729; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12759 = 3'h3 == state ? ram_0_40 : _GEN_11730; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12760 = 3'h3 == state ? ram_0_41 : _GEN_11731; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12761 = 3'h3 == state ? ram_0_42 : _GEN_11732; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12762 = 3'h3 == state ? ram_0_43 : _GEN_11733; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12763 = 3'h3 == state ? ram_0_44 : _GEN_11734; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12764 = 3'h3 == state ? ram_0_45 : _GEN_11735; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12765 = 3'h3 == state ? ram_0_46 : _GEN_11736; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12766 = 3'h3 == state ? ram_0_47 : _GEN_11737; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12767 = 3'h3 == state ? ram_0_48 : _GEN_11738; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12768 = 3'h3 == state ? ram_0_49 : _GEN_11739; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12769 = 3'h3 == state ? ram_0_50 : _GEN_11740; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12770 = 3'h3 == state ? ram_0_51 : _GEN_11741; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12771 = 3'h3 == state ? ram_0_52 : _GEN_11742; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12772 = 3'h3 == state ? ram_0_53 : _GEN_11743; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12773 = 3'h3 == state ? ram_0_54 : _GEN_11744; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12774 = 3'h3 == state ? ram_0_55 : _GEN_11745; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12775 = 3'h3 == state ? ram_0_56 : _GEN_11746; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12776 = 3'h3 == state ? ram_0_57 : _GEN_11747; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12777 = 3'h3 == state ? ram_0_58 : _GEN_11748; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12778 = 3'h3 == state ? ram_0_59 : _GEN_11749; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12779 = 3'h3 == state ? ram_0_60 : _GEN_11750; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12780 = 3'h3 == state ? ram_0_61 : _GEN_11751; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12781 = 3'h3 == state ? ram_0_62 : _GEN_11752; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12782 = 3'h3 == state ? ram_0_63 : _GEN_11753; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12783 = 3'h3 == state ? ram_0_64 : _GEN_11754; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12784 = 3'h3 == state ? ram_0_65 : _GEN_11755; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12785 = 3'h3 == state ? ram_0_66 : _GEN_11756; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12786 = 3'h3 == state ? ram_0_67 : _GEN_11757; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12787 = 3'h3 == state ? ram_0_68 : _GEN_11758; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12788 = 3'h3 == state ? ram_0_69 : _GEN_11759; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12789 = 3'h3 == state ? ram_0_70 : _GEN_11760; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12790 = 3'h3 == state ? ram_0_71 : _GEN_11761; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12791 = 3'h3 == state ? ram_0_72 : _GEN_11762; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12792 = 3'h3 == state ? ram_0_73 : _GEN_11763; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12793 = 3'h3 == state ? ram_0_74 : _GEN_11764; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12794 = 3'h3 == state ? ram_0_75 : _GEN_11765; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12795 = 3'h3 == state ? ram_0_76 : _GEN_11766; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12796 = 3'h3 == state ? ram_0_77 : _GEN_11767; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12797 = 3'h3 == state ? ram_0_78 : _GEN_11768; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12798 = 3'h3 == state ? ram_0_79 : _GEN_11769; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12799 = 3'h3 == state ? ram_0_80 : _GEN_11770; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12800 = 3'h3 == state ? ram_0_81 : _GEN_11771; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12801 = 3'h3 == state ? ram_0_82 : _GEN_11772; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12802 = 3'h3 == state ? ram_0_83 : _GEN_11773; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12803 = 3'h3 == state ? ram_0_84 : _GEN_11774; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12804 = 3'h3 == state ? ram_0_85 : _GEN_11775; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12805 = 3'h3 == state ? ram_0_86 : _GEN_11776; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12806 = 3'h3 == state ? ram_0_87 : _GEN_11777; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12807 = 3'h3 == state ? ram_0_88 : _GEN_11778; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12808 = 3'h3 == state ? ram_0_89 : _GEN_11779; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12809 = 3'h3 == state ? ram_0_90 : _GEN_11780; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12810 = 3'h3 == state ? ram_0_91 : _GEN_11781; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12811 = 3'h3 == state ? ram_0_92 : _GEN_11782; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12812 = 3'h3 == state ? ram_0_93 : _GEN_11783; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12813 = 3'h3 == state ? ram_0_94 : _GEN_11784; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12814 = 3'h3 == state ? ram_0_95 : _GEN_11785; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12815 = 3'h3 == state ? ram_0_96 : _GEN_11786; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12816 = 3'h3 == state ? ram_0_97 : _GEN_11787; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12817 = 3'h3 == state ? ram_0_98 : _GEN_11788; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12818 = 3'h3 == state ? ram_0_99 : _GEN_11789; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12819 = 3'h3 == state ? ram_0_100 : _GEN_11790; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12820 = 3'h3 == state ? ram_0_101 : _GEN_11791; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12821 = 3'h3 == state ? ram_0_102 : _GEN_11792; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12822 = 3'h3 == state ? ram_0_103 : _GEN_11793; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12823 = 3'h3 == state ? ram_0_104 : _GEN_11794; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12824 = 3'h3 == state ? ram_0_105 : _GEN_11795; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12825 = 3'h3 == state ? ram_0_106 : _GEN_11796; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12826 = 3'h3 == state ? ram_0_107 : _GEN_11797; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12827 = 3'h3 == state ? ram_0_108 : _GEN_11798; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12828 = 3'h3 == state ? ram_0_109 : _GEN_11799; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12829 = 3'h3 == state ? ram_0_110 : _GEN_11800; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12830 = 3'h3 == state ? ram_0_111 : _GEN_11801; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12831 = 3'h3 == state ? ram_0_112 : _GEN_11802; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12832 = 3'h3 == state ? ram_0_113 : _GEN_11803; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12833 = 3'h3 == state ? ram_0_114 : _GEN_11804; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12834 = 3'h3 == state ? ram_0_115 : _GEN_11805; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12835 = 3'h3 == state ? ram_0_116 : _GEN_11806; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12836 = 3'h3 == state ? ram_0_117 : _GEN_11807; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12837 = 3'h3 == state ? ram_0_118 : _GEN_11808; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12838 = 3'h3 == state ? ram_0_119 : _GEN_11809; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12839 = 3'h3 == state ? ram_0_120 : _GEN_11810; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12840 = 3'h3 == state ? ram_0_121 : _GEN_11811; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12841 = 3'h3 == state ? ram_0_122 : _GEN_11812; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12842 = 3'h3 == state ? ram_0_123 : _GEN_11813; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12843 = 3'h3 == state ? ram_0_124 : _GEN_11814; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12844 = 3'h3 == state ? ram_0_125 : _GEN_11815; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12845 = 3'h3 == state ? ram_0_126 : _GEN_11816; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_12846 = 3'h3 == state ? ram_0_127 : _GEN_11817; // @[d_cache.scala 81:18 18:24]
  wire [31:0] _GEN_12847 = 3'h3 == state ? tag_0_0 : _GEN_11818; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12848 = 3'h3 == state ? tag_0_1 : _GEN_11819; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12849 = 3'h3 == state ? tag_0_2 : _GEN_11820; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12850 = 3'h3 == state ? tag_0_3 : _GEN_11821; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12851 = 3'h3 == state ? tag_0_4 : _GEN_11822; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12852 = 3'h3 == state ? tag_0_5 : _GEN_11823; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12853 = 3'h3 == state ? tag_0_6 : _GEN_11824; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12854 = 3'h3 == state ? tag_0_7 : _GEN_11825; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12855 = 3'h3 == state ? tag_0_8 : _GEN_11826; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12856 = 3'h3 == state ? tag_0_9 : _GEN_11827; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12857 = 3'h3 == state ? tag_0_10 : _GEN_11828; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12858 = 3'h3 == state ? tag_0_11 : _GEN_11829; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12859 = 3'h3 == state ? tag_0_12 : _GEN_11830; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12860 = 3'h3 == state ? tag_0_13 : _GEN_11831; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12861 = 3'h3 == state ? tag_0_14 : _GEN_11832; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12862 = 3'h3 == state ? tag_0_15 : _GEN_11833; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12863 = 3'h3 == state ? tag_0_16 : _GEN_11834; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12864 = 3'h3 == state ? tag_0_17 : _GEN_11835; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12865 = 3'h3 == state ? tag_0_18 : _GEN_11836; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12866 = 3'h3 == state ? tag_0_19 : _GEN_11837; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12867 = 3'h3 == state ? tag_0_20 : _GEN_11838; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12868 = 3'h3 == state ? tag_0_21 : _GEN_11839; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12869 = 3'h3 == state ? tag_0_22 : _GEN_11840; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12870 = 3'h3 == state ? tag_0_23 : _GEN_11841; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12871 = 3'h3 == state ? tag_0_24 : _GEN_11842; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12872 = 3'h3 == state ? tag_0_25 : _GEN_11843; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12873 = 3'h3 == state ? tag_0_26 : _GEN_11844; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12874 = 3'h3 == state ? tag_0_27 : _GEN_11845; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12875 = 3'h3 == state ? tag_0_28 : _GEN_11846; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12876 = 3'h3 == state ? tag_0_29 : _GEN_11847; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12877 = 3'h3 == state ? tag_0_30 : _GEN_11848; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12878 = 3'h3 == state ? tag_0_31 : _GEN_11849; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12879 = 3'h3 == state ? tag_0_32 : _GEN_11850; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12880 = 3'h3 == state ? tag_0_33 : _GEN_11851; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12881 = 3'h3 == state ? tag_0_34 : _GEN_11852; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12882 = 3'h3 == state ? tag_0_35 : _GEN_11853; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12883 = 3'h3 == state ? tag_0_36 : _GEN_11854; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12884 = 3'h3 == state ? tag_0_37 : _GEN_11855; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12885 = 3'h3 == state ? tag_0_38 : _GEN_11856; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12886 = 3'h3 == state ? tag_0_39 : _GEN_11857; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12887 = 3'h3 == state ? tag_0_40 : _GEN_11858; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12888 = 3'h3 == state ? tag_0_41 : _GEN_11859; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12889 = 3'h3 == state ? tag_0_42 : _GEN_11860; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12890 = 3'h3 == state ? tag_0_43 : _GEN_11861; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12891 = 3'h3 == state ? tag_0_44 : _GEN_11862; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12892 = 3'h3 == state ? tag_0_45 : _GEN_11863; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12893 = 3'h3 == state ? tag_0_46 : _GEN_11864; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12894 = 3'h3 == state ? tag_0_47 : _GEN_11865; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12895 = 3'h3 == state ? tag_0_48 : _GEN_11866; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12896 = 3'h3 == state ? tag_0_49 : _GEN_11867; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12897 = 3'h3 == state ? tag_0_50 : _GEN_11868; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12898 = 3'h3 == state ? tag_0_51 : _GEN_11869; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12899 = 3'h3 == state ? tag_0_52 : _GEN_11870; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12900 = 3'h3 == state ? tag_0_53 : _GEN_11871; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12901 = 3'h3 == state ? tag_0_54 : _GEN_11872; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12902 = 3'h3 == state ? tag_0_55 : _GEN_11873; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12903 = 3'h3 == state ? tag_0_56 : _GEN_11874; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12904 = 3'h3 == state ? tag_0_57 : _GEN_11875; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12905 = 3'h3 == state ? tag_0_58 : _GEN_11876; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12906 = 3'h3 == state ? tag_0_59 : _GEN_11877; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12907 = 3'h3 == state ? tag_0_60 : _GEN_11878; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12908 = 3'h3 == state ? tag_0_61 : _GEN_11879; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12909 = 3'h3 == state ? tag_0_62 : _GEN_11880; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12910 = 3'h3 == state ? tag_0_63 : _GEN_11881; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12911 = 3'h3 == state ? tag_0_64 : _GEN_11882; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12912 = 3'h3 == state ? tag_0_65 : _GEN_11883; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12913 = 3'h3 == state ? tag_0_66 : _GEN_11884; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12914 = 3'h3 == state ? tag_0_67 : _GEN_11885; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12915 = 3'h3 == state ? tag_0_68 : _GEN_11886; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12916 = 3'h3 == state ? tag_0_69 : _GEN_11887; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12917 = 3'h3 == state ? tag_0_70 : _GEN_11888; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12918 = 3'h3 == state ? tag_0_71 : _GEN_11889; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12919 = 3'h3 == state ? tag_0_72 : _GEN_11890; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12920 = 3'h3 == state ? tag_0_73 : _GEN_11891; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12921 = 3'h3 == state ? tag_0_74 : _GEN_11892; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12922 = 3'h3 == state ? tag_0_75 : _GEN_11893; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12923 = 3'h3 == state ? tag_0_76 : _GEN_11894; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12924 = 3'h3 == state ? tag_0_77 : _GEN_11895; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12925 = 3'h3 == state ? tag_0_78 : _GEN_11896; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12926 = 3'h3 == state ? tag_0_79 : _GEN_11897; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12927 = 3'h3 == state ? tag_0_80 : _GEN_11898; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12928 = 3'h3 == state ? tag_0_81 : _GEN_11899; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12929 = 3'h3 == state ? tag_0_82 : _GEN_11900; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12930 = 3'h3 == state ? tag_0_83 : _GEN_11901; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12931 = 3'h3 == state ? tag_0_84 : _GEN_11902; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12932 = 3'h3 == state ? tag_0_85 : _GEN_11903; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12933 = 3'h3 == state ? tag_0_86 : _GEN_11904; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12934 = 3'h3 == state ? tag_0_87 : _GEN_11905; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12935 = 3'h3 == state ? tag_0_88 : _GEN_11906; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12936 = 3'h3 == state ? tag_0_89 : _GEN_11907; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12937 = 3'h3 == state ? tag_0_90 : _GEN_11908; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12938 = 3'h3 == state ? tag_0_91 : _GEN_11909; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12939 = 3'h3 == state ? tag_0_92 : _GEN_11910; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12940 = 3'h3 == state ? tag_0_93 : _GEN_11911; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12941 = 3'h3 == state ? tag_0_94 : _GEN_11912; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12942 = 3'h3 == state ? tag_0_95 : _GEN_11913; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12943 = 3'h3 == state ? tag_0_96 : _GEN_11914; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12944 = 3'h3 == state ? tag_0_97 : _GEN_11915; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12945 = 3'h3 == state ? tag_0_98 : _GEN_11916; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12946 = 3'h3 == state ? tag_0_99 : _GEN_11917; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12947 = 3'h3 == state ? tag_0_100 : _GEN_11918; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12948 = 3'h3 == state ? tag_0_101 : _GEN_11919; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12949 = 3'h3 == state ? tag_0_102 : _GEN_11920; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12950 = 3'h3 == state ? tag_0_103 : _GEN_11921; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12951 = 3'h3 == state ? tag_0_104 : _GEN_11922; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12952 = 3'h3 == state ? tag_0_105 : _GEN_11923; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12953 = 3'h3 == state ? tag_0_106 : _GEN_11924; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12954 = 3'h3 == state ? tag_0_107 : _GEN_11925; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12955 = 3'h3 == state ? tag_0_108 : _GEN_11926; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12956 = 3'h3 == state ? tag_0_109 : _GEN_11927; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12957 = 3'h3 == state ? tag_0_110 : _GEN_11928; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12958 = 3'h3 == state ? tag_0_111 : _GEN_11929; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12959 = 3'h3 == state ? tag_0_112 : _GEN_11930; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12960 = 3'h3 == state ? tag_0_113 : _GEN_11931; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12961 = 3'h3 == state ? tag_0_114 : _GEN_11932; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12962 = 3'h3 == state ? tag_0_115 : _GEN_11933; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12963 = 3'h3 == state ? tag_0_116 : _GEN_11934; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12964 = 3'h3 == state ? tag_0_117 : _GEN_11935; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12965 = 3'h3 == state ? tag_0_118 : _GEN_11936; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12966 = 3'h3 == state ? tag_0_119 : _GEN_11937; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12967 = 3'h3 == state ? tag_0_120 : _GEN_11938; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12968 = 3'h3 == state ? tag_0_121 : _GEN_11939; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12969 = 3'h3 == state ? tag_0_122 : _GEN_11940; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12970 = 3'h3 == state ? tag_0_123 : _GEN_11941; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12971 = 3'h3 == state ? tag_0_124 : _GEN_11942; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12972 = 3'h3 == state ? tag_0_125 : _GEN_11943; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12973 = 3'h3 == state ? tag_0_126 : _GEN_11944; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_12974 = 3'h3 == state ? tag_0_127 : _GEN_11945; // @[d_cache.scala 81:18 22:24]
  wire  _GEN_12975 = 3'h3 == state ? valid_0_0 : _GEN_11946; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12976 = 3'h3 == state ? valid_0_1 : _GEN_11947; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12977 = 3'h3 == state ? valid_0_2 : _GEN_11948; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12978 = 3'h3 == state ? valid_0_3 : _GEN_11949; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12979 = 3'h3 == state ? valid_0_4 : _GEN_11950; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12980 = 3'h3 == state ? valid_0_5 : _GEN_11951; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12981 = 3'h3 == state ? valid_0_6 : _GEN_11952; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12982 = 3'h3 == state ? valid_0_7 : _GEN_11953; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12983 = 3'h3 == state ? valid_0_8 : _GEN_11954; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12984 = 3'h3 == state ? valid_0_9 : _GEN_11955; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12985 = 3'h3 == state ? valid_0_10 : _GEN_11956; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12986 = 3'h3 == state ? valid_0_11 : _GEN_11957; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12987 = 3'h3 == state ? valid_0_12 : _GEN_11958; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12988 = 3'h3 == state ? valid_0_13 : _GEN_11959; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12989 = 3'h3 == state ? valid_0_14 : _GEN_11960; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12990 = 3'h3 == state ? valid_0_15 : _GEN_11961; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12991 = 3'h3 == state ? valid_0_16 : _GEN_11962; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12992 = 3'h3 == state ? valid_0_17 : _GEN_11963; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12993 = 3'h3 == state ? valid_0_18 : _GEN_11964; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12994 = 3'h3 == state ? valid_0_19 : _GEN_11965; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12995 = 3'h3 == state ? valid_0_20 : _GEN_11966; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12996 = 3'h3 == state ? valid_0_21 : _GEN_11967; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12997 = 3'h3 == state ? valid_0_22 : _GEN_11968; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12998 = 3'h3 == state ? valid_0_23 : _GEN_11969; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_12999 = 3'h3 == state ? valid_0_24 : _GEN_11970; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13000 = 3'h3 == state ? valid_0_25 : _GEN_11971; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13001 = 3'h3 == state ? valid_0_26 : _GEN_11972; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13002 = 3'h3 == state ? valid_0_27 : _GEN_11973; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13003 = 3'h3 == state ? valid_0_28 : _GEN_11974; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13004 = 3'h3 == state ? valid_0_29 : _GEN_11975; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13005 = 3'h3 == state ? valid_0_30 : _GEN_11976; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13006 = 3'h3 == state ? valid_0_31 : _GEN_11977; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13007 = 3'h3 == state ? valid_0_32 : _GEN_11978; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13008 = 3'h3 == state ? valid_0_33 : _GEN_11979; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13009 = 3'h3 == state ? valid_0_34 : _GEN_11980; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13010 = 3'h3 == state ? valid_0_35 : _GEN_11981; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13011 = 3'h3 == state ? valid_0_36 : _GEN_11982; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13012 = 3'h3 == state ? valid_0_37 : _GEN_11983; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13013 = 3'h3 == state ? valid_0_38 : _GEN_11984; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13014 = 3'h3 == state ? valid_0_39 : _GEN_11985; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13015 = 3'h3 == state ? valid_0_40 : _GEN_11986; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13016 = 3'h3 == state ? valid_0_41 : _GEN_11987; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13017 = 3'h3 == state ? valid_0_42 : _GEN_11988; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13018 = 3'h3 == state ? valid_0_43 : _GEN_11989; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13019 = 3'h3 == state ? valid_0_44 : _GEN_11990; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13020 = 3'h3 == state ? valid_0_45 : _GEN_11991; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13021 = 3'h3 == state ? valid_0_46 : _GEN_11992; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13022 = 3'h3 == state ? valid_0_47 : _GEN_11993; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13023 = 3'h3 == state ? valid_0_48 : _GEN_11994; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13024 = 3'h3 == state ? valid_0_49 : _GEN_11995; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13025 = 3'h3 == state ? valid_0_50 : _GEN_11996; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13026 = 3'h3 == state ? valid_0_51 : _GEN_11997; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13027 = 3'h3 == state ? valid_0_52 : _GEN_11998; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13028 = 3'h3 == state ? valid_0_53 : _GEN_11999; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13029 = 3'h3 == state ? valid_0_54 : _GEN_12000; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13030 = 3'h3 == state ? valid_0_55 : _GEN_12001; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13031 = 3'h3 == state ? valid_0_56 : _GEN_12002; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13032 = 3'h3 == state ? valid_0_57 : _GEN_12003; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13033 = 3'h3 == state ? valid_0_58 : _GEN_12004; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13034 = 3'h3 == state ? valid_0_59 : _GEN_12005; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13035 = 3'h3 == state ? valid_0_60 : _GEN_12006; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13036 = 3'h3 == state ? valid_0_61 : _GEN_12007; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13037 = 3'h3 == state ? valid_0_62 : _GEN_12008; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13038 = 3'h3 == state ? valid_0_63 : _GEN_12009; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13039 = 3'h3 == state ? valid_0_64 : _GEN_12010; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13040 = 3'h3 == state ? valid_0_65 : _GEN_12011; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13041 = 3'h3 == state ? valid_0_66 : _GEN_12012; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13042 = 3'h3 == state ? valid_0_67 : _GEN_12013; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13043 = 3'h3 == state ? valid_0_68 : _GEN_12014; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13044 = 3'h3 == state ? valid_0_69 : _GEN_12015; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13045 = 3'h3 == state ? valid_0_70 : _GEN_12016; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13046 = 3'h3 == state ? valid_0_71 : _GEN_12017; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13047 = 3'h3 == state ? valid_0_72 : _GEN_12018; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13048 = 3'h3 == state ? valid_0_73 : _GEN_12019; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13049 = 3'h3 == state ? valid_0_74 : _GEN_12020; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13050 = 3'h3 == state ? valid_0_75 : _GEN_12021; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13051 = 3'h3 == state ? valid_0_76 : _GEN_12022; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13052 = 3'h3 == state ? valid_0_77 : _GEN_12023; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13053 = 3'h3 == state ? valid_0_78 : _GEN_12024; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13054 = 3'h3 == state ? valid_0_79 : _GEN_12025; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13055 = 3'h3 == state ? valid_0_80 : _GEN_12026; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13056 = 3'h3 == state ? valid_0_81 : _GEN_12027; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13057 = 3'h3 == state ? valid_0_82 : _GEN_12028; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13058 = 3'h3 == state ? valid_0_83 : _GEN_12029; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13059 = 3'h3 == state ? valid_0_84 : _GEN_12030; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13060 = 3'h3 == state ? valid_0_85 : _GEN_12031; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13061 = 3'h3 == state ? valid_0_86 : _GEN_12032; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13062 = 3'h3 == state ? valid_0_87 : _GEN_12033; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13063 = 3'h3 == state ? valid_0_88 : _GEN_12034; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13064 = 3'h3 == state ? valid_0_89 : _GEN_12035; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13065 = 3'h3 == state ? valid_0_90 : _GEN_12036; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13066 = 3'h3 == state ? valid_0_91 : _GEN_12037; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13067 = 3'h3 == state ? valid_0_92 : _GEN_12038; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13068 = 3'h3 == state ? valid_0_93 : _GEN_12039; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13069 = 3'h3 == state ? valid_0_94 : _GEN_12040; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13070 = 3'h3 == state ? valid_0_95 : _GEN_12041; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13071 = 3'h3 == state ? valid_0_96 : _GEN_12042; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13072 = 3'h3 == state ? valid_0_97 : _GEN_12043; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13073 = 3'h3 == state ? valid_0_98 : _GEN_12044; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13074 = 3'h3 == state ? valid_0_99 : _GEN_12045; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13075 = 3'h3 == state ? valid_0_100 : _GEN_12046; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13076 = 3'h3 == state ? valid_0_101 : _GEN_12047; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13077 = 3'h3 == state ? valid_0_102 : _GEN_12048; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13078 = 3'h3 == state ? valid_0_103 : _GEN_12049; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13079 = 3'h3 == state ? valid_0_104 : _GEN_12050; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13080 = 3'h3 == state ? valid_0_105 : _GEN_12051; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13081 = 3'h3 == state ? valid_0_106 : _GEN_12052; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13082 = 3'h3 == state ? valid_0_107 : _GEN_12053; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13083 = 3'h3 == state ? valid_0_108 : _GEN_12054; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13084 = 3'h3 == state ? valid_0_109 : _GEN_12055; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13085 = 3'h3 == state ? valid_0_110 : _GEN_12056; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13086 = 3'h3 == state ? valid_0_111 : _GEN_12057; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13087 = 3'h3 == state ? valid_0_112 : _GEN_12058; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13088 = 3'h3 == state ? valid_0_113 : _GEN_12059; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13089 = 3'h3 == state ? valid_0_114 : _GEN_12060; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13090 = 3'h3 == state ? valid_0_115 : _GEN_12061; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13091 = 3'h3 == state ? valid_0_116 : _GEN_12062; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13092 = 3'h3 == state ? valid_0_117 : _GEN_12063; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13093 = 3'h3 == state ? valid_0_118 : _GEN_12064; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13094 = 3'h3 == state ? valid_0_119 : _GEN_12065; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13095 = 3'h3 == state ? valid_0_120 : _GEN_12066; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13096 = 3'h3 == state ? valid_0_121 : _GEN_12067; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13097 = 3'h3 == state ? valid_0_122 : _GEN_12068; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13098 = 3'h3 == state ? valid_0_123 : _GEN_12069; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13099 = 3'h3 == state ? valid_0_124 : _GEN_12070; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13100 = 3'h3 == state ? valid_0_125 : _GEN_12071; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13101 = 3'h3 == state ? valid_0_126 : _GEN_12072; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13102 = 3'h3 == state ? valid_0_127 : _GEN_12073; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_13103 = 3'h3 == state ? quene : _GEN_12074; // @[d_cache.scala 81:18 37:24]
  wire [63:0] _GEN_13104 = 3'h3 == state ? ram_1_0 : _GEN_12075; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13105 = 3'h3 == state ? ram_1_1 : _GEN_12076; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13106 = 3'h3 == state ? ram_1_2 : _GEN_12077; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13107 = 3'h3 == state ? ram_1_3 : _GEN_12078; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13108 = 3'h3 == state ? ram_1_4 : _GEN_12079; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13109 = 3'h3 == state ? ram_1_5 : _GEN_12080; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13110 = 3'h3 == state ? ram_1_6 : _GEN_12081; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13111 = 3'h3 == state ? ram_1_7 : _GEN_12082; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13112 = 3'h3 == state ? ram_1_8 : _GEN_12083; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13113 = 3'h3 == state ? ram_1_9 : _GEN_12084; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13114 = 3'h3 == state ? ram_1_10 : _GEN_12085; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13115 = 3'h3 == state ? ram_1_11 : _GEN_12086; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13116 = 3'h3 == state ? ram_1_12 : _GEN_12087; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13117 = 3'h3 == state ? ram_1_13 : _GEN_12088; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13118 = 3'h3 == state ? ram_1_14 : _GEN_12089; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13119 = 3'h3 == state ? ram_1_15 : _GEN_12090; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13120 = 3'h3 == state ? ram_1_16 : _GEN_12091; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13121 = 3'h3 == state ? ram_1_17 : _GEN_12092; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13122 = 3'h3 == state ? ram_1_18 : _GEN_12093; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13123 = 3'h3 == state ? ram_1_19 : _GEN_12094; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13124 = 3'h3 == state ? ram_1_20 : _GEN_12095; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13125 = 3'h3 == state ? ram_1_21 : _GEN_12096; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13126 = 3'h3 == state ? ram_1_22 : _GEN_12097; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13127 = 3'h3 == state ? ram_1_23 : _GEN_12098; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13128 = 3'h3 == state ? ram_1_24 : _GEN_12099; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13129 = 3'h3 == state ? ram_1_25 : _GEN_12100; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13130 = 3'h3 == state ? ram_1_26 : _GEN_12101; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13131 = 3'h3 == state ? ram_1_27 : _GEN_12102; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13132 = 3'h3 == state ? ram_1_28 : _GEN_12103; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13133 = 3'h3 == state ? ram_1_29 : _GEN_12104; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13134 = 3'h3 == state ? ram_1_30 : _GEN_12105; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13135 = 3'h3 == state ? ram_1_31 : _GEN_12106; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13136 = 3'h3 == state ? ram_1_32 : _GEN_12107; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13137 = 3'h3 == state ? ram_1_33 : _GEN_12108; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13138 = 3'h3 == state ? ram_1_34 : _GEN_12109; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13139 = 3'h3 == state ? ram_1_35 : _GEN_12110; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13140 = 3'h3 == state ? ram_1_36 : _GEN_12111; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13141 = 3'h3 == state ? ram_1_37 : _GEN_12112; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13142 = 3'h3 == state ? ram_1_38 : _GEN_12113; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13143 = 3'h3 == state ? ram_1_39 : _GEN_12114; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13144 = 3'h3 == state ? ram_1_40 : _GEN_12115; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13145 = 3'h3 == state ? ram_1_41 : _GEN_12116; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13146 = 3'h3 == state ? ram_1_42 : _GEN_12117; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13147 = 3'h3 == state ? ram_1_43 : _GEN_12118; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13148 = 3'h3 == state ? ram_1_44 : _GEN_12119; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13149 = 3'h3 == state ? ram_1_45 : _GEN_12120; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13150 = 3'h3 == state ? ram_1_46 : _GEN_12121; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13151 = 3'h3 == state ? ram_1_47 : _GEN_12122; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13152 = 3'h3 == state ? ram_1_48 : _GEN_12123; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13153 = 3'h3 == state ? ram_1_49 : _GEN_12124; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13154 = 3'h3 == state ? ram_1_50 : _GEN_12125; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13155 = 3'h3 == state ? ram_1_51 : _GEN_12126; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13156 = 3'h3 == state ? ram_1_52 : _GEN_12127; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13157 = 3'h3 == state ? ram_1_53 : _GEN_12128; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13158 = 3'h3 == state ? ram_1_54 : _GEN_12129; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13159 = 3'h3 == state ? ram_1_55 : _GEN_12130; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13160 = 3'h3 == state ? ram_1_56 : _GEN_12131; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13161 = 3'h3 == state ? ram_1_57 : _GEN_12132; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13162 = 3'h3 == state ? ram_1_58 : _GEN_12133; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13163 = 3'h3 == state ? ram_1_59 : _GEN_12134; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13164 = 3'h3 == state ? ram_1_60 : _GEN_12135; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13165 = 3'h3 == state ? ram_1_61 : _GEN_12136; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13166 = 3'h3 == state ? ram_1_62 : _GEN_12137; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13167 = 3'h3 == state ? ram_1_63 : _GEN_12138; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13168 = 3'h3 == state ? ram_1_64 : _GEN_12139; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13169 = 3'h3 == state ? ram_1_65 : _GEN_12140; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13170 = 3'h3 == state ? ram_1_66 : _GEN_12141; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13171 = 3'h3 == state ? ram_1_67 : _GEN_12142; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13172 = 3'h3 == state ? ram_1_68 : _GEN_12143; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13173 = 3'h3 == state ? ram_1_69 : _GEN_12144; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13174 = 3'h3 == state ? ram_1_70 : _GEN_12145; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13175 = 3'h3 == state ? ram_1_71 : _GEN_12146; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13176 = 3'h3 == state ? ram_1_72 : _GEN_12147; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13177 = 3'h3 == state ? ram_1_73 : _GEN_12148; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13178 = 3'h3 == state ? ram_1_74 : _GEN_12149; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13179 = 3'h3 == state ? ram_1_75 : _GEN_12150; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13180 = 3'h3 == state ? ram_1_76 : _GEN_12151; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13181 = 3'h3 == state ? ram_1_77 : _GEN_12152; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13182 = 3'h3 == state ? ram_1_78 : _GEN_12153; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13183 = 3'h3 == state ? ram_1_79 : _GEN_12154; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13184 = 3'h3 == state ? ram_1_80 : _GEN_12155; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13185 = 3'h3 == state ? ram_1_81 : _GEN_12156; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13186 = 3'h3 == state ? ram_1_82 : _GEN_12157; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13187 = 3'h3 == state ? ram_1_83 : _GEN_12158; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13188 = 3'h3 == state ? ram_1_84 : _GEN_12159; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13189 = 3'h3 == state ? ram_1_85 : _GEN_12160; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13190 = 3'h3 == state ? ram_1_86 : _GEN_12161; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13191 = 3'h3 == state ? ram_1_87 : _GEN_12162; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13192 = 3'h3 == state ? ram_1_88 : _GEN_12163; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13193 = 3'h3 == state ? ram_1_89 : _GEN_12164; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13194 = 3'h3 == state ? ram_1_90 : _GEN_12165; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13195 = 3'h3 == state ? ram_1_91 : _GEN_12166; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13196 = 3'h3 == state ? ram_1_92 : _GEN_12167; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13197 = 3'h3 == state ? ram_1_93 : _GEN_12168; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13198 = 3'h3 == state ? ram_1_94 : _GEN_12169; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13199 = 3'h3 == state ? ram_1_95 : _GEN_12170; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13200 = 3'h3 == state ? ram_1_96 : _GEN_12171; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13201 = 3'h3 == state ? ram_1_97 : _GEN_12172; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13202 = 3'h3 == state ? ram_1_98 : _GEN_12173; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13203 = 3'h3 == state ? ram_1_99 : _GEN_12174; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13204 = 3'h3 == state ? ram_1_100 : _GEN_12175; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13205 = 3'h3 == state ? ram_1_101 : _GEN_12176; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13206 = 3'h3 == state ? ram_1_102 : _GEN_12177; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13207 = 3'h3 == state ? ram_1_103 : _GEN_12178; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13208 = 3'h3 == state ? ram_1_104 : _GEN_12179; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13209 = 3'h3 == state ? ram_1_105 : _GEN_12180; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13210 = 3'h3 == state ? ram_1_106 : _GEN_12181; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13211 = 3'h3 == state ? ram_1_107 : _GEN_12182; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13212 = 3'h3 == state ? ram_1_108 : _GEN_12183; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13213 = 3'h3 == state ? ram_1_109 : _GEN_12184; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13214 = 3'h3 == state ? ram_1_110 : _GEN_12185; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13215 = 3'h3 == state ? ram_1_111 : _GEN_12186; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13216 = 3'h3 == state ? ram_1_112 : _GEN_12187; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13217 = 3'h3 == state ? ram_1_113 : _GEN_12188; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13218 = 3'h3 == state ? ram_1_114 : _GEN_12189; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13219 = 3'h3 == state ? ram_1_115 : _GEN_12190; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13220 = 3'h3 == state ? ram_1_116 : _GEN_12191; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13221 = 3'h3 == state ? ram_1_117 : _GEN_12192; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13222 = 3'h3 == state ? ram_1_118 : _GEN_12193; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13223 = 3'h3 == state ? ram_1_119 : _GEN_12194; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13224 = 3'h3 == state ? ram_1_120 : _GEN_12195; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13225 = 3'h3 == state ? ram_1_121 : _GEN_12196; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13226 = 3'h3 == state ? ram_1_122 : _GEN_12197; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13227 = 3'h3 == state ? ram_1_123 : _GEN_12198; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13228 = 3'h3 == state ? ram_1_124 : _GEN_12199; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13229 = 3'h3 == state ? ram_1_125 : _GEN_12200; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13230 = 3'h3 == state ? ram_1_126 : _GEN_12201; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_13231 = 3'h3 == state ? ram_1_127 : _GEN_12202; // @[d_cache.scala 81:18 19:24]
  wire [31:0] _GEN_13232 = 3'h3 == state ? tag_1_0 : _GEN_12203; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13233 = 3'h3 == state ? tag_1_1 : _GEN_12204; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13234 = 3'h3 == state ? tag_1_2 : _GEN_12205; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13235 = 3'h3 == state ? tag_1_3 : _GEN_12206; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13236 = 3'h3 == state ? tag_1_4 : _GEN_12207; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13237 = 3'h3 == state ? tag_1_5 : _GEN_12208; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13238 = 3'h3 == state ? tag_1_6 : _GEN_12209; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13239 = 3'h3 == state ? tag_1_7 : _GEN_12210; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13240 = 3'h3 == state ? tag_1_8 : _GEN_12211; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13241 = 3'h3 == state ? tag_1_9 : _GEN_12212; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13242 = 3'h3 == state ? tag_1_10 : _GEN_12213; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13243 = 3'h3 == state ? tag_1_11 : _GEN_12214; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13244 = 3'h3 == state ? tag_1_12 : _GEN_12215; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13245 = 3'h3 == state ? tag_1_13 : _GEN_12216; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13246 = 3'h3 == state ? tag_1_14 : _GEN_12217; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13247 = 3'h3 == state ? tag_1_15 : _GEN_12218; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13248 = 3'h3 == state ? tag_1_16 : _GEN_12219; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13249 = 3'h3 == state ? tag_1_17 : _GEN_12220; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13250 = 3'h3 == state ? tag_1_18 : _GEN_12221; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13251 = 3'h3 == state ? tag_1_19 : _GEN_12222; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13252 = 3'h3 == state ? tag_1_20 : _GEN_12223; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13253 = 3'h3 == state ? tag_1_21 : _GEN_12224; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13254 = 3'h3 == state ? tag_1_22 : _GEN_12225; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13255 = 3'h3 == state ? tag_1_23 : _GEN_12226; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13256 = 3'h3 == state ? tag_1_24 : _GEN_12227; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13257 = 3'h3 == state ? tag_1_25 : _GEN_12228; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13258 = 3'h3 == state ? tag_1_26 : _GEN_12229; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13259 = 3'h3 == state ? tag_1_27 : _GEN_12230; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13260 = 3'h3 == state ? tag_1_28 : _GEN_12231; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13261 = 3'h3 == state ? tag_1_29 : _GEN_12232; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13262 = 3'h3 == state ? tag_1_30 : _GEN_12233; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13263 = 3'h3 == state ? tag_1_31 : _GEN_12234; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13264 = 3'h3 == state ? tag_1_32 : _GEN_12235; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13265 = 3'h3 == state ? tag_1_33 : _GEN_12236; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13266 = 3'h3 == state ? tag_1_34 : _GEN_12237; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13267 = 3'h3 == state ? tag_1_35 : _GEN_12238; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13268 = 3'h3 == state ? tag_1_36 : _GEN_12239; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13269 = 3'h3 == state ? tag_1_37 : _GEN_12240; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13270 = 3'h3 == state ? tag_1_38 : _GEN_12241; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13271 = 3'h3 == state ? tag_1_39 : _GEN_12242; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13272 = 3'h3 == state ? tag_1_40 : _GEN_12243; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13273 = 3'h3 == state ? tag_1_41 : _GEN_12244; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13274 = 3'h3 == state ? tag_1_42 : _GEN_12245; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13275 = 3'h3 == state ? tag_1_43 : _GEN_12246; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13276 = 3'h3 == state ? tag_1_44 : _GEN_12247; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13277 = 3'h3 == state ? tag_1_45 : _GEN_12248; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13278 = 3'h3 == state ? tag_1_46 : _GEN_12249; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13279 = 3'h3 == state ? tag_1_47 : _GEN_12250; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13280 = 3'h3 == state ? tag_1_48 : _GEN_12251; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13281 = 3'h3 == state ? tag_1_49 : _GEN_12252; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13282 = 3'h3 == state ? tag_1_50 : _GEN_12253; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13283 = 3'h3 == state ? tag_1_51 : _GEN_12254; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13284 = 3'h3 == state ? tag_1_52 : _GEN_12255; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13285 = 3'h3 == state ? tag_1_53 : _GEN_12256; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13286 = 3'h3 == state ? tag_1_54 : _GEN_12257; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13287 = 3'h3 == state ? tag_1_55 : _GEN_12258; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13288 = 3'h3 == state ? tag_1_56 : _GEN_12259; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13289 = 3'h3 == state ? tag_1_57 : _GEN_12260; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13290 = 3'h3 == state ? tag_1_58 : _GEN_12261; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13291 = 3'h3 == state ? tag_1_59 : _GEN_12262; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13292 = 3'h3 == state ? tag_1_60 : _GEN_12263; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13293 = 3'h3 == state ? tag_1_61 : _GEN_12264; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13294 = 3'h3 == state ? tag_1_62 : _GEN_12265; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13295 = 3'h3 == state ? tag_1_63 : _GEN_12266; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13296 = 3'h3 == state ? tag_1_64 : _GEN_12267; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13297 = 3'h3 == state ? tag_1_65 : _GEN_12268; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13298 = 3'h3 == state ? tag_1_66 : _GEN_12269; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13299 = 3'h3 == state ? tag_1_67 : _GEN_12270; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13300 = 3'h3 == state ? tag_1_68 : _GEN_12271; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13301 = 3'h3 == state ? tag_1_69 : _GEN_12272; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13302 = 3'h3 == state ? tag_1_70 : _GEN_12273; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13303 = 3'h3 == state ? tag_1_71 : _GEN_12274; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13304 = 3'h3 == state ? tag_1_72 : _GEN_12275; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13305 = 3'h3 == state ? tag_1_73 : _GEN_12276; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13306 = 3'h3 == state ? tag_1_74 : _GEN_12277; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13307 = 3'h3 == state ? tag_1_75 : _GEN_12278; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13308 = 3'h3 == state ? tag_1_76 : _GEN_12279; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13309 = 3'h3 == state ? tag_1_77 : _GEN_12280; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13310 = 3'h3 == state ? tag_1_78 : _GEN_12281; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13311 = 3'h3 == state ? tag_1_79 : _GEN_12282; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13312 = 3'h3 == state ? tag_1_80 : _GEN_12283; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13313 = 3'h3 == state ? tag_1_81 : _GEN_12284; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13314 = 3'h3 == state ? tag_1_82 : _GEN_12285; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13315 = 3'h3 == state ? tag_1_83 : _GEN_12286; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13316 = 3'h3 == state ? tag_1_84 : _GEN_12287; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13317 = 3'h3 == state ? tag_1_85 : _GEN_12288; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13318 = 3'h3 == state ? tag_1_86 : _GEN_12289; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13319 = 3'h3 == state ? tag_1_87 : _GEN_12290; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13320 = 3'h3 == state ? tag_1_88 : _GEN_12291; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13321 = 3'h3 == state ? tag_1_89 : _GEN_12292; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13322 = 3'h3 == state ? tag_1_90 : _GEN_12293; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13323 = 3'h3 == state ? tag_1_91 : _GEN_12294; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13324 = 3'h3 == state ? tag_1_92 : _GEN_12295; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13325 = 3'h3 == state ? tag_1_93 : _GEN_12296; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13326 = 3'h3 == state ? tag_1_94 : _GEN_12297; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13327 = 3'h3 == state ? tag_1_95 : _GEN_12298; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13328 = 3'h3 == state ? tag_1_96 : _GEN_12299; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13329 = 3'h3 == state ? tag_1_97 : _GEN_12300; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13330 = 3'h3 == state ? tag_1_98 : _GEN_12301; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13331 = 3'h3 == state ? tag_1_99 : _GEN_12302; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13332 = 3'h3 == state ? tag_1_100 : _GEN_12303; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13333 = 3'h3 == state ? tag_1_101 : _GEN_12304; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13334 = 3'h3 == state ? tag_1_102 : _GEN_12305; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13335 = 3'h3 == state ? tag_1_103 : _GEN_12306; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13336 = 3'h3 == state ? tag_1_104 : _GEN_12307; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13337 = 3'h3 == state ? tag_1_105 : _GEN_12308; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13338 = 3'h3 == state ? tag_1_106 : _GEN_12309; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13339 = 3'h3 == state ? tag_1_107 : _GEN_12310; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13340 = 3'h3 == state ? tag_1_108 : _GEN_12311; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13341 = 3'h3 == state ? tag_1_109 : _GEN_12312; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13342 = 3'h3 == state ? tag_1_110 : _GEN_12313; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13343 = 3'h3 == state ? tag_1_111 : _GEN_12314; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13344 = 3'h3 == state ? tag_1_112 : _GEN_12315; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13345 = 3'h3 == state ? tag_1_113 : _GEN_12316; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13346 = 3'h3 == state ? tag_1_114 : _GEN_12317; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13347 = 3'h3 == state ? tag_1_115 : _GEN_12318; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13348 = 3'h3 == state ? tag_1_116 : _GEN_12319; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13349 = 3'h3 == state ? tag_1_117 : _GEN_12320; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13350 = 3'h3 == state ? tag_1_118 : _GEN_12321; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13351 = 3'h3 == state ? tag_1_119 : _GEN_12322; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13352 = 3'h3 == state ? tag_1_120 : _GEN_12323; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13353 = 3'h3 == state ? tag_1_121 : _GEN_12324; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13354 = 3'h3 == state ? tag_1_122 : _GEN_12325; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13355 = 3'h3 == state ? tag_1_123 : _GEN_12326; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13356 = 3'h3 == state ? tag_1_124 : _GEN_12327; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13357 = 3'h3 == state ? tag_1_125 : _GEN_12328; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13358 = 3'h3 == state ? tag_1_126 : _GEN_12329; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_13359 = 3'h3 == state ? tag_1_127 : _GEN_12330; // @[d_cache.scala 81:18 23:24]
  wire  _GEN_13360 = 3'h3 == state ? valid_1_0 : _GEN_12331; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13361 = 3'h3 == state ? valid_1_1 : _GEN_12332; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13362 = 3'h3 == state ? valid_1_2 : _GEN_12333; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13363 = 3'h3 == state ? valid_1_3 : _GEN_12334; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13364 = 3'h3 == state ? valid_1_4 : _GEN_12335; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13365 = 3'h3 == state ? valid_1_5 : _GEN_12336; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13366 = 3'h3 == state ? valid_1_6 : _GEN_12337; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13367 = 3'h3 == state ? valid_1_7 : _GEN_12338; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13368 = 3'h3 == state ? valid_1_8 : _GEN_12339; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13369 = 3'h3 == state ? valid_1_9 : _GEN_12340; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13370 = 3'h3 == state ? valid_1_10 : _GEN_12341; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13371 = 3'h3 == state ? valid_1_11 : _GEN_12342; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13372 = 3'h3 == state ? valid_1_12 : _GEN_12343; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13373 = 3'h3 == state ? valid_1_13 : _GEN_12344; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13374 = 3'h3 == state ? valid_1_14 : _GEN_12345; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13375 = 3'h3 == state ? valid_1_15 : _GEN_12346; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13376 = 3'h3 == state ? valid_1_16 : _GEN_12347; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13377 = 3'h3 == state ? valid_1_17 : _GEN_12348; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13378 = 3'h3 == state ? valid_1_18 : _GEN_12349; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13379 = 3'h3 == state ? valid_1_19 : _GEN_12350; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13380 = 3'h3 == state ? valid_1_20 : _GEN_12351; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13381 = 3'h3 == state ? valid_1_21 : _GEN_12352; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13382 = 3'h3 == state ? valid_1_22 : _GEN_12353; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13383 = 3'h3 == state ? valid_1_23 : _GEN_12354; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13384 = 3'h3 == state ? valid_1_24 : _GEN_12355; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13385 = 3'h3 == state ? valid_1_25 : _GEN_12356; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13386 = 3'h3 == state ? valid_1_26 : _GEN_12357; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13387 = 3'h3 == state ? valid_1_27 : _GEN_12358; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13388 = 3'h3 == state ? valid_1_28 : _GEN_12359; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13389 = 3'h3 == state ? valid_1_29 : _GEN_12360; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13390 = 3'h3 == state ? valid_1_30 : _GEN_12361; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13391 = 3'h3 == state ? valid_1_31 : _GEN_12362; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13392 = 3'h3 == state ? valid_1_32 : _GEN_12363; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13393 = 3'h3 == state ? valid_1_33 : _GEN_12364; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13394 = 3'h3 == state ? valid_1_34 : _GEN_12365; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13395 = 3'h3 == state ? valid_1_35 : _GEN_12366; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13396 = 3'h3 == state ? valid_1_36 : _GEN_12367; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13397 = 3'h3 == state ? valid_1_37 : _GEN_12368; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13398 = 3'h3 == state ? valid_1_38 : _GEN_12369; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13399 = 3'h3 == state ? valid_1_39 : _GEN_12370; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13400 = 3'h3 == state ? valid_1_40 : _GEN_12371; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13401 = 3'h3 == state ? valid_1_41 : _GEN_12372; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13402 = 3'h3 == state ? valid_1_42 : _GEN_12373; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13403 = 3'h3 == state ? valid_1_43 : _GEN_12374; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13404 = 3'h3 == state ? valid_1_44 : _GEN_12375; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13405 = 3'h3 == state ? valid_1_45 : _GEN_12376; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13406 = 3'h3 == state ? valid_1_46 : _GEN_12377; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13407 = 3'h3 == state ? valid_1_47 : _GEN_12378; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13408 = 3'h3 == state ? valid_1_48 : _GEN_12379; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13409 = 3'h3 == state ? valid_1_49 : _GEN_12380; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13410 = 3'h3 == state ? valid_1_50 : _GEN_12381; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13411 = 3'h3 == state ? valid_1_51 : _GEN_12382; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13412 = 3'h3 == state ? valid_1_52 : _GEN_12383; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13413 = 3'h3 == state ? valid_1_53 : _GEN_12384; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13414 = 3'h3 == state ? valid_1_54 : _GEN_12385; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13415 = 3'h3 == state ? valid_1_55 : _GEN_12386; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13416 = 3'h3 == state ? valid_1_56 : _GEN_12387; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13417 = 3'h3 == state ? valid_1_57 : _GEN_12388; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13418 = 3'h3 == state ? valid_1_58 : _GEN_12389; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13419 = 3'h3 == state ? valid_1_59 : _GEN_12390; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13420 = 3'h3 == state ? valid_1_60 : _GEN_12391; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13421 = 3'h3 == state ? valid_1_61 : _GEN_12392; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13422 = 3'h3 == state ? valid_1_62 : _GEN_12393; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13423 = 3'h3 == state ? valid_1_63 : _GEN_12394; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13424 = 3'h3 == state ? valid_1_64 : _GEN_12395; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13425 = 3'h3 == state ? valid_1_65 : _GEN_12396; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13426 = 3'h3 == state ? valid_1_66 : _GEN_12397; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13427 = 3'h3 == state ? valid_1_67 : _GEN_12398; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13428 = 3'h3 == state ? valid_1_68 : _GEN_12399; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13429 = 3'h3 == state ? valid_1_69 : _GEN_12400; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13430 = 3'h3 == state ? valid_1_70 : _GEN_12401; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13431 = 3'h3 == state ? valid_1_71 : _GEN_12402; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13432 = 3'h3 == state ? valid_1_72 : _GEN_12403; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13433 = 3'h3 == state ? valid_1_73 : _GEN_12404; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13434 = 3'h3 == state ? valid_1_74 : _GEN_12405; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13435 = 3'h3 == state ? valid_1_75 : _GEN_12406; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13436 = 3'h3 == state ? valid_1_76 : _GEN_12407; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13437 = 3'h3 == state ? valid_1_77 : _GEN_12408; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13438 = 3'h3 == state ? valid_1_78 : _GEN_12409; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13439 = 3'h3 == state ? valid_1_79 : _GEN_12410; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13440 = 3'h3 == state ? valid_1_80 : _GEN_12411; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13441 = 3'h3 == state ? valid_1_81 : _GEN_12412; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13442 = 3'h3 == state ? valid_1_82 : _GEN_12413; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13443 = 3'h3 == state ? valid_1_83 : _GEN_12414; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13444 = 3'h3 == state ? valid_1_84 : _GEN_12415; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13445 = 3'h3 == state ? valid_1_85 : _GEN_12416; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13446 = 3'h3 == state ? valid_1_86 : _GEN_12417; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13447 = 3'h3 == state ? valid_1_87 : _GEN_12418; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13448 = 3'h3 == state ? valid_1_88 : _GEN_12419; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13449 = 3'h3 == state ? valid_1_89 : _GEN_12420; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13450 = 3'h3 == state ? valid_1_90 : _GEN_12421; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13451 = 3'h3 == state ? valid_1_91 : _GEN_12422; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13452 = 3'h3 == state ? valid_1_92 : _GEN_12423; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13453 = 3'h3 == state ? valid_1_93 : _GEN_12424; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13454 = 3'h3 == state ? valid_1_94 : _GEN_12425; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13455 = 3'h3 == state ? valid_1_95 : _GEN_12426; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13456 = 3'h3 == state ? valid_1_96 : _GEN_12427; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13457 = 3'h3 == state ? valid_1_97 : _GEN_12428; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13458 = 3'h3 == state ? valid_1_98 : _GEN_12429; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13459 = 3'h3 == state ? valid_1_99 : _GEN_12430; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13460 = 3'h3 == state ? valid_1_100 : _GEN_12431; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13461 = 3'h3 == state ? valid_1_101 : _GEN_12432; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13462 = 3'h3 == state ? valid_1_102 : _GEN_12433; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13463 = 3'h3 == state ? valid_1_103 : _GEN_12434; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13464 = 3'h3 == state ? valid_1_104 : _GEN_12435; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13465 = 3'h3 == state ? valid_1_105 : _GEN_12436; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13466 = 3'h3 == state ? valid_1_106 : _GEN_12437; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13467 = 3'h3 == state ? valid_1_107 : _GEN_12438; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13468 = 3'h3 == state ? valid_1_108 : _GEN_12439; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13469 = 3'h3 == state ? valid_1_109 : _GEN_12440; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13470 = 3'h3 == state ? valid_1_110 : _GEN_12441; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13471 = 3'h3 == state ? valid_1_111 : _GEN_12442; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13472 = 3'h3 == state ? valid_1_112 : _GEN_12443; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13473 = 3'h3 == state ? valid_1_113 : _GEN_12444; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13474 = 3'h3 == state ? valid_1_114 : _GEN_12445; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13475 = 3'h3 == state ? valid_1_115 : _GEN_12446; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13476 = 3'h3 == state ? valid_1_116 : _GEN_12447; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13477 = 3'h3 == state ? valid_1_117 : _GEN_12448; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13478 = 3'h3 == state ? valid_1_118 : _GEN_12449; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13479 = 3'h3 == state ? valid_1_119 : _GEN_12450; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13480 = 3'h3 == state ? valid_1_120 : _GEN_12451; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13481 = 3'h3 == state ? valid_1_121 : _GEN_12452; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13482 = 3'h3 == state ? valid_1_122 : _GEN_12453; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13483 = 3'h3 == state ? valid_1_123 : _GEN_12454; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13484 = 3'h3 == state ? valid_1_124 : _GEN_12455; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13485 = 3'h3 == state ? valid_1_125 : _GEN_12456; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13486 = 3'h3 == state ? valid_1_126 : _GEN_12457; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_13487 = 3'h3 == state ? valid_1_127 : _GEN_12458; // @[d_cache.scala 81:18 25:26]
  wire [63:0] _GEN_13488 = 3'h3 == state ? write_back_data : _GEN_12459; // @[d_cache.scala 81:18 31:34]
  wire [41:0] _GEN_13489 = 3'h3 == state ? {{10'd0}, write_back_addr} : _GEN_12460; // @[d_cache.scala 81:18 32:34]
  wire  _GEN_13490 = 3'h3 == state ? dirty_0_0 : _GEN_12461; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13491 = 3'h3 == state ? dirty_0_1 : _GEN_12462; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13492 = 3'h3 == state ? dirty_0_2 : _GEN_12463; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13493 = 3'h3 == state ? dirty_0_3 : _GEN_12464; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13494 = 3'h3 == state ? dirty_0_4 : _GEN_12465; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13495 = 3'h3 == state ? dirty_0_5 : _GEN_12466; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13496 = 3'h3 == state ? dirty_0_6 : _GEN_12467; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13497 = 3'h3 == state ? dirty_0_7 : _GEN_12468; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13498 = 3'h3 == state ? dirty_0_8 : _GEN_12469; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13499 = 3'h3 == state ? dirty_0_9 : _GEN_12470; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13500 = 3'h3 == state ? dirty_0_10 : _GEN_12471; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13501 = 3'h3 == state ? dirty_0_11 : _GEN_12472; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13502 = 3'h3 == state ? dirty_0_12 : _GEN_12473; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13503 = 3'h3 == state ? dirty_0_13 : _GEN_12474; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13504 = 3'h3 == state ? dirty_0_14 : _GEN_12475; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13505 = 3'h3 == state ? dirty_0_15 : _GEN_12476; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13506 = 3'h3 == state ? dirty_0_16 : _GEN_12477; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13507 = 3'h3 == state ? dirty_0_17 : _GEN_12478; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13508 = 3'h3 == state ? dirty_0_18 : _GEN_12479; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13509 = 3'h3 == state ? dirty_0_19 : _GEN_12480; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13510 = 3'h3 == state ? dirty_0_20 : _GEN_12481; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13511 = 3'h3 == state ? dirty_0_21 : _GEN_12482; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13512 = 3'h3 == state ? dirty_0_22 : _GEN_12483; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13513 = 3'h3 == state ? dirty_0_23 : _GEN_12484; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13514 = 3'h3 == state ? dirty_0_24 : _GEN_12485; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13515 = 3'h3 == state ? dirty_0_25 : _GEN_12486; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13516 = 3'h3 == state ? dirty_0_26 : _GEN_12487; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13517 = 3'h3 == state ? dirty_0_27 : _GEN_12488; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13518 = 3'h3 == state ? dirty_0_28 : _GEN_12489; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13519 = 3'h3 == state ? dirty_0_29 : _GEN_12490; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13520 = 3'h3 == state ? dirty_0_30 : _GEN_12491; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13521 = 3'h3 == state ? dirty_0_31 : _GEN_12492; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13522 = 3'h3 == state ? dirty_0_32 : _GEN_12493; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13523 = 3'h3 == state ? dirty_0_33 : _GEN_12494; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13524 = 3'h3 == state ? dirty_0_34 : _GEN_12495; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13525 = 3'h3 == state ? dirty_0_35 : _GEN_12496; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13526 = 3'h3 == state ? dirty_0_36 : _GEN_12497; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13527 = 3'h3 == state ? dirty_0_37 : _GEN_12498; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13528 = 3'h3 == state ? dirty_0_38 : _GEN_12499; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13529 = 3'h3 == state ? dirty_0_39 : _GEN_12500; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13530 = 3'h3 == state ? dirty_0_40 : _GEN_12501; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13531 = 3'h3 == state ? dirty_0_41 : _GEN_12502; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13532 = 3'h3 == state ? dirty_0_42 : _GEN_12503; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13533 = 3'h3 == state ? dirty_0_43 : _GEN_12504; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13534 = 3'h3 == state ? dirty_0_44 : _GEN_12505; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13535 = 3'h3 == state ? dirty_0_45 : _GEN_12506; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13536 = 3'h3 == state ? dirty_0_46 : _GEN_12507; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13537 = 3'h3 == state ? dirty_0_47 : _GEN_12508; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13538 = 3'h3 == state ? dirty_0_48 : _GEN_12509; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13539 = 3'h3 == state ? dirty_0_49 : _GEN_12510; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13540 = 3'h3 == state ? dirty_0_50 : _GEN_12511; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13541 = 3'h3 == state ? dirty_0_51 : _GEN_12512; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13542 = 3'h3 == state ? dirty_0_52 : _GEN_12513; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13543 = 3'h3 == state ? dirty_0_53 : _GEN_12514; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13544 = 3'h3 == state ? dirty_0_54 : _GEN_12515; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13545 = 3'h3 == state ? dirty_0_55 : _GEN_12516; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13546 = 3'h3 == state ? dirty_0_56 : _GEN_12517; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13547 = 3'h3 == state ? dirty_0_57 : _GEN_12518; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13548 = 3'h3 == state ? dirty_0_58 : _GEN_12519; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13549 = 3'h3 == state ? dirty_0_59 : _GEN_12520; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13550 = 3'h3 == state ? dirty_0_60 : _GEN_12521; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13551 = 3'h3 == state ? dirty_0_61 : _GEN_12522; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13552 = 3'h3 == state ? dirty_0_62 : _GEN_12523; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13553 = 3'h3 == state ? dirty_0_63 : _GEN_12524; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13554 = 3'h3 == state ? dirty_0_64 : _GEN_12525; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13555 = 3'h3 == state ? dirty_0_65 : _GEN_12526; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13556 = 3'h3 == state ? dirty_0_66 : _GEN_12527; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13557 = 3'h3 == state ? dirty_0_67 : _GEN_12528; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13558 = 3'h3 == state ? dirty_0_68 : _GEN_12529; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13559 = 3'h3 == state ? dirty_0_69 : _GEN_12530; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13560 = 3'h3 == state ? dirty_0_70 : _GEN_12531; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13561 = 3'h3 == state ? dirty_0_71 : _GEN_12532; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13562 = 3'h3 == state ? dirty_0_72 : _GEN_12533; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13563 = 3'h3 == state ? dirty_0_73 : _GEN_12534; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13564 = 3'h3 == state ? dirty_0_74 : _GEN_12535; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13565 = 3'h3 == state ? dirty_0_75 : _GEN_12536; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13566 = 3'h3 == state ? dirty_0_76 : _GEN_12537; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13567 = 3'h3 == state ? dirty_0_77 : _GEN_12538; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13568 = 3'h3 == state ? dirty_0_78 : _GEN_12539; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13569 = 3'h3 == state ? dirty_0_79 : _GEN_12540; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13570 = 3'h3 == state ? dirty_0_80 : _GEN_12541; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13571 = 3'h3 == state ? dirty_0_81 : _GEN_12542; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13572 = 3'h3 == state ? dirty_0_82 : _GEN_12543; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13573 = 3'h3 == state ? dirty_0_83 : _GEN_12544; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13574 = 3'h3 == state ? dirty_0_84 : _GEN_12545; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13575 = 3'h3 == state ? dirty_0_85 : _GEN_12546; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13576 = 3'h3 == state ? dirty_0_86 : _GEN_12547; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13577 = 3'h3 == state ? dirty_0_87 : _GEN_12548; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13578 = 3'h3 == state ? dirty_0_88 : _GEN_12549; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13579 = 3'h3 == state ? dirty_0_89 : _GEN_12550; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13580 = 3'h3 == state ? dirty_0_90 : _GEN_12551; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13581 = 3'h3 == state ? dirty_0_91 : _GEN_12552; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13582 = 3'h3 == state ? dirty_0_92 : _GEN_12553; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13583 = 3'h3 == state ? dirty_0_93 : _GEN_12554; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13584 = 3'h3 == state ? dirty_0_94 : _GEN_12555; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13585 = 3'h3 == state ? dirty_0_95 : _GEN_12556; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13586 = 3'h3 == state ? dirty_0_96 : _GEN_12557; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13587 = 3'h3 == state ? dirty_0_97 : _GEN_12558; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13588 = 3'h3 == state ? dirty_0_98 : _GEN_12559; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13589 = 3'h3 == state ? dirty_0_99 : _GEN_12560; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13590 = 3'h3 == state ? dirty_0_100 : _GEN_12561; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13591 = 3'h3 == state ? dirty_0_101 : _GEN_12562; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13592 = 3'h3 == state ? dirty_0_102 : _GEN_12563; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13593 = 3'h3 == state ? dirty_0_103 : _GEN_12564; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13594 = 3'h3 == state ? dirty_0_104 : _GEN_12565; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13595 = 3'h3 == state ? dirty_0_105 : _GEN_12566; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13596 = 3'h3 == state ? dirty_0_106 : _GEN_12567; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13597 = 3'h3 == state ? dirty_0_107 : _GEN_12568; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13598 = 3'h3 == state ? dirty_0_108 : _GEN_12569; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13599 = 3'h3 == state ? dirty_0_109 : _GEN_12570; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13600 = 3'h3 == state ? dirty_0_110 : _GEN_12571; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13601 = 3'h3 == state ? dirty_0_111 : _GEN_12572; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13602 = 3'h3 == state ? dirty_0_112 : _GEN_12573; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13603 = 3'h3 == state ? dirty_0_113 : _GEN_12574; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13604 = 3'h3 == state ? dirty_0_114 : _GEN_12575; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13605 = 3'h3 == state ? dirty_0_115 : _GEN_12576; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13606 = 3'h3 == state ? dirty_0_116 : _GEN_12577; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13607 = 3'h3 == state ? dirty_0_117 : _GEN_12578; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13608 = 3'h3 == state ? dirty_0_118 : _GEN_12579; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13609 = 3'h3 == state ? dirty_0_119 : _GEN_12580; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13610 = 3'h3 == state ? dirty_0_120 : _GEN_12581; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13611 = 3'h3 == state ? dirty_0_121 : _GEN_12582; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13612 = 3'h3 == state ? dirty_0_122 : _GEN_12583; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13613 = 3'h3 == state ? dirty_0_123 : _GEN_12584; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13614 = 3'h3 == state ? dirty_0_124 : _GEN_12585; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13615 = 3'h3 == state ? dirty_0_125 : _GEN_12586; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13616 = 3'h3 == state ? dirty_0_126 : _GEN_12587; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13617 = 3'h3 == state ? dirty_0_127 : _GEN_12588; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_13618 = 3'h3 == state ? dirty_1_0 : _GEN_12589; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13619 = 3'h3 == state ? dirty_1_1 : _GEN_12590; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13620 = 3'h3 == state ? dirty_1_2 : _GEN_12591; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13621 = 3'h3 == state ? dirty_1_3 : _GEN_12592; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13622 = 3'h3 == state ? dirty_1_4 : _GEN_12593; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13623 = 3'h3 == state ? dirty_1_5 : _GEN_12594; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13624 = 3'h3 == state ? dirty_1_6 : _GEN_12595; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13625 = 3'h3 == state ? dirty_1_7 : _GEN_12596; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13626 = 3'h3 == state ? dirty_1_8 : _GEN_12597; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13627 = 3'h3 == state ? dirty_1_9 : _GEN_12598; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13628 = 3'h3 == state ? dirty_1_10 : _GEN_12599; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13629 = 3'h3 == state ? dirty_1_11 : _GEN_12600; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13630 = 3'h3 == state ? dirty_1_12 : _GEN_12601; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13631 = 3'h3 == state ? dirty_1_13 : _GEN_12602; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13632 = 3'h3 == state ? dirty_1_14 : _GEN_12603; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13633 = 3'h3 == state ? dirty_1_15 : _GEN_12604; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13634 = 3'h3 == state ? dirty_1_16 : _GEN_12605; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13635 = 3'h3 == state ? dirty_1_17 : _GEN_12606; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13636 = 3'h3 == state ? dirty_1_18 : _GEN_12607; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13637 = 3'h3 == state ? dirty_1_19 : _GEN_12608; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13638 = 3'h3 == state ? dirty_1_20 : _GEN_12609; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13639 = 3'h3 == state ? dirty_1_21 : _GEN_12610; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13640 = 3'h3 == state ? dirty_1_22 : _GEN_12611; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13641 = 3'h3 == state ? dirty_1_23 : _GEN_12612; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13642 = 3'h3 == state ? dirty_1_24 : _GEN_12613; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13643 = 3'h3 == state ? dirty_1_25 : _GEN_12614; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13644 = 3'h3 == state ? dirty_1_26 : _GEN_12615; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13645 = 3'h3 == state ? dirty_1_27 : _GEN_12616; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13646 = 3'h3 == state ? dirty_1_28 : _GEN_12617; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13647 = 3'h3 == state ? dirty_1_29 : _GEN_12618; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13648 = 3'h3 == state ? dirty_1_30 : _GEN_12619; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13649 = 3'h3 == state ? dirty_1_31 : _GEN_12620; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13650 = 3'h3 == state ? dirty_1_32 : _GEN_12621; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13651 = 3'h3 == state ? dirty_1_33 : _GEN_12622; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13652 = 3'h3 == state ? dirty_1_34 : _GEN_12623; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13653 = 3'h3 == state ? dirty_1_35 : _GEN_12624; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13654 = 3'h3 == state ? dirty_1_36 : _GEN_12625; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13655 = 3'h3 == state ? dirty_1_37 : _GEN_12626; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13656 = 3'h3 == state ? dirty_1_38 : _GEN_12627; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13657 = 3'h3 == state ? dirty_1_39 : _GEN_12628; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13658 = 3'h3 == state ? dirty_1_40 : _GEN_12629; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13659 = 3'h3 == state ? dirty_1_41 : _GEN_12630; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13660 = 3'h3 == state ? dirty_1_42 : _GEN_12631; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13661 = 3'h3 == state ? dirty_1_43 : _GEN_12632; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13662 = 3'h3 == state ? dirty_1_44 : _GEN_12633; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13663 = 3'h3 == state ? dirty_1_45 : _GEN_12634; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13664 = 3'h3 == state ? dirty_1_46 : _GEN_12635; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13665 = 3'h3 == state ? dirty_1_47 : _GEN_12636; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13666 = 3'h3 == state ? dirty_1_48 : _GEN_12637; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13667 = 3'h3 == state ? dirty_1_49 : _GEN_12638; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13668 = 3'h3 == state ? dirty_1_50 : _GEN_12639; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13669 = 3'h3 == state ? dirty_1_51 : _GEN_12640; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13670 = 3'h3 == state ? dirty_1_52 : _GEN_12641; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13671 = 3'h3 == state ? dirty_1_53 : _GEN_12642; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13672 = 3'h3 == state ? dirty_1_54 : _GEN_12643; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13673 = 3'h3 == state ? dirty_1_55 : _GEN_12644; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13674 = 3'h3 == state ? dirty_1_56 : _GEN_12645; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13675 = 3'h3 == state ? dirty_1_57 : _GEN_12646; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13676 = 3'h3 == state ? dirty_1_58 : _GEN_12647; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13677 = 3'h3 == state ? dirty_1_59 : _GEN_12648; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13678 = 3'h3 == state ? dirty_1_60 : _GEN_12649; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13679 = 3'h3 == state ? dirty_1_61 : _GEN_12650; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13680 = 3'h3 == state ? dirty_1_62 : _GEN_12651; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13681 = 3'h3 == state ? dirty_1_63 : _GEN_12652; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13682 = 3'h3 == state ? dirty_1_64 : _GEN_12653; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13683 = 3'h3 == state ? dirty_1_65 : _GEN_12654; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13684 = 3'h3 == state ? dirty_1_66 : _GEN_12655; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13685 = 3'h3 == state ? dirty_1_67 : _GEN_12656; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13686 = 3'h3 == state ? dirty_1_68 : _GEN_12657; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13687 = 3'h3 == state ? dirty_1_69 : _GEN_12658; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13688 = 3'h3 == state ? dirty_1_70 : _GEN_12659; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13689 = 3'h3 == state ? dirty_1_71 : _GEN_12660; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13690 = 3'h3 == state ? dirty_1_72 : _GEN_12661; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13691 = 3'h3 == state ? dirty_1_73 : _GEN_12662; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13692 = 3'h3 == state ? dirty_1_74 : _GEN_12663; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13693 = 3'h3 == state ? dirty_1_75 : _GEN_12664; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13694 = 3'h3 == state ? dirty_1_76 : _GEN_12665; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13695 = 3'h3 == state ? dirty_1_77 : _GEN_12666; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13696 = 3'h3 == state ? dirty_1_78 : _GEN_12667; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13697 = 3'h3 == state ? dirty_1_79 : _GEN_12668; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13698 = 3'h3 == state ? dirty_1_80 : _GEN_12669; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13699 = 3'h3 == state ? dirty_1_81 : _GEN_12670; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13700 = 3'h3 == state ? dirty_1_82 : _GEN_12671; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13701 = 3'h3 == state ? dirty_1_83 : _GEN_12672; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13702 = 3'h3 == state ? dirty_1_84 : _GEN_12673; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13703 = 3'h3 == state ? dirty_1_85 : _GEN_12674; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13704 = 3'h3 == state ? dirty_1_86 : _GEN_12675; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13705 = 3'h3 == state ? dirty_1_87 : _GEN_12676; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13706 = 3'h3 == state ? dirty_1_88 : _GEN_12677; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13707 = 3'h3 == state ? dirty_1_89 : _GEN_12678; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13708 = 3'h3 == state ? dirty_1_90 : _GEN_12679; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13709 = 3'h3 == state ? dirty_1_91 : _GEN_12680; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13710 = 3'h3 == state ? dirty_1_92 : _GEN_12681; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13711 = 3'h3 == state ? dirty_1_93 : _GEN_12682; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13712 = 3'h3 == state ? dirty_1_94 : _GEN_12683; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13713 = 3'h3 == state ? dirty_1_95 : _GEN_12684; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13714 = 3'h3 == state ? dirty_1_96 : _GEN_12685; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13715 = 3'h3 == state ? dirty_1_97 : _GEN_12686; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13716 = 3'h3 == state ? dirty_1_98 : _GEN_12687; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13717 = 3'h3 == state ? dirty_1_99 : _GEN_12688; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13718 = 3'h3 == state ? dirty_1_100 : _GEN_12689; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13719 = 3'h3 == state ? dirty_1_101 : _GEN_12690; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13720 = 3'h3 == state ? dirty_1_102 : _GEN_12691; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13721 = 3'h3 == state ? dirty_1_103 : _GEN_12692; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13722 = 3'h3 == state ? dirty_1_104 : _GEN_12693; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13723 = 3'h3 == state ? dirty_1_105 : _GEN_12694; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13724 = 3'h3 == state ? dirty_1_106 : _GEN_12695; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13725 = 3'h3 == state ? dirty_1_107 : _GEN_12696; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13726 = 3'h3 == state ? dirty_1_108 : _GEN_12697; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13727 = 3'h3 == state ? dirty_1_109 : _GEN_12698; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13728 = 3'h3 == state ? dirty_1_110 : _GEN_12699; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13729 = 3'h3 == state ? dirty_1_111 : _GEN_12700; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13730 = 3'h3 == state ? dirty_1_112 : _GEN_12701; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13731 = 3'h3 == state ? dirty_1_113 : _GEN_12702; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13732 = 3'h3 == state ? dirty_1_114 : _GEN_12703; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13733 = 3'h3 == state ? dirty_1_115 : _GEN_12704; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13734 = 3'h3 == state ? dirty_1_116 : _GEN_12705; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13735 = 3'h3 == state ? dirty_1_117 : _GEN_12706; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13736 = 3'h3 == state ? dirty_1_118 : _GEN_12707; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13737 = 3'h3 == state ? dirty_1_119 : _GEN_12708; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13738 = 3'h3 == state ? dirty_1_120 : _GEN_12709; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13739 = 3'h3 == state ? dirty_1_121 : _GEN_12710; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13740 = 3'h3 == state ? dirty_1_122 : _GEN_12711; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13741 = 3'h3 == state ? dirty_1_123 : _GEN_12712; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13742 = 3'h3 == state ? dirty_1_124 : _GEN_12713; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13743 = 3'h3 == state ? dirty_1_125 : _GEN_12714; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13744 = 3'h3 == state ? dirty_1_126 : _GEN_12715; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_13745 = 3'h3 == state ? dirty_1_127 : _GEN_12716; // @[d_cache.scala 81:18 27:26]
  wire [41:0] _GEN_15030 = 3'h2 == state ? {{10'd0}, write_back_addr} : _GEN_13489; // @[d_cache.scala 81:18 32:34]
  wire [41:0] _GEN_16315 = 3'h1 == state ? {{10'd0}, write_back_addr} : _GEN_15030; // @[d_cache.scala 81:18 32:34]
  wire [41:0] _GEN_17600 = 3'h0 == state ? {{10'd0}, write_back_addr} : _GEN_16315; // @[d_cache.scala 81:18 32:34]
  wire [63:0] _io_to_lsu_rdata_T_1 = _GEN_1160 >> shift_bit; // @[d_cache.scala 226:49]
  wire [63:0] _io_to_lsu_rdata_T_3 = _GEN_1672 >> shift_bit; // @[d_cache.scala 233:49]
  wire [63:0] _GEN_17857 = way1_hit ? _io_to_lsu_rdata_T_3 : 64'h0; // @[d_cache.scala 232:33 233:33 240:33]
  wire [63:0] _GEN_17861 = way0_hit ? _io_to_lsu_rdata_T_1 : _GEN_17857; // @[d_cache.scala 225:23 226:33]
  wire  _GEN_17863 = way0_hit | way1_hit; // @[d_cache.scala 225:23 228:34]
  wire  _GEN_17865 = way1_hit ? 1'h0 : 1'h1; // @[d_cache.scala 264:33 266:35 273:35]
  wire  _GEN_17866 = way0_hit ? 1'h0 : _GEN_17865; // @[d_cache.scala 257:23 259:35]
  wire  _T_70 = state == 3'h3; // @[d_cache.scala 279:21]
  wire [63:0] _GEN_19499 = {{32'd0}, io_from_lsu_araddr}; // @[d_cache.scala 287:48]
  wire [63:0] _io_to_axi_araddr_T = _GEN_19499 & 64'hfffffffffffffff8; // @[d_cache.scala 287:48]
  wire  _T_73 = state == 3'h6; // @[d_cache.scala 328:21]
  wire [31:0] _GEN_17869 = state == 3'h6 ? 32'h0 : io_from_lsu_araddr; // @[d_cache.scala 328:35 336:26 352:26]
  wire  _GEN_17870 = state == 3'h6 ? 1'h0 : io_from_lsu_rready; // @[d_cache.scala 328:35 337:26 353:26]
  wire [31:0] _GEN_17871 = state == 3'h6 ? write_back_addr : 32'h0; // @[d_cache.scala 328:35 338:26 354:26]
  wire [63:0] _GEN_17872 = state == 3'h6 ? write_back_data : 64'h0; // @[d_cache.scala 328:35 340:25 356:25]
  wire [7:0] _GEN_17873 = state == 3'h6 ? 8'hff : 8'h0; // @[d_cache.scala 328:35 341:25 357:25]
  wire  _GEN_17875 = state == 3'h5 | _T_73; // @[d_cache.scala 312:31 314:27]
  wire [31:0] _GEN_17876 = state == 3'h5 ? io_from_lsu_araddr : _GEN_17869; // @[d_cache.scala 312:31 320:26]
  wire  _GEN_17877 = state == 3'h5 ? io_from_lsu_rready : _GEN_17870; // @[d_cache.scala 312:31 321:26]
  wire [31:0] _GEN_17878 = state == 3'h5 ? 32'h0 : _GEN_17871; // @[d_cache.scala 312:31 322:26]
  wire  _GEN_17879 = state == 3'h5 ? 1'h0 : _T_73; // @[d_cache.scala 312:31 323:27]
  wire [63:0] _GEN_17880 = state == 3'h5 ? 64'h0 : _GEN_17872; // @[d_cache.scala 312:31 324:25]
  wire [7:0] _GEN_17881 = state == 3'h5 ? 8'h0 : _GEN_17873; // @[d_cache.scala 312:31 325:25]
  wire  _GEN_17883 = state == 3'h4 | _GEN_17875; // @[d_cache.scala 295:31 297:27]
  wire  _GEN_17884 = state == 3'h4 & io_from_axi_wready; // @[d_cache.scala 295:31 299:26]
  wire  _GEN_17885 = state == 3'h4 & io_from_axi_bvalid; // @[d_cache.scala 295:31 300:26]
  wire  _GEN_17886 = state == 3'h4 & io_from_axi_awready; // @[d_cache.scala 295:31 301:27]
  wire [31:0] _GEN_17887 = state == 3'h4 ? 32'h0 : _GEN_17876; // @[d_cache.scala 295:31 303:26]
  wire  _GEN_17888 = state == 3'h4 ? io_from_lsu_rready : _GEN_17877; // @[d_cache.scala 295:31 304:26]
  wire [31:0] _GEN_17889 = state == 3'h4 ? io_from_lsu_awaddr : _GEN_17878; // @[d_cache.scala 295:31 305:26]
  wire  _GEN_17890 = state == 3'h4 ? io_from_lsu_awvalid : _GEN_17879; // @[d_cache.scala 295:31 306:27]
  wire [63:0] _GEN_17891 = state == 3'h4 ? {{32'd0}, io_from_lsu_wdata} : _GEN_17880; // @[d_cache.scala 295:31 307:25]
  wire [7:0] _GEN_17892 = state == 3'h4 ? io_from_lsu_wstrb : _GEN_17881; // @[d_cache.scala 295:31 308:25]
  wire  _GEN_17893 = state == 3'h4 ? io_from_lsu_wvalid : _GEN_17879; // @[d_cache.scala 295:31 309:26]
  wire  _GEN_17894 = state == 3'h4 ? io_from_lsu_bready : _GEN_17879; // @[d_cache.scala 295:31 310:26]
  wire  _GEN_17896 = state == 3'h3 | _GEN_17883; // @[d_cache.scala 279:31 281:27]
  wire  _GEN_17897 = state == 3'h3 ? 1'h0 : _GEN_17884; // @[d_cache.scala 279:31 283:26]
  wire  _GEN_17898 = state == 3'h3 ? 1'h0 : _GEN_17885; // @[d_cache.scala 279:31 284:26]
  wire  _GEN_17899 = state == 3'h3 ? 1'h0 : _GEN_17886; // @[d_cache.scala 279:31 285:27]
  wire [63:0] _GEN_17901 = state == 3'h3 ? _io_to_axi_araddr_T : {{32'd0}, _GEN_17887}; // @[d_cache.scala 279:31 287:26]
  wire  _GEN_17902 = state == 3'h3 ? io_from_lsu_rready : _GEN_17888; // @[d_cache.scala 279:31 288:26]
  wire [31:0] _GEN_17903 = state == 3'h3 ? 32'h0 : _GEN_17889; // @[d_cache.scala 279:31 289:26]
  wire  _GEN_17904 = state == 3'h3 ? 1'h0 : _GEN_17890; // @[d_cache.scala 279:31 290:27]
  wire [63:0] _GEN_17905 = state == 3'h3 ? 64'h0 : _GEN_17891; // @[d_cache.scala 279:31 291:25]
  wire [7:0] _GEN_17906 = state == 3'h3 ? 8'h0 : _GEN_17892; // @[d_cache.scala 279:31 292:25]
  wire  _GEN_17907 = state == 3'h3 ? 1'h0 : _GEN_17893; // @[d_cache.scala 279:31 293:26]
  wire  _GEN_17908 = state == 3'h3 ? 1'h0 : _GEN_17894; // @[d_cache.scala 279:31 294:26]
  wire  _GEN_17909 = state == 3'h2 ? 1'h0 : _T_70; // @[d_cache.scala 247:33 248:27]
  wire [63:0] _GEN_17910 = state == 3'h2 ? {{32'd0}, io_from_lsu_araddr} : _GEN_17901; // @[d_cache.scala 247:33 249:26]
  wire  _GEN_17911 = state == 3'h2 ? 1'h0 : _GEN_17902; // @[d_cache.scala 247:33 250:26]
  wire [31:0] _GEN_17912 = state == 3'h2 ? 32'h0 : _GEN_17903; // @[d_cache.scala 247:33 251:26]
  wire  _GEN_17913 = state == 3'h2 ? 1'h0 : _GEN_17904; // @[d_cache.scala 247:33 252:27]
  wire [63:0] _GEN_17914 = state == 3'h2 ? 64'h0 : _GEN_17905; // @[d_cache.scala 247:33 253:25]
  wire [7:0] _GEN_17915 = state == 3'h2 ? 8'h0 : _GEN_17906; // @[d_cache.scala 247:33 254:25]
  wire  _GEN_17916 = state == 3'h2 ? 1'h0 : _GEN_17907; // @[d_cache.scala 247:33 255:26]
  wire  _GEN_17917 = state == 3'h2 ? 1'h0 : _GEN_17908; // @[d_cache.scala 247:33 256:26]
  wire  _GEN_17919 = state == 3'h2 ? _GEN_17866 : _GEN_17896; // @[d_cache.scala 247:33]
  wire  _GEN_17920 = state == 3'h2 ? _GEN_17863 : _GEN_17897; // @[d_cache.scala 247:33]
  wire  _GEN_17921 = state == 3'h2 ? _GEN_17863 : _GEN_17899; // @[d_cache.scala 247:33]
  wire  _GEN_17922 = state == 3'h2 ? _GEN_17863 : _GEN_17898; // @[d_cache.scala 247:33]
  wire  _GEN_17923 = state == 3'h1 ? 1'h0 : _GEN_17909; // @[d_cache.scala 215:33 216:27]
  wire [63:0] _GEN_17924 = state == 3'h1 ? {{32'd0}, io_from_lsu_araddr} : _GEN_17910; // @[d_cache.scala 215:33 217:26]
  wire  _GEN_17925 = state == 3'h1 ? io_from_lsu_rready : _GEN_17911; // @[d_cache.scala 215:33 218:26]
  wire [31:0] _GEN_17926 = state == 3'h1 ? 32'h0 : _GEN_17912; // @[d_cache.scala 215:33 219:26]
  wire  _GEN_17927 = state == 3'h1 ? 1'h0 : _GEN_17913; // @[d_cache.scala 215:33 220:27]
  wire [63:0] _GEN_17928 = state == 3'h1 ? 64'h0 : _GEN_17914; // @[d_cache.scala 215:33 221:25]
  wire [7:0] _GEN_17929 = state == 3'h1 ? 8'h0 : _GEN_17915; // @[d_cache.scala 215:33 222:25]
  wire  _GEN_17930 = state == 3'h1 ? 1'h0 : _GEN_17916; // @[d_cache.scala 215:33 223:26]
  wire  _GEN_17931 = state == 3'h1 ? io_from_lsu_bready : _GEN_17917; // @[d_cache.scala 215:33 224:26]
  wire [63:0] _GEN_17932 = state == 3'h1 ? _GEN_17861 : 64'h0; // @[d_cache.scala 215:33]
  wire  _GEN_17933 = state == 3'h1 | _GEN_17919; // @[d_cache.scala 215:33]
  wire  _GEN_17934 = state == 3'h1 & _GEN_17863; // @[d_cache.scala 215:33]
  wire  _GEN_17935 = state == 3'h1 ? 1'h0 : _GEN_17920; // @[d_cache.scala 215:33]
  wire  _GEN_17936 = state == 3'h1 ? 1'h0 : _GEN_17921; // @[d_cache.scala 215:33]
  wire  _GEN_17937 = state == 3'h1 ? 1'h0 : _GEN_17922; // @[d_cache.scala 215:33]
  wire [63:0] _GEN_17945 = state == 3'h0 ? {{32'd0}, io_from_lsu_araddr} : _GEN_17924; // @[d_cache.scala 199:23 207:26]
  wire [63:0] _GEN_17949 = state == 3'h0 ? 64'h0 : _GEN_17928; // @[d_cache.scala 199:23 211:25]
  wire [63:0] _GEN_18210 = 7'h1 == index[6:0] ? recent_wdata0_1 : recent_wdata0_0; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18211 = 7'h2 == index[6:0] ? recent_wdata0_2 : _GEN_18210; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18212 = 7'h3 == index[6:0] ? recent_wdata0_3 : _GEN_18211; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18213 = 7'h4 == index[6:0] ? recent_wdata0_4 : _GEN_18212; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18214 = 7'h5 == index[6:0] ? recent_wdata0_5 : _GEN_18213; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18215 = 7'h6 == index[6:0] ? recent_wdata0_6 : _GEN_18214; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18216 = 7'h7 == index[6:0] ? recent_wdata0_7 : _GEN_18215; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18217 = 7'h8 == index[6:0] ? recent_wdata0_8 : _GEN_18216; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18218 = 7'h9 == index[6:0] ? recent_wdata0_9 : _GEN_18217; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18219 = 7'ha == index[6:0] ? recent_wdata0_10 : _GEN_18218; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18220 = 7'hb == index[6:0] ? recent_wdata0_11 : _GEN_18219; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18221 = 7'hc == index[6:0] ? recent_wdata0_12 : _GEN_18220; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18222 = 7'hd == index[6:0] ? recent_wdata0_13 : _GEN_18221; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18223 = 7'he == index[6:0] ? recent_wdata0_14 : _GEN_18222; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18224 = 7'hf == index[6:0] ? recent_wdata0_15 : _GEN_18223; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18225 = 7'h10 == index[6:0] ? recent_wdata0_16 : _GEN_18224; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18226 = 7'h11 == index[6:0] ? recent_wdata0_17 : _GEN_18225; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18227 = 7'h12 == index[6:0] ? recent_wdata0_18 : _GEN_18226; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18228 = 7'h13 == index[6:0] ? recent_wdata0_19 : _GEN_18227; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18229 = 7'h14 == index[6:0] ? recent_wdata0_20 : _GEN_18228; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18230 = 7'h15 == index[6:0] ? recent_wdata0_21 : _GEN_18229; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18231 = 7'h16 == index[6:0] ? recent_wdata0_22 : _GEN_18230; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18232 = 7'h17 == index[6:0] ? recent_wdata0_23 : _GEN_18231; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18233 = 7'h18 == index[6:0] ? recent_wdata0_24 : _GEN_18232; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18234 = 7'h19 == index[6:0] ? recent_wdata0_25 : _GEN_18233; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18235 = 7'h1a == index[6:0] ? recent_wdata0_26 : _GEN_18234; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18236 = 7'h1b == index[6:0] ? recent_wdata0_27 : _GEN_18235; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18237 = 7'h1c == index[6:0] ? recent_wdata0_28 : _GEN_18236; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18238 = 7'h1d == index[6:0] ? recent_wdata0_29 : _GEN_18237; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18239 = 7'h1e == index[6:0] ? recent_wdata0_30 : _GEN_18238; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18240 = 7'h1f == index[6:0] ? recent_wdata0_31 : _GEN_18239; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18241 = 7'h20 == index[6:0] ? recent_wdata0_32 : _GEN_18240; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18242 = 7'h21 == index[6:0] ? recent_wdata0_33 : _GEN_18241; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18243 = 7'h22 == index[6:0] ? recent_wdata0_34 : _GEN_18242; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18244 = 7'h23 == index[6:0] ? recent_wdata0_35 : _GEN_18243; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18245 = 7'h24 == index[6:0] ? recent_wdata0_36 : _GEN_18244; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18246 = 7'h25 == index[6:0] ? recent_wdata0_37 : _GEN_18245; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18247 = 7'h26 == index[6:0] ? recent_wdata0_38 : _GEN_18246; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18248 = 7'h27 == index[6:0] ? recent_wdata0_39 : _GEN_18247; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18249 = 7'h28 == index[6:0] ? recent_wdata0_40 : _GEN_18248; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18250 = 7'h29 == index[6:0] ? recent_wdata0_41 : _GEN_18249; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18251 = 7'h2a == index[6:0] ? recent_wdata0_42 : _GEN_18250; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18252 = 7'h2b == index[6:0] ? recent_wdata0_43 : _GEN_18251; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18253 = 7'h2c == index[6:0] ? recent_wdata0_44 : _GEN_18252; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18254 = 7'h2d == index[6:0] ? recent_wdata0_45 : _GEN_18253; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18255 = 7'h2e == index[6:0] ? recent_wdata0_46 : _GEN_18254; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18256 = 7'h2f == index[6:0] ? recent_wdata0_47 : _GEN_18255; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18257 = 7'h30 == index[6:0] ? recent_wdata0_48 : _GEN_18256; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18258 = 7'h31 == index[6:0] ? recent_wdata0_49 : _GEN_18257; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18259 = 7'h32 == index[6:0] ? recent_wdata0_50 : _GEN_18258; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18260 = 7'h33 == index[6:0] ? recent_wdata0_51 : _GEN_18259; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18261 = 7'h34 == index[6:0] ? recent_wdata0_52 : _GEN_18260; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18262 = 7'h35 == index[6:0] ? recent_wdata0_53 : _GEN_18261; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18263 = 7'h36 == index[6:0] ? recent_wdata0_54 : _GEN_18262; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18264 = 7'h37 == index[6:0] ? recent_wdata0_55 : _GEN_18263; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18265 = 7'h38 == index[6:0] ? recent_wdata0_56 : _GEN_18264; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18266 = 7'h39 == index[6:0] ? recent_wdata0_57 : _GEN_18265; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18267 = 7'h3a == index[6:0] ? recent_wdata0_58 : _GEN_18266; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18268 = 7'h3b == index[6:0] ? recent_wdata0_59 : _GEN_18267; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18269 = 7'h3c == index[6:0] ? recent_wdata0_60 : _GEN_18268; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18270 = 7'h3d == index[6:0] ? recent_wdata0_61 : _GEN_18269; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18271 = 7'h3e == index[6:0] ? recent_wdata0_62 : _GEN_18270; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18272 = 7'h3f == index[6:0] ? recent_wdata0_63 : _GEN_18271; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18273 = 7'h40 == index[6:0] ? recent_wdata0_64 : _GEN_18272; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18274 = 7'h41 == index[6:0] ? recent_wdata0_65 : _GEN_18273; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18275 = 7'h42 == index[6:0] ? recent_wdata0_66 : _GEN_18274; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18276 = 7'h43 == index[6:0] ? recent_wdata0_67 : _GEN_18275; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18277 = 7'h44 == index[6:0] ? recent_wdata0_68 : _GEN_18276; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18278 = 7'h45 == index[6:0] ? recent_wdata0_69 : _GEN_18277; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18279 = 7'h46 == index[6:0] ? recent_wdata0_70 : _GEN_18278; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18280 = 7'h47 == index[6:0] ? recent_wdata0_71 : _GEN_18279; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18281 = 7'h48 == index[6:0] ? recent_wdata0_72 : _GEN_18280; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18282 = 7'h49 == index[6:0] ? recent_wdata0_73 : _GEN_18281; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18283 = 7'h4a == index[6:0] ? recent_wdata0_74 : _GEN_18282; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18284 = 7'h4b == index[6:0] ? recent_wdata0_75 : _GEN_18283; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18285 = 7'h4c == index[6:0] ? recent_wdata0_76 : _GEN_18284; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18286 = 7'h4d == index[6:0] ? recent_wdata0_77 : _GEN_18285; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18287 = 7'h4e == index[6:0] ? recent_wdata0_78 : _GEN_18286; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18288 = 7'h4f == index[6:0] ? recent_wdata0_79 : _GEN_18287; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18289 = 7'h50 == index[6:0] ? recent_wdata0_80 : _GEN_18288; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18290 = 7'h51 == index[6:0] ? recent_wdata0_81 : _GEN_18289; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18291 = 7'h52 == index[6:0] ? recent_wdata0_82 : _GEN_18290; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18292 = 7'h53 == index[6:0] ? recent_wdata0_83 : _GEN_18291; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18293 = 7'h54 == index[6:0] ? recent_wdata0_84 : _GEN_18292; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18294 = 7'h55 == index[6:0] ? recent_wdata0_85 : _GEN_18293; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18295 = 7'h56 == index[6:0] ? recent_wdata0_86 : _GEN_18294; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18296 = 7'h57 == index[6:0] ? recent_wdata0_87 : _GEN_18295; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18297 = 7'h58 == index[6:0] ? recent_wdata0_88 : _GEN_18296; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18298 = 7'h59 == index[6:0] ? recent_wdata0_89 : _GEN_18297; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18299 = 7'h5a == index[6:0] ? recent_wdata0_90 : _GEN_18298; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18300 = 7'h5b == index[6:0] ? recent_wdata0_91 : _GEN_18299; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18301 = 7'h5c == index[6:0] ? recent_wdata0_92 : _GEN_18300; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18302 = 7'h5d == index[6:0] ? recent_wdata0_93 : _GEN_18301; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18303 = 7'h5e == index[6:0] ? recent_wdata0_94 : _GEN_18302; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18304 = 7'h5f == index[6:0] ? recent_wdata0_95 : _GEN_18303; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18305 = 7'h60 == index[6:0] ? recent_wdata0_96 : _GEN_18304; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18306 = 7'h61 == index[6:0] ? recent_wdata0_97 : _GEN_18305; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18307 = 7'h62 == index[6:0] ? recent_wdata0_98 : _GEN_18306; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18308 = 7'h63 == index[6:0] ? recent_wdata0_99 : _GEN_18307; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18309 = 7'h64 == index[6:0] ? recent_wdata0_100 : _GEN_18308; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18310 = 7'h65 == index[6:0] ? recent_wdata0_101 : _GEN_18309; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18311 = 7'h66 == index[6:0] ? recent_wdata0_102 : _GEN_18310; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18312 = 7'h67 == index[6:0] ? recent_wdata0_103 : _GEN_18311; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18313 = 7'h68 == index[6:0] ? recent_wdata0_104 : _GEN_18312; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18314 = 7'h69 == index[6:0] ? recent_wdata0_105 : _GEN_18313; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18315 = 7'h6a == index[6:0] ? recent_wdata0_106 : _GEN_18314; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18316 = 7'h6b == index[6:0] ? recent_wdata0_107 : _GEN_18315; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18317 = 7'h6c == index[6:0] ? recent_wdata0_108 : _GEN_18316; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18318 = 7'h6d == index[6:0] ? recent_wdata0_109 : _GEN_18317; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18319 = 7'h6e == index[6:0] ? recent_wdata0_110 : _GEN_18318; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18320 = 7'h6f == index[6:0] ? recent_wdata0_111 : _GEN_18319; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18321 = 7'h70 == index[6:0] ? recent_wdata0_112 : _GEN_18320; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18322 = 7'h71 == index[6:0] ? recent_wdata0_113 : _GEN_18321; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18323 = 7'h72 == index[6:0] ? recent_wdata0_114 : _GEN_18322; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18324 = 7'h73 == index[6:0] ? recent_wdata0_115 : _GEN_18323; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18325 = 7'h74 == index[6:0] ? recent_wdata0_116 : _GEN_18324; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18326 = 7'h75 == index[6:0] ? recent_wdata0_117 : _GEN_18325; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18327 = 7'h76 == index[6:0] ? recent_wdata0_118 : _GEN_18326; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18328 = 7'h77 == index[6:0] ? recent_wdata0_119 : _GEN_18327; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18329 = 7'h78 == index[6:0] ? recent_wdata0_120 : _GEN_18328; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18330 = 7'h79 == index[6:0] ? recent_wdata0_121 : _GEN_18329; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18331 = 7'h7a == index[6:0] ? recent_wdata0_122 : _GEN_18330; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18332 = 7'h7b == index[6:0] ? recent_wdata0_123 : _GEN_18331; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18333 = 7'h7c == index[6:0] ? recent_wdata0_124 : _GEN_18332; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18334 = 7'h7d == index[6:0] ? recent_wdata0_125 : _GEN_18333; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18335 = 7'h7e == index[6:0] ? recent_wdata0_126 : _GEN_18334; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18338 = 7'h1 == index[6:0] ? recent_wdata1_1 : recent_wdata1_0; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18339 = 7'h2 == index[6:0] ? recent_wdata1_2 : _GEN_18338; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18340 = 7'h3 == index[6:0] ? recent_wdata1_3 : _GEN_18339; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18341 = 7'h4 == index[6:0] ? recent_wdata1_4 : _GEN_18340; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18342 = 7'h5 == index[6:0] ? recent_wdata1_5 : _GEN_18341; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18343 = 7'h6 == index[6:0] ? recent_wdata1_6 : _GEN_18342; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18344 = 7'h7 == index[6:0] ? recent_wdata1_7 : _GEN_18343; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18345 = 7'h8 == index[6:0] ? recent_wdata1_8 : _GEN_18344; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18346 = 7'h9 == index[6:0] ? recent_wdata1_9 : _GEN_18345; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18347 = 7'ha == index[6:0] ? recent_wdata1_10 : _GEN_18346; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18348 = 7'hb == index[6:0] ? recent_wdata1_11 : _GEN_18347; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18349 = 7'hc == index[6:0] ? recent_wdata1_12 : _GEN_18348; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18350 = 7'hd == index[6:0] ? recent_wdata1_13 : _GEN_18349; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18351 = 7'he == index[6:0] ? recent_wdata1_14 : _GEN_18350; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18352 = 7'hf == index[6:0] ? recent_wdata1_15 : _GEN_18351; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18353 = 7'h10 == index[6:0] ? recent_wdata1_16 : _GEN_18352; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18354 = 7'h11 == index[6:0] ? recent_wdata1_17 : _GEN_18353; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18355 = 7'h12 == index[6:0] ? recent_wdata1_18 : _GEN_18354; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18356 = 7'h13 == index[6:0] ? recent_wdata1_19 : _GEN_18355; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18357 = 7'h14 == index[6:0] ? recent_wdata1_20 : _GEN_18356; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18358 = 7'h15 == index[6:0] ? recent_wdata1_21 : _GEN_18357; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18359 = 7'h16 == index[6:0] ? recent_wdata1_22 : _GEN_18358; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18360 = 7'h17 == index[6:0] ? recent_wdata1_23 : _GEN_18359; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18361 = 7'h18 == index[6:0] ? recent_wdata1_24 : _GEN_18360; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18362 = 7'h19 == index[6:0] ? recent_wdata1_25 : _GEN_18361; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18363 = 7'h1a == index[6:0] ? recent_wdata1_26 : _GEN_18362; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18364 = 7'h1b == index[6:0] ? recent_wdata1_27 : _GEN_18363; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18365 = 7'h1c == index[6:0] ? recent_wdata1_28 : _GEN_18364; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18366 = 7'h1d == index[6:0] ? recent_wdata1_29 : _GEN_18365; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18367 = 7'h1e == index[6:0] ? recent_wdata1_30 : _GEN_18366; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18368 = 7'h1f == index[6:0] ? recent_wdata1_31 : _GEN_18367; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18369 = 7'h20 == index[6:0] ? recent_wdata1_32 : _GEN_18368; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18370 = 7'h21 == index[6:0] ? recent_wdata1_33 : _GEN_18369; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18371 = 7'h22 == index[6:0] ? recent_wdata1_34 : _GEN_18370; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18372 = 7'h23 == index[6:0] ? recent_wdata1_35 : _GEN_18371; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18373 = 7'h24 == index[6:0] ? recent_wdata1_36 : _GEN_18372; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18374 = 7'h25 == index[6:0] ? recent_wdata1_37 : _GEN_18373; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18375 = 7'h26 == index[6:0] ? recent_wdata1_38 : _GEN_18374; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18376 = 7'h27 == index[6:0] ? recent_wdata1_39 : _GEN_18375; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18377 = 7'h28 == index[6:0] ? recent_wdata1_40 : _GEN_18376; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18378 = 7'h29 == index[6:0] ? recent_wdata1_41 : _GEN_18377; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18379 = 7'h2a == index[6:0] ? recent_wdata1_42 : _GEN_18378; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18380 = 7'h2b == index[6:0] ? recent_wdata1_43 : _GEN_18379; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18381 = 7'h2c == index[6:0] ? recent_wdata1_44 : _GEN_18380; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18382 = 7'h2d == index[6:0] ? recent_wdata1_45 : _GEN_18381; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18383 = 7'h2e == index[6:0] ? recent_wdata1_46 : _GEN_18382; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18384 = 7'h2f == index[6:0] ? recent_wdata1_47 : _GEN_18383; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18385 = 7'h30 == index[6:0] ? recent_wdata1_48 : _GEN_18384; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18386 = 7'h31 == index[6:0] ? recent_wdata1_49 : _GEN_18385; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18387 = 7'h32 == index[6:0] ? recent_wdata1_50 : _GEN_18386; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18388 = 7'h33 == index[6:0] ? recent_wdata1_51 : _GEN_18387; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18389 = 7'h34 == index[6:0] ? recent_wdata1_52 : _GEN_18388; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18390 = 7'h35 == index[6:0] ? recent_wdata1_53 : _GEN_18389; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18391 = 7'h36 == index[6:0] ? recent_wdata1_54 : _GEN_18390; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18392 = 7'h37 == index[6:0] ? recent_wdata1_55 : _GEN_18391; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18393 = 7'h38 == index[6:0] ? recent_wdata1_56 : _GEN_18392; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18394 = 7'h39 == index[6:0] ? recent_wdata1_57 : _GEN_18393; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18395 = 7'h3a == index[6:0] ? recent_wdata1_58 : _GEN_18394; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18396 = 7'h3b == index[6:0] ? recent_wdata1_59 : _GEN_18395; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18397 = 7'h3c == index[6:0] ? recent_wdata1_60 : _GEN_18396; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18398 = 7'h3d == index[6:0] ? recent_wdata1_61 : _GEN_18397; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18399 = 7'h3e == index[6:0] ? recent_wdata1_62 : _GEN_18398; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18400 = 7'h3f == index[6:0] ? recent_wdata1_63 : _GEN_18399; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18401 = 7'h40 == index[6:0] ? recent_wdata1_64 : _GEN_18400; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18402 = 7'h41 == index[6:0] ? recent_wdata1_65 : _GEN_18401; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18403 = 7'h42 == index[6:0] ? recent_wdata1_66 : _GEN_18402; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18404 = 7'h43 == index[6:0] ? recent_wdata1_67 : _GEN_18403; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18405 = 7'h44 == index[6:0] ? recent_wdata1_68 : _GEN_18404; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18406 = 7'h45 == index[6:0] ? recent_wdata1_69 : _GEN_18405; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18407 = 7'h46 == index[6:0] ? recent_wdata1_70 : _GEN_18406; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18408 = 7'h47 == index[6:0] ? recent_wdata1_71 : _GEN_18407; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18409 = 7'h48 == index[6:0] ? recent_wdata1_72 : _GEN_18408; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18410 = 7'h49 == index[6:0] ? recent_wdata1_73 : _GEN_18409; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18411 = 7'h4a == index[6:0] ? recent_wdata1_74 : _GEN_18410; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18412 = 7'h4b == index[6:0] ? recent_wdata1_75 : _GEN_18411; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18413 = 7'h4c == index[6:0] ? recent_wdata1_76 : _GEN_18412; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18414 = 7'h4d == index[6:0] ? recent_wdata1_77 : _GEN_18413; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18415 = 7'h4e == index[6:0] ? recent_wdata1_78 : _GEN_18414; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18416 = 7'h4f == index[6:0] ? recent_wdata1_79 : _GEN_18415; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18417 = 7'h50 == index[6:0] ? recent_wdata1_80 : _GEN_18416; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18418 = 7'h51 == index[6:0] ? recent_wdata1_81 : _GEN_18417; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18419 = 7'h52 == index[6:0] ? recent_wdata1_82 : _GEN_18418; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18420 = 7'h53 == index[6:0] ? recent_wdata1_83 : _GEN_18419; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18421 = 7'h54 == index[6:0] ? recent_wdata1_84 : _GEN_18420; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18422 = 7'h55 == index[6:0] ? recent_wdata1_85 : _GEN_18421; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18423 = 7'h56 == index[6:0] ? recent_wdata1_86 : _GEN_18422; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18424 = 7'h57 == index[6:0] ? recent_wdata1_87 : _GEN_18423; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18425 = 7'h58 == index[6:0] ? recent_wdata1_88 : _GEN_18424; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18426 = 7'h59 == index[6:0] ? recent_wdata1_89 : _GEN_18425; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18427 = 7'h5a == index[6:0] ? recent_wdata1_90 : _GEN_18426; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18428 = 7'h5b == index[6:0] ? recent_wdata1_91 : _GEN_18427; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18429 = 7'h5c == index[6:0] ? recent_wdata1_92 : _GEN_18428; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18430 = 7'h5d == index[6:0] ? recent_wdata1_93 : _GEN_18429; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18431 = 7'h5e == index[6:0] ? recent_wdata1_94 : _GEN_18430; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18432 = 7'h5f == index[6:0] ? recent_wdata1_95 : _GEN_18431; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18433 = 7'h60 == index[6:0] ? recent_wdata1_96 : _GEN_18432; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18434 = 7'h61 == index[6:0] ? recent_wdata1_97 : _GEN_18433; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18435 = 7'h62 == index[6:0] ? recent_wdata1_98 : _GEN_18434; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18436 = 7'h63 == index[6:0] ? recent_wdata1_99 : _GEN_18435; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18437 = 7'h64 == index[6:0] ? recent_wdata1_100 : _GEN_18436; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18438 = 7'h65 == index[6:0] ? recent_wdata1_101 : _GEN_18437; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18439 = 7'h66 == index[6:0] ? recent_wdata1_102 : _GEN_18438; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18440 = 7'h67 == index[6:0] ? recent_wdata1_103 : _GEN_18439; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18441 = 7'h68 == index[6:0] ? recent_wdata1_104 : _GEN_18440; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18442 = 7'h69 == index[6:0] ? recent_wdata1_105 : _GEN_18441; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18443 = 7'h6a == index[6:0] ? recent_wdata1_106 : _GEN_18442; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18444 = 7'h6b == index[6:0] ? recent_wdata1_107 : _GEN_18443; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18445 = 7'h6c == index[6:0] ? recent_wdata1_108 : _GEN_18444; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18446 = 7'h6d == index[6:0] ? recent_wdata1_109 : _GEN_18445; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18447 = 7'h6e == index[6:0] ? recent_wdata1_110 : _GEN_18446; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18448 = 7'h6f == index[6:0] ? recent_wdata1_111 : _GEN_18447; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18449 = 7'h70 == index[6:0] ? recent_wdata1_112 : _GEN_18448; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18450 = 7'h71 == index[6:0] ? recent_wdata1_113 : _GEN_18449; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18451 = 7'h72 == index[6:0] ? recent_wdata1_114 : _GEN_18450; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18452 = 7'h73 == index[6:0] ? recent_wdata1_115 : _GEN_18451; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18453 = 7'h74 == index[6:0] ? recent_wdata1_116 : _GEN_18452; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18454 = 7'h75 == index[6:0] ? recent_wdata1_117 : _GEN_18453; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18455 = 7'h76 == index[6:0] ? recent_wdata1_118 : _GEN_18454; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18456 = 7'h77 == index[6:0] ? recent_wdata1_119 : _GEN_18455; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18457 = 7'h78 == index[6:0] ? recent_wdata1_120 : _GEN_18456; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18458 = 7'h79 == index[6:0] ? recent_wdata1_121 : _GEN_18457; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18459 = 7'h7a == index[6:0] ? recent_wdata1_122 : _GEN_18458; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18460 = 7'h7b == index[6:0] ? recent_wdata1_123 : _GEN_18459; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18461 = 7'h7c == index[6:0] ? recent_wdata1_124 : _GEN_18460; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18462 = 7'h7d == index[6:0] ? recent_wdata1_125 : _GEN_18461; // @[d_cache.scala 363:{11,11}]
  wire [63:0] _GEN_18463 = 7'h7e == index[6:0] ? recent_wdata1_126 : _GEN_18462; // @[d_cache.scala 363:{11,11}]
  wire [41:0] _GEN_19500 = reset ? 42'h0 : _GEN_17600; // @[d_cache.scala 32:{34,34}]
  wire  _GEN_19502 = ~_T_20 & _T_21; // @[d_cache.scala 93:27]
  assign io_to_lsu_arready = state == 3'h0 ? io_from_axi_arready : _GEN_17933; // @[d_cache.scala 199:23 201:27]
  assign io_to_lsu_rdata = state == 3'h0 ? 64'h0 : _GEN_17932; // @[d_cache.scala 199:23 200:25]
  assign io_to_lsu_rvalid = state == 3'h0 ? 1'h0 : _GEN_17934; // @[d_cache.scala 199:23 202:26]
  assign io_to_lsu_awready = state == 3'h0 ? io_from_axi_awready : _GEN_17936; // @[d_cache.scala 199:23 205:27]
  assign io_to_lsu_wready = state == 3'h0 ? 1'h0 : _GEN_17935; // @[d_cache.scala 199:23 203:26]
  assign io_to_lsu_bvalid = state == 3'h0 ? 1'h0 : _GEN_17937; // @[d_cache.scala 199:23 204:26]
  assign io_to_axi_araddr = _GEN_17945[31:0];
  assign io_to_axi_arvalid = state == 3'h0 ? 1'h0 : _GEN_17923; // @[d_cache.scala 199:23 206:27]
  assign io_to_axi_rready = state == 3'h0 ? io_from_lsu_rready : _GEN_17925; // @[d_cache.scala 199:23 208:26]
  assign io_to_axi_awaddr = state == 3'h0 ? 32'h0 : _GEN_17926; // @[d_cache.scala 199:23 209:26]
  assign io_to_axi_awvalid = state == 3'h0 ? 1'h0 : _GEN_17927; // @[d_cache.scala 199:23 210:27]
  assign io_to_axi_wdata = _GEN_17949[31:0];
  assign io_to_axi_wstrb = state == 3'h0 ? 8'h0 : _GEN_17929; // @[d_cache.scala 199:23 212:25]
  assign io_to_axi_wvalid = state == 3'h0 ? 1'h0 : _GEN_17930; // @[d_cache.scala 199:23 213:26]
  assign io_to_axi_bready = state == 3'h0 ? io_from_lsu_bready : _GEN_17931; // @[d_cache.scala 199:23 214:26]
  always @(posedge clock) begin
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_0 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_0 <= _GEN_2443;
        end else begin
          ram_0_0 <= _GEN_12719;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_1 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_1 <= _GEN_2444;
        end else begin
          ram_0_1 <= _GEN_12720;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_2 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_2 <= _GEN_2445;
        end else begin
          ram_0_2 <= _GEN_12721;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_3 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_3 <= _GEN_2446;
        end else begin
          ram_0_3 <= _GEN_12722;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_4 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_4 <= _GEN_2447;
        end else begin
          ram_0_4 <= _GEN_12723;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_5 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_5 <= _GEN_2448;
        end else begin
          ram_0_5 <= _GEN_12724;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_6 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_6 <= _GEN_2449;
        end else begin
          ram_0_6 <= _GEN_12725;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_7 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_7 <= _GEN_2450;
        end else begin
          ram_0_7 <= _GEN_12726;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_8 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_8 <= _GEN_2451;
        end else begin
          ram_0_8 <= _GEN_12727;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_9 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_9 <= _GEN_2452;
        end else begin
          ram_0_9 <= _GEN_12728;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_10 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_10 <= _GEN_2453;
        end else begin
          ram_0_10 <= _GEN_12729;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_11 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_11 <= _GEN_2454;
        end else begin
          ram_0_11 <= _GEN_12730;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_12 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_12 <= _GEN_2455;
        end else begin
          ram_0_12 <= _GEN_12731;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_13 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_13 <= _GEN_2456;
        end else begin
          ram_0_13 <= _GEN_12732;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_14 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_14 <= _GEN_2457;
        end else begin
          ram_0_14 <= _GEN_12733;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_15 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_15 <= _GEN_2458;
        end else begin
          ram_0_15 <= _GEN_12734;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_16 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_16 <= _GEN_2459;
        end else begin
          ram_0_16 <= _GEN_12735;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_17 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_17 <= _GEN_2460;
        end else begin
          ram_0_17 <= _GEN_12736;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_18 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_18 <= _GEN_2461;
        end else begin
          ram_0_18 <= _GEN_12737;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_19 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_19 <= _GEN_2462;
        end else begin
          ram_0_19 <= _GEN_12738;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_20 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_20 <= _GEN_2463;
        end else begin
          ram_0_20 <= _GEN_12739;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_21 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_21 <= _GEN_2464;
        end else begin
          ram_0_21 <= _GEN_12740;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_22 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_22 <= _GEN_2465;
        end else begin
          ram_0_22 <= _GEN_12741;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_23 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_23 <= _GEN_2466;
        end else begin
          ram_0_23 <= _GEN_12742;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_24 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_24 <= _GEN_2467;
        end else begin
          ram_0_24 <= _GEN_12743;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_25 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_25 <= _GEN_2468;
        end else begin
          ram_0_25 <= _GEN_12744;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_26 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_26 <= _GEN_2469;
        end else begin
          ram_0_26 <= _GEN_12745;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_27 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_27 <= _GEN_2470;
        end else begin
          ram_0_27 <= _GEN_12746;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_28 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_28 <= _GEN_2471;
        end else begin
          ram_0_28 <= _GEN_12747;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_29 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_29 <= _GEN_2472;
        end else begin
          ram_0_29 <= _GEN_12748;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_30 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_30 <= _GEN_2473;
        end else begin
          ram_0_30 <= _GEN_12749;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_31 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_31 <= _GEN_2474;
        end else begin
          ram_0_31 <= _GEN_12750;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_32 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_32 <= _GEN_2475;
        end else begin
          ram_0_32 <= _GEN_12751;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_33 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_33 <= _GEN_2476;
        end else begin
          ram_0_33 <= _GEN_12752;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_34 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_34 <= _GEN_2477;
        end else begin
          ram_0_34 <= _GEN_12753;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_35 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_35 <= _GEN_2478;
        end else begin
          ram_0_35 <= _GEN_12754;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_36 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_36 <= _GEN_2479;
        end else begin
          ram_0_36 <= _GEN_12755;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_37 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_37 <= _GEN_2480;
        end else begin
          ram_0_37 <= _GEN_12756;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_38 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_38 <= _GEN_2481;
        end else begin
          ram_0_38 <= _GEN_12757;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_39 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_39 <= _GEN_2482;
        end else begin
          ram_0_39 <= _GEN_12758;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_40 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_40 <= _GEN_2483;
        end else begin
          ram_0_40 <= _GEN_12759;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_41 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_41 <= _GEN_2484;
        end else begin
          ram_0_41 <= _GEN_12760;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_42 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_42 <= _GEN_2485;
        end else begin
          ram_0_42 <= _GEN_12761;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_43 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_43 <= _GEN_2486;
        end else begin
          ram_0_43 <= _GEN_12762;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_44 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_44 <= _GEN_2487;
        end else begin
          ram_0_44 <= _GEN_12763;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_45 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_45 <= _GEN_2488;
        end else begin
          ram_0_45 <= _GEN_12764;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_46 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_46 <= _GEN_2489;
        end else begin
          ram_0_46 <= _GEN_12765;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_47 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_47 <= _GEN_2490;
        end else begin
          ram_0_47 <= _GEN_12766;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_48 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_48 <= _GEN_2491;
        end else begin
          ram_0_48 <= _GEN_12767;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_49 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_49 <= _GEN_2492;
        end else begin
          ram_0_49 <= _GEN_12768;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_50 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_50 <= _GEN_2493;
        end else begin
          ram_0_50 <= _GEN_12769;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_51 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_51 <= _GEN_2494;
        end else begin
          ram_0_51 <= _GEN_12770;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_52 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_52 <= _GEN_2495;
        end else begin
          ram_0_52 <= _GEN_12771;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_53 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_53 <= _GEN_2496;
        end else begin
          ram_0_53 <= _GEN_12772;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_54 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_54 <= _GEN_2497;
        end else begin
          ram_0_54 <= _GEN_12773;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_55 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_55 <= _GEN_2498;
        end else begin
          ram_0_55 <= _GEN_12774;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_56 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_56 <= _GEN_2499;
        end else begin
          ram_0_56 <= _GEN_12775;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_57 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_57 <= _GEN_2500;
        end else begin
          ram_0_57 <= _GEN_12776;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_58 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_58 <= _GEN_2501;
        end else begin
          ram_0_58 <= _GEN_12777;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_59 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_59 <= _GEN_2502;
        end else begin
          ram_0_59 <= _GEN_12778;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_60 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_60 <= _GEN_2503;
        end else begin
          ram_0_60 <= _GEN_12779;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_61 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_61 <= _GEN_2504;
        end else begin
          ram_0_61 <= _GEN_12780;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_62 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_62 <= _GEN_2505;
        end else begin
          ram_0_62 <= _GEN_12781;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_63 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_63 <= _GEN_2506;
        end else begin
          ram_0_63 <= _GEN_12782;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_64 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_64 <= _GEN_2507;
        end else begin
          ram_0_64 <= _GEN_12783;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_65 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_65 <= _GEN_2508;
        end else begin
          ram_0_65 <= _GEN_12784;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_66 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_66 <= _GEN_2509;
        end else begin
          ram_0_66 <= _GEN_12785;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_67 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_67 <= _GEN_2510;
        end else begin
          ram_0_67 <= _GEN_12786;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_68 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_68 <= _GEN_2511;
        end else begin
          ram_0_68 <= _GEN_12787;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_69 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_69 <= _GEN_2512;
        end else begin
          ram_0_69 <= _GEN_12788;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_70 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_70 <= _GEN_2513;
        end else begin
          ram_0_70 <= _GEN_12789;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_71 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_71 <= _GEN_2514;
        end else begin
          ram_0_71 <= _GEN_12790;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_72 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_72 <= _GEN_2515;
        end else begin
          ram_0_72 <= _GEN_12791;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_73 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_73 <= _GEN_2516;
        end else begin
          ram_0_73 <= _GEN_12792;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_74 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_74 <= _GEN_2517;
        end else begin
          ram_0_74 <= _GEN_12793;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_75 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_75 <= _GEN_2518;
        end else begin
          ram_0_75 <= _GEN_12794;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_76 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_76 <= _GEN_2519;
        end else begin
          ram_0_76 <= _GEN_12795;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_77 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_77 <= _GEN_2520;
        end else begin
          ram_0_77 <= _GEN_12796;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_78 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_78 <= _GEN_2521;
        end else begin
          ram_0_78 <= _GEN_12797;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_79 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_79 <= _GEN_2522;
        end else begin
          ram_0_79 <= _GEN_12798;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_80 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_80 <= _GEN_2523;
        end else begin
          ram_0_80 <= _GEN_12799;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_81 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_81 <= _GEN_2524;
        end else begin
          ram_0_81 <= _GEN_12800;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_82 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_82 <= _GEN_2525;
        end else begin
          ram_0_82 <= _GEN_12801;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_83 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_83 <= _GEN_2526;
        end else begin
          ram_0_83 <= _GEN_12802;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_84 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_84 <= _GEN_2527;
        end else begin
          ram_0_84 <= _GEN_12803;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_85 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_85 <= _GEN_2528;
        end else begin
          ram_0_85 <= _GEN_12804;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_86 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_86 <= _GEN_2529;
        end else begin
          ram_0_86 <= _GEN_12805;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_87 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_87 <= _GEN_2530;
        end else begin
          ram_0_87 <= _GEN_12806;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_88 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_88 <= _GEN_2531;
        end else begin
          ram_0_88 <= _GEN_12807;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_89 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_89 <= _GEN_2532;
        end else begin
          ram_0_89 <= _GEN_12808;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_90 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_90 <= _GEN_2533;
        end else begin
          ram_0_90 <= _GEN_12809;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_91 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_91 <= _GEN_2534;
        end else begin
          ram_0_91 <= _GEN_12810;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_92 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_92 <= _GEN_2535;
        end else begin
          ram_0_92 <= _GEN_12811;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_93 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_93 <= _GEN_2536;
        end else begin
          ram_0_93 <= _GEN_12812;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_94 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_94 <= _GEN_2537;
        end else begin
          ram_0_94 <= _GEN_12813;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_95 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_95 <= _GEN_2538;
        end else begin
          ram_0_95 <= _GEN_12814;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_96 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_96 <= _GEN_2539;
        end else begin
          ram_0_96 <= _GEN_12815;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_97 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_97 <= _GEN_2540;
        end else begin
          ram_0_97 <= _GEN_12816;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_98 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_98 <= _GEN_2541;
        end else begin
          ram_0_98 <= _GEN_12817;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_99 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_99 <= _GEN_2542;
        end else begin
          ram_0_99 <= _GEN_12818;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_100 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_100 <= _GEN_2543;
        end else begin
          ram_0_100 <= _GEN_12819;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_101 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_101 <= _GEN_2544;
        end else begin
          ram_0_101 <= _GEN_12820;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_102 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_102 <= _GEN_2545;
        end else begin
          ram_0_102 <= _GEN_12821;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_103 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_103 <= _GEN_2546;
        end else begin
          ram_0_103 <= _GEN_12822;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_104 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_104 <= _GEN_2547;
        end else begin
          ram_0_104 <= _GEN_12823;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_105 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_105 <= _GEN_2548;
        end else begin
          ram_0_105 <= _GEN_12824;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_106 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_106 <= _GEN_2549;
        end else begin
          ram_0_106 <= _GEN_12825;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_107 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_107 <= _GEN_2550;
        end else begin
          ram_0_107 <= _GEN_12826;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_108 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_108 <= _GEN_2551;
        end else begin
          ram_0_108 <= _GEN_12827;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_109 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_109 <= _GEN_2552;
        end else begin
          ram_0_109 <= _GEN_12828;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_110 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_110 <= _GEN_2553;
        end else begin
          ram_0_110 <= _GEN_12829;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_111 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_111 <= _GEN_2554;
        end else begin
          ram_0_111 <= _GEN_12830;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_112 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_112 <= _GEN_2555;
        end else begin
          ram_0_112 <= _GEN_12831;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_113 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_113 <= _GEN_2556;
        end else begin
          ram_0_113 <= _GEN_12832;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_114 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_114 <= _GEN_2557;
        end else begin
          ram_0_114 <= _GEN_12833;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_115 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_115 <= _GEN_2558;
        end else begin
          ram_0_115 <= _GEN_12834;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_116 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_116 <= _GEN_2559;
        end else begin
          ram_0_116 <= _GEN_12835;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_117 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_117 <= _GEN_2560;
        end else begin
          ram_0_117 <= _GEN_12836;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_118 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_118 <= _GEN_2561;
        end else begin
          ram_0_118 <= _GEN_12837;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_119 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_119 <= _GEN_2562;
        end else begin
          ram_0_119 <= _GEN_12838;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_120 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_120 <= _GEN_2563;
        end else begin
          ram_0_120 <= _GEN_12839;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_121 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_121 <= _GEN_2564;
        end else begin
          ram_0_121 <= _GEN_12840;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_122 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_122 <= _GEN_2565;
        end else begin
          ram_0_122 <= _GEN_12841;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_123 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_123 <= _GEN_2566;
        end else begin
          ram_0_123 <= _GEN_12842;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_124 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_124 <= _GEN_2567;
        end else begin
          ram_0_124 <= _GEN_12843;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_125 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_125 <= _GEN_2568;
        end else begin
          ram_0_125 <= _GEN_12844;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_126 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_126 <= _GEN_2569;
        end else begin
          ram_0_126 <= _GEN_12845;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_127 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_127 <= _GEN_2570;
        end else begin
          ram_0_127 <= _GEN_12846;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_0 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_0 <= _GEN_2827;
        end else begin
          ram_1_0 <= _GEN_13104;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_1 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_1 <= _GEN_2828;
        end else begin
          ram_1_1 <= _GEN_13105;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_2 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_2 <= _GEN_2829;
        end else begin
          ram_1_2 <= _GEN_13106;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_3 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_3 <= _GEN_2830;
        end else begin
          ram_1_3 <= _GEN_13107;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_4 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_4 <= _GEN_2831;
        end else begin
          ram_1_4 <= _GEN_13108;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_5 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_5 <= _GEN_2832;
        end else begin
          ram_1_5 <= _GEN_13109;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_6 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_6 <= _GEN_2833;
        end else begin
          ram_1_6 <= _GEN_13110;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_7 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_7 <= _GEN_2834;
        end else begin
          ram_1_7 <= _GEN_13111;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_8 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_8 <= _GEN_2835;
        end else begin
          ram_1_8 <= _GEN_13112;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_9 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_9 <= _GEN_2836;
        end else begin
          ram_1_9 <= _GEN_13113;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_10 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_10 <= _GEN_2837;
        end else begin
          ram_1_10 <= _GEN_13114;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_11 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_11 <= _GEN_2838;
        end else begin
          ram_1_11 <= _GEN_13115;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_12 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_12 <= _GEN_2839;
        end else begin
          ram_1_12 <= _GEN_13116;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_13 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_13 <= _GEN_2840;
        end else begin
          ram_1_13 <= _GEN_13117;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_14 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_14 <= _GEN_2841;
        end else begin
          ram_1_14 <= _GEN_13118;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_15 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_15 <= _GEN_2842;
        end else begin
          ram_1_15 <= _GEN_13119;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_16 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_16 <= _GEN_2843;
        end else begin
          ram_1_16 <= _GEN_13120;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_17 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_17 <= _GEN_2844;
        end else begin
          ram_1_17 <= _GEN_13121;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_18 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_18 <= _GEN_2845;
        end else begin
          ram_1_18 <= _GEN_13122;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_19 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_19 <= _GEN_2846;
        end else begin
          ram_1_19 <= _GEN_13123;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_20 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_20 <= _GEN_2847;
        end else begin
          ram_1_20 <= _GEN_13124;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_21 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_21 <= _GEN_2848;
        end else begin
          ram_1_21 <= _GEN_13125;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_22 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_22 <= _GEN_2849;
        end else begin
          ram_1_22 <= _GEN_13126;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_23 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_23 <= _GEN_2850;
        end else begin
          ram_1_23 <= _GEN_13127;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_24 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_24 <= _GEN_2851;
        end else begin
          ram_1_24 <= _GEN_13128;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_25 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_25 <= _GEN_2852;
        end else begin
          ram_1_25 <= _GEN_13129;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_26 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_26 <= _GEN_2853;
        end else begin
          ram_1_26 <= _GEN_13130;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_27 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_27 <= _GEN_2854;
        end else begin
          ram_1_27 <= _GEN_13131;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_28 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_28 <= _GEN_2855;
        end else begin
          ram_1_28 <= _GEN_13132;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_29 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_29 <= _GEN_2856;
        end else begin
          ram_1_29 <= _GEN_13133;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_30 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_30 <= _GEN_2857;
        end else begin
          ram_1_30 <= _GEN_13134;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_31 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_31 <= _GEN_2858;
        end else begin
          ram_1_31 <= _GEN_13135;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_32 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_32 <= _GEN_2859;
        end else begin
          ram_1_32 <= _GEN_13136;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_33 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_33 <= _GEN_2860;
        end else begin
          ram_1_33 <= _GEN_13137;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_34 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_34 <= _GEN_2861;
        end else begin
          ram_1_34 <= _GEN_13138;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_35 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_35 <= _GEN_2862;
        end else begin
          ram_1_35 <= _GEN_13139;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_36 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_36 <= _GEN_2863;
        end else begin
          ram_1_36 <= _GEN_13140;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_37 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_37 <= _GEN_2864;
        end else begin
          ram_1_37 <= _GEN_13141;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_38 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_38 <= _GEN_2865;
        end else begin
          ram_1_38 <= _GEN_13142;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_39 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_39 <= _GEN_2866;
        end else begin
          ram_1_39 <= _GEN_13143;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_40 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_40 <= _GEN_2867;
        end else begin
          ram_1_40 <= _GEN_13144;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_41 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_41 <= _GEN_2868;
        end else begin
          ram_1_41 <= _GEN_13145;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_42 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_42 <= _GEN_2869;
        end else begin
          ram_1_42 <= _GEN_13146;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_43 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_43 <= _GEN_2870;
        end else begin
          ram_1_43 <= _GEN_13147;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_44 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_44 <= _GEN_2871;
        end else begin
          ram_1_44 <= _GEN_13148;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_45 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_45 <= _GEN_2872;
        end else begin
          ram_1_45 <= _GEN_13149;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_46 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_46 <= _GEN_2873;
        end else begin
          ram_1_46 <= _GEN_13150;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_47 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_47 <= _GEN_2874;
        end else begin
          ram_1_47 <= _GEN_13151;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_48 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_48 <= _GEN_2875;
        end else begin
          ram_1_48 <= _GEN_13152;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_49 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_49 <= _GEN_2876;
        end else begin
          ram_1_49 <= _GEN_13153;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_50 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_50 <= _GEN_2877;
        end else begin
          ram_1_50 <= _GEN_13154;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_51 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_51 <= _GEN_2878;
        end else begin
          ram_1_51 <= _GEN_13155;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_52 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_52 <= _GEN_2879;
        end else begin
          ram_1_52 <= _GEN_13156;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_53 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_53 <= _GEN_2880;
        end else begin
          ram_1_53 <= _GEN_13157;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_54 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_54 <= _GEN_2881;
        end else begin
          ram_1_54 <= _GEN_13158;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_55 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_55 <= _GEN_2882;
        end else begin
          ram_1_55 <= _GEN_13159;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_56 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_56 <= _GEN_2883;
        end else begin
          ram_1_56 <= _GEN_13160;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_57 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_57 <= _GEN_2884;
        end else begin
          ram_1_57 <= _GEN_13161;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_58 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_58 <= _GEN_2885;
        end else begin
          ram_1_58 <= _GEN_13162;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_59 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_59 <= _GEN_2886;
        end else begin
          ram_1_59 <= _GEN_13163;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_60 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_60 <= _GEN_2887;
        end else begin
          ram_1_60 <= _GEN_13164;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_61 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_61 <= _GEN_2888;
        end else begin
          ram_1_61 <= _GEN_13165;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_62 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_62 <= _GEN_2889;
        end else begin
          ram_1_62 <= _GEN_13166;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_63 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_63 <= _GEN_2890;
        end else begin
          ram_1_63 <= _GEN_13167;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_64 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_64 <= _GEN_2891;
        end else begin
          ram_1_64 <= _GEN_13168;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_65 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_65 <= _GEN_2892;
        end else begin
          ram_1_65 <= _GEN_13169;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_66 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_66 <= _GEN_2893;
        end else begin
          ram_1_66 <= _GEN_13170;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_67 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_67 <= _GEN_2894;
        end else begin
          ram_1_67 <= _GEN_13171;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_68 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_68 <= _GEN_2895;
        end else begin
          ram_1_68 <= _GEN_13172;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_69 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_69 <= _GEN_2896;
        end else begin
          ram_1_69 <= _GEN_13173;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_70 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_70 <= _GEN_2897;
        end else begin
          ram_1_70 <= _GEN_13174;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_71 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_71 <= _GEN_2898;
        end else begin
          ram_1_71 <= _GEN_13175;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_72 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_72 <= _GEN_2899;
        end else begin
          ram_1_72 <= _GEN_13176;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_73 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_73 <= _GEN_2900;
        end else begin
          ram_1_73 <= _GEN_13177;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_74 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_74 <= _GEN_2901;
        end else begin
          ram_1_74 <= _GEN_13178;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_75 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_75 <= _GEN_2902;
        end else begin
          ram_1_75 <= _GEN_13179;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_76 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_76 <= _GEN_2903;
        end else begin
          ram_1_76 <= _GEN_13180;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_77 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_77 <= _GEN_2904;
        end else begin
          ram_1_77 <= _GEN_13181;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_78 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_78 <= _GEN_2905;
        end else begin
          ram_1_78 <= _GEN_13182;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_79 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_79 <= _GEN_2906;
        end else begin
          ram_1_79 <= _GEN_13183;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_80 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_80 <= _GEN_2907;
        end else begin
          ram_1_80 <= _GEN_13184;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_81 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_81 <= _GEN_2908;
        end else begin
          ram_1_81 <= _GEN_13185;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_82 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_82 <= _GEN_2909;
        end else begin
          ram_1_82 <= _GEN_13186;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_83 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_83 <= _GEN_2910;
        end else begin
          ram_1_83 <= _GEN_13187;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_84 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_84 <= _GEN_2911;
        end else begin
          ram_1_84 <= _GEN_13188;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_85 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_85 <= _GEN_2912;
        end else begin
          ram_1_85 <= _GEN_13189;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_86 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_86 <= _GEN_2913;
        end else begin
          ram_1_86 <= _GEN_13190;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_87 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_87 <= _GEN_2914;
        end else begin
          ram_1_87 <= _GEN_13191;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_88 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_88 <= _GEN_2915;
        end else begin
          ram_1_88 <= _GEN_13192;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_89 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_89 <= _GEN_2916;
        end else begin
          ram_1_89 <= _GEN_13193;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_90 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_90 <= _GEN_2917;
        end else begin
          ram_1_90 <= _GEN_13194;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_91 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_91 <= _GEN_2918;
        end else begin
          ram_1_91 <= _GEN_13195;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_92 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_92 <= _GEN_2919;
        end else begin
          ram_1_92 <= _GEN_13196;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_93 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_93 <= _GEN_2920;
        end else begin
          ram_1_93 <= _GEN_13197;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_94 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_94 <= _GEN_2921;
        end else begin
          ram_1_94 <= _GEN_13198;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_95 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_95 <= _GEN_2922;
        end else begin
          ram_1_95 <= _GEN_13199;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_96 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_96 <= _GEN_2923;
        end else begin
          ram_1_96 <= _GEN_13200;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_97 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_97 <= _GEN_2924;
        end else begin
          ram_1_97 <= _GEN_13201;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_98 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_98 <= _GEN_2925;
        end else begin
          ram_1_98 <= _GEN_13202;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_99 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_99 <= _GEN_2926;
        end else begin
          ram_1_99 <= _GEN_13203;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_100 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_100 <= _GEN_2927;
        end else begin
          ram_1_100 <= _GEN_13204;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_101 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_101 <= _GEN_2928;
        end else begin
          ram_1_101 <= _GEN_13205;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_102 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_102 <= _GEN_2929;
        end else begin
          ram_1_102 <= _GEN_13206;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_103 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_103 <= _GEN_2930;
        end else begin
          ram_1_103 <= _GEN_13207;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_104 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_104 <= _GEN_2931;
        end else begin
          ram_1_104 <= _GEN_13208;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_105 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_105 <= _GEN_2932;
        end else begin
          ram_1_105 <= _GEN_13209;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_106 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_106 <= _GEN_2933;
        end else begin
          ram_1_106 <= _GEN_13210;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_107 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_107 <= _GEN_2934;
        end else begin
          ram_1_107 <= _GEN_13211;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_108 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_108 <= _GEN_2935;
        end else begin
          ram_1_108 <= _GEN_13212;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_109 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_109 <= _GEN_2936;
        end else begin
          ram_1_109 <= _GEN_13213;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_110 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_110 <= _GEN_2937;
        end else begin
          ram_1_110 <= _GEN_13214;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_111 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_111 <= _GEN_2938;
        end else begin
          ram_1_111 <= _GEN_13215;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_112 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_112 <= _GEN_2939;
        end else begin
          ram_1_112 <= _GEN_13216;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_113 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_113 <= _GEN_2940;
        end else begin
          ram_1_113 <= _GEN_13217;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_114 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_114 <= _GEN_2941;
        end else begin
          ram_1_114 <= _GEN_13218;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_115 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_115 <= _GEN_2942;
        end else begin
          ram_1_115 <= _GEN_13219;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_116 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_116 <= _GEN_2943;
        end else begin
          ram_1_116 <= _GEN_13220;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_117 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_117 <= _GEN_2944;
        end else begin
          ram_1_117 <= _GEN_13221;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_118 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_118 <= _GEN_2945;
        end else begin
          ram_1_118 <= _GEN_13222;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_119 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_119 <= _GEN_2946;
        end else begin
          ram_1_119 <= _GEN_13223;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_120 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_120 <= _GEN_2947;
        end else begin
          ram_1_120 <= _GEN_13224;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_121 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_121 <= _GEN_2948;
        end else begin
          ram_1_121 <= _GEN_13225;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_122 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_122 <= _GEN_2949;
        end else begin
          ram_1_122 <= _GEN_13226;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_123 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_123 <= _GEN_2950;
        end else begin
          ram_1_123 <= _GEN_13227;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_124 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_124 <= _GEN_2951;
        end else begin
          ram_1_124 <= _GEN_13228;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_125 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_125 <= _GEN_2952;
        end else begin
          ram_1_125 <= _GEN_13229;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_126 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_126 <= _GEN_2953;
        end else begin
          ram_1_126 <= _GEN_13230;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_127 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_127 <= _GEN_2954;
        end else begin
          ram_1_127 <= _GEN_13231;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_0 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_0 <= _GEN_2571;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_1 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_1 <= _GEN_2572;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_2 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_2 <= _GEN_2573;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_3 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_3 <= _GEN_2574;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_4 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_4 <= _GEN_2575;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_5 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_5 <= _GEN_2576;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_6 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_6 <= _GEN_2577;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_7 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_7 <= _GEN_2578;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_8 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_8 <= _GEN_2579;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_9 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_9 <= _GEN_2580;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_10 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_10 <= _GEN_2581;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_11 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_11 <= _GEN_2582;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_12 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_12 <= _GEN_2583;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_13 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_13 <= _GEN_2584;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_14 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_14 <= _GEN_2585;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_15 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_15 <= _GEN_2586;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_16 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_16 <= _GEN_2587;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_17 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_17 <= _GEN_2588;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_18 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_18 <= _GEN_2589;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_19 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_19 <= _GEN_2590;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_20 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_20 <= _GEN_2591;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_21 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_21 <= _GEN_2592;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_22 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_22 <= _GEN_2593;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_23 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_23 <= _GEN_2594;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_24 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_24 <= _GEN_2595;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_25 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_25 <= _GEN_2596;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_26 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_26 <= _GEN_2597;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_27 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_27 <= _GEN_2598;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_28 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_28 <= _GEN_2599;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_29 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_29 <= _GEN_2600;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_30 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_30 <= _GEN_2601;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_31 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_31 <= _GEN_2602;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_32 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_32 <= _GEN_2603;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_33 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_33 <= _GEN_2604;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_34 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_34 <= _GEN_2605;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_35 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_35 <= _GEN_2606;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_36 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_36 <= _GEN_2607;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_37 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_37 <= _GEN_2608;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_38 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_38 <= _GEN_2609;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_39 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_39 <= _GEN_2610;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_40 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_40 <= _GEN_2611;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_41 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_41 <= _GEN_2612;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_42 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_42 <= _GEN_2613;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_43 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_43 <= _GEN_2614;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_44 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_44 <= _GEN_2615;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_45 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_45 <= _GEN_2616;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_46 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_46 <= _GEN_2617;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_47 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_47 <= _GEN_2618;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_48 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_48 <= _GEN_2619;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_49 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_49 <= _GEN_2620;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_50 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_50 <= _GEN_2621;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_51 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_51 <= _GEN_2622;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_52 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_52 <= _GEN_2623;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_53 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_53 <= _GEN_2624;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_54 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_54 <= _GEN_2625;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_55 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_55 <= _GEN_2626;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_56 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_56 <= _GEN_2627;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_57 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_57 <= _GEN_2628;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_58 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_58 <= _GEN_2629;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_59 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_59 <= _GEN_2630;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_60 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_60 <= _GEN_2631;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_61 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_61 <= _GEN_2632;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_62 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_62 <= _GEN_2633;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_63 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_63 <= _GEN_2634;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_64 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_64 <= _GEN_2635;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_65 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_65 <= _GEN_2636;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_66 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_66 <= _GEN_2637;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_67 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_67 <= _GEN_2638;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_68 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_68 <= _GEN_2639;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_69 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_69 <= _GEN_2640;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_70 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_70 <= _GEN_2641;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_71 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_71 <= _GEN_2642;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_72 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_72 <= _GEN_2643;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_73 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_73 <= _GEN_2644;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_74 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_74 <= _GEN_2645;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_75 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_75 <= _GEN_2646;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_76 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_76 <= _GEN_2647;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_77 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_77 <= _GEN_2648;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_78 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_78 <= _GEN_2649;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_79 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_79 <= _GEN_2650;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_80 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_80 <= _GEN_2651;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_81 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_81 <= _GEN_2652;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_82 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_82 <= _GEN_2653;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_83 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_83 <= _GEN_2654;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_84 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_84 <= _GEN_2655;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_85 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_85 <= _GEN_2656;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_86 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_86 <= _GEN_2657;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_87 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_87 <= _GEN_2658;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_88 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_88 <= _GEN_2659;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_89 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_89 <= _GEN_2660;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_90 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_90 <= _GEN_2661;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_91 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_91 <= _GEN_2662;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_92 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_92 <= _GEN_2663;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_93 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_93 <= _GEN_2664;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_94 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_94 <= _GEN_2665;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_95 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_95 <= _GEN_2666;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_96 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_96 <= _GEN_2667;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_97 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_97 <= _GEN_2668;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_98 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_98 <= _GEN_2669;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_99 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_99 <= _GEN_2670;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_100 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_100 <= _GEN_2671;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_101 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_101 <= _GEN_2672;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_102 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_102 <= _GEN_2673;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_103 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_103 <= _GEN_2674;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_104 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_104 <= _GEN_2675;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_105 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_105 <= _GEN_2676;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_106 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_106 <= _GEN_2677;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_107 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_107 <= _GEN_2678;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_108 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_108 <= _GEN_2679;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_109 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_109 <= _GEN_2680;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_110 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_110 <= _GEN_2681;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_111 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_111 <= _GEN_2682;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_112 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_112 <= _GEN_2683;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_113 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_113 <= _GEN_2684;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_114 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_114 <= _GEN_2685;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_115 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_115 <= _GEN_2686;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_116 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_116 <= _GEN_2687;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_117 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_117 <= _GEN_2688;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_118 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_118 <= _GEN_2689;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_119 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_119 <= _GEN_2690;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_120 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_120 <= _GEN_2691;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_121 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_121 <= _GEN_2692;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_122 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_122 <= _GEN_2693;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_123 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_123 <= _GEN_2694;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_124 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_124 <= _GEN_2695;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_125 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_125 <= _GEN_2696;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_126 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_126 <= _GEN_2697;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:32]
      recent_wdata0_127 <= 64'h0; // @[d_cache.scala 20:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata0_127 <= _GEN_2698;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_0 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_0 <= _GEN_2955;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_1 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_1 <= _GEN_2956;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_2 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_2 <= _GEN_2957;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_3 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_3 <= _GEN_2958;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_4 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_4 <= _GEN_2959;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_5 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_5 <= _GEN_2960;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_6 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_6 <= _GEN_2961;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_7 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_7 <= _GEN_2962;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_8 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_8 <= _GEN_2963;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_9 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_9 <= _GEN_2964;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_10 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_10 <= _GEN_2965;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_11 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_11 <= _GEN_2966;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_12 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_12 <= _GEN_2967;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_13 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_13 <= _GEN_2968;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_14 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_14 <= _GEN_2969;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_15 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_15 <= _GEN_2970;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_16 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_16 <= _GEN_2971;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_17 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_17 <= _GEN_2972;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_18 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_18 <= _GEN_2973;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_19 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_19 <= _GEN_2974;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_20 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_20 <= _GEN_2975;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_21 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_21 <= _GEN_2976;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_22 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_22 <= _GEN_2977;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_23 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_23 <= _GEN_2978;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_24 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_24 <= _GEN_2979;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_25 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_25 <= _GEN_2980;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_26 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_26 <= _GEN_2981;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_27 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_27 <= _GEN_2982;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_28 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_28 <= _GEN_2983;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_29 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_29 <= _GEN_2984;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_30 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_30 <= _GEN_2985;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_31 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_31 <= _GEN_2986;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_32 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_32 <= _GEN_2987;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_33 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_33 <= _GEN_2988;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_34 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_34 <= _GEN_2989;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_35 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_35 <= _GEN_2990;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_36 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_36 <= _GEN_2991;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_37 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_37 <= _GEN_2992;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_38 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_38 <= _GEN_2993;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_39 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_39 <= _GEN_2994;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_40 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_40 <= _GEN_2995;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_41 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_41 <= _GEN_2996;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_42 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_42 <= _GEN_2997;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_43 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_43 <= _GEN_2998;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_44 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_44 <= _GEN_2999;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_45 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_45 <= _GEN_3000;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_46 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_46 <= _GEN_3001;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_47 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_47 <= _GEN_3002;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_48 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_48 <= _GEN_3003;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_49 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_49 <= _GEN_3004;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_50 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_50 <= _GEN_3005;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_51 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_51 <= _GEN_3006;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_52 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_52 <= _GEN_3007;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_53 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_53 <= _GEN_3008;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_54 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_54 <= _GEN_3009;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_55 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_55 <= _GEN_3010;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_56 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_56 <= _GEN_3011;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_57 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_57 <= _GEN_3012;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_58 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_58 <= _GEN_3013;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_59 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_59 <= _GEN_3014;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_60 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_60 <= _GEN_3015;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_61 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_61 <= _GEN_3016;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_62 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_62 <= _GEN_3017;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_63 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_63 <= _GEN_3018;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_64 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_64 <= _GEN_3019;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_65 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_65 <= _GEN_3020;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_66 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_66 <= _GEN_3021;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_67 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_67 <= _GEN_3022;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_68 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_68 <= _GEN_3023;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_69 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_69 <= _GEN_3024;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_70 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_70 <= _GEN_3025;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_71 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_71 <= _GEN_3026;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_72 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_72 <= _GEN_3027;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_73 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_73 <= _GEN_3028;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_74 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_74 <= _GEN_3029;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_75 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_75 <= _GEN_3030;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_76 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_76 <= _GEN_3031;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_77 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_77 <= _GEN_3032;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_78 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_78 <= _GEN_3033;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_79 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_79 <= _GEN_3034;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_80 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_80 <= _GEN_3035;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_81 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_81 <= _GEN_3036;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_82 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_82 <= _GEN_3037;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_83 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_83 <= _GEN_3038;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_84 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_84 <= _GEN_3039;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_85 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_85 <= _GEN_3040;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_86 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_86 <= _GEN_3041;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_87 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_87 <= _GEN_3042;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_88 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_88 <= _GEN_3043;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_89 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_89 <= _GEN_3044;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_90 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_90 <= _GEN_3045;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_91 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_91 <= _GEN_3046;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_92 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_92 <= _GEN_3047;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_93 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_93 <= _GEN_3048;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_94 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_94 <= _GEN_3049;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_95 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_95 <= _GEN_3050;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_96 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_96 <= _GEN_3051;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_97 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_97 <= _GEN_3052;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_98 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_98 <= _GEN_3053;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_99 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_99 <= _GEN_3054;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_100 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_100 <= _GEN_3055;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_101 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_101 <= _GEN_3056;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_102 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_102 <= _GEN_3057;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_103 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_103 <= _GEN_3058;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_104 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_104 <= _GEN_3059;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_105 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_105 <= _GEN_3060;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_106 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_106 <= _GEN_3061;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_107 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_107 <= _GEN_3062;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_108 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_108 <= _GEN_3063;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_109 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_109 <= _GEN_3064;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_110 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_110 <= _GEN_3065;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_111 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_111 <= _GEN_3066;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_112 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_112 <= _GEN_3067;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_113 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_113 <= _GEN_3068;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_114 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_114 <= _GEN_3069;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_115 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_115 <= _GEN_3070;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_116 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_116 <= _GEN_3071;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_117 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_117 <= _GEN_3072;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_118 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_118 <= _GEN_3073;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_119 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_119 <= _GEN_3074;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_120 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_120 <= _GEN_3075;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_121 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_121 <= _GEN_3076;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_122 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_122 <= _GEN_3077;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_123 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_123 <= _GEN_3078;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_124 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_124 <= _GEN_3079;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_125 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_125 <= _GEN_3080;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_126 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_126 <= _GEN_3081;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      recent_wdata1_127 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          recent_wdata1_127 <= _GEN_3082;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_0 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_0 <= _GEN_12847;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_1 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_1 <= _GEN_12848;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_2 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_2 <= _GEN_12849;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_3 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_3 <= _GEN_12850;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_4 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_4 <= _GEN_12851;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_5 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_5 <= _GEN_12852;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_6 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_6 <= _GEN_12853;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_7 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_7 <= _GEN_12854;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_8 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_8 <= _GEN_12855;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_9 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_9 <= _GEN_12856;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_10 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_10 <= _GEN_12857;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_11 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_11 <= _GEN_12858;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_12 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_12 <= _GEN_12859;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_13 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_13 <= _GEN_12860;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_14 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_14 <= _GEN_12861;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_15 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_15 <= _GEN_12862;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_16 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_16 <= _GEN_12863;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_17 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_17 <= _GEN_12864;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_18 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_18 <= _GEN_12865;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_19 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_19 <= _GEN_12866;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_20 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_20 <= _GEN_12867;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_21 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_21 <= _GEN_12868;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_22 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_22 <= _GEN_12869;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_23 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_23 <= _GEN_12870;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_24 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_24 <= _GEN_12871;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_25 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_25 <= _GEN_12872;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_26 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_26 <= _GEN_12873;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_27 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_27 <= _GEN_12874;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_28 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_28 <= _GEN_12875;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_29 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_29 <= _GEN_12876;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_30 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_30 <= _GEN_12877;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_31 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_31 <= _GEN_12878;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_32 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_32 <= _GEN_12879;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_33 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_33 <= _GEN_12880;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_34 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_34 <= _GEN_12881;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_35 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_35 <= _GEN_12882;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_36 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_36 <= _GEN_12883;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_37 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_37 <= _GEN_12884;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_38 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_38 <= _GEN_12885;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_39 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_39 <= _GEN_12886;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_40 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_40 <= _GEN_12887;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_41 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_41 <= _GEN_12888;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_42 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_42 <= _GEN_12889;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_43 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_43 <= _GEN_12890;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_44 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_44 <= _GEN_12891;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_45 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_45 <= _GEN_12892;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_46 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_46 <= _GEN_12893;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_47 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_47 <= _GEN_12894;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_48 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_48 <= _GEN_12895;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_49 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_49 <= _GEN_12896;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_50 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_50 <= _GEN_12897;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_51 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_51 <= _GEN_12898;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_52 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_52 <= _GEN_12899;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_53 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_53 <= _GEN_12900;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_54 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_54 <= _GEN_12901;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_55 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_55 <= _GEN_12902;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_56 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_56 <= _GEN_12903;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_57 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_57 <= _GEN_12904;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_58 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_58 <= _GEN_12905;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_59 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_59 <= _GEN_12906;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_60 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_60 <= _GEN_12907;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_61 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_61 <= _GEN_12908;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_62 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_62 <= _GEN_12909;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_63 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_63 <= _GEN_12910;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_64 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_64 <= _GEN_12911;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_65 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_65 <= _GEN_12912;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_66 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_66 <= _GEN_12913;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_67 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_67 <= _GEN_12914;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_68 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_68 <= _GEN_12915;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_69 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_69 <= _GEN_12916;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_70 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_70 <= _GEN_12917;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_71 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_71 <= _GEN_12918;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_72 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_72 <= _GEN_12919;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_73 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_73 <= _GEN_12920;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_74 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_74 <= _GEN_12921;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_75 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_75 <= _GEN_12922;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_76 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_76 <= _GEN_12923;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_77 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_77 <= _GEN_12924;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_78 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_78 <= _GEN_12925;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_79 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_79 <= _GEN_12926;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_80 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_80 <= _GEN_12927;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_81 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_81 <= _GEN_12928;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_82 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_82 <= _GEN_12929;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_83 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_83 <= _GEN_12930;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_84 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_84 <= _GEN_12931;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_85 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_85 <= _GEN_12932;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_86 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_86 <= _GEN_12933;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_87 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_87 <= _GEN_12934;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_88 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_88 <= _GEN_12935;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_89 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_89 <= _GEN_12936;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_90 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_90 <= _GEN_12937;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_91 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_91 <= _GEN_12938;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_92 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_92 <= _GEN_12939;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_93 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_93 <= _GEN_12940;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_94 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_94 <= _GEN_12941;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_95 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_95 <= _GEN_12942;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_96 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_96 <= _GEN_12943;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_97 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_97 <= _GEN_12944;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_98 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_98 <= _GEN_12945;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_99 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_99 <= _GEN_12946;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_100 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_100 <= _GEN_12947;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_101 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_101 <= _GEN_12948;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_102 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_102 <= _GEN_12949;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_103 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_103 <= _GEN_12950;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_104 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_104 <= _GEN_12951;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_105 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_105 <= _GEN_12952;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_106 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_106 <= _GEN_12953;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_107 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_107 <= _GEN_12954;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_108 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_108 <= _GEN_12955;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_109 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_109 <= _GEN_12956;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_110 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_110 <= _GEN_12957;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_111 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_111 <= _GEN_12958;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_112 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_112 <= _GEN_12959;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_113 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_113 <= _GEN_12960;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_114 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_114 <= _GEN_12961;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_115 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_115 <= _GEN_12962;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_116 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_116 <= _GEN_12963;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_117 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_117 <= _GEN_12964;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_118 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_118 <= _GEN_12965;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_119 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_119 <= _GEN_12966;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_120 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_120 <= _GEN_12967;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_121 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_121 <= _GEN_12968;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_122 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_122 <= _GEN_12969;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_123 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_123 <= _GEN_12970;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_124 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_124 <= _GEN_12971;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_125 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_125 <= _GEN_12972;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_126 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_126 <= _GEN_12973;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_127 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_127 <= _GEN_12974;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_0 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_0 <= _GEN_13232;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_1 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_1 <= _GEN_13233;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_2 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_2 <= _GEN_13234;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_3 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_3 <= _GEN_13235;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_4 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_4 <= _GEN_13236;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_5 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_5 <= _GEN_13237;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_6 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_6 <= _GEN_13238;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_7 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_7 <= _GEN_13239;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_8 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_8 <= _GEN_13240;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_9 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_9 <= _GEN_13241;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_10 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_10 <= _GEN_13242;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_11 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_11 <= _GEN_13243;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_12 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_12 <= _GEN_13244;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_13 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_13 <= _GEN_13245;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_14 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_14 <= _GEN_13246;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_15 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_15 <= _GEN_13247;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_16 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_16 <= _GEN_13248;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_17 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_17 <= _GEN_13249;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_18 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_18 <= _GEN_13250;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_19 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_19 <= _GEN_13251;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_20 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_20 <= _GEN_13252;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_21 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_21 <= _GEN_13253;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_22 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_22 <= _GEN_13254;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_23 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_23 <= _GEN_13255;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_24 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_24 <= _GEN_13256;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_25 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_25 <= _GEN_13257;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_26 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_26 <= _GEN_13258;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_27 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_27 <= _GEN_13259;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_28 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_28 <= _GEN_13260;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_29 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_29 <= _GEN_13261;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_30 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_30 <= _GEN_13262;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_31 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_31 <= _GEN_13263;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_32 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_32 <= _GEN_13264;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_33 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_33 <= _GEN_13265;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_34 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_34 <= _GEN_13266;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_35 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_35 <= _GEN_13267;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_36 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_36 <= _GEN_13268;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_37 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_37 <= _GEN_13269;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_38 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_38 <= _GEN_13270;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_39 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_39 <= _GEN_13271;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_40 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_40 <= _GEN_13272;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_41 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_41 <= _GEN_13273;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_42 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_42 <= _GEN_13274;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_43 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_43 <= _GEN_13275;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_44 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_44 <= _GEN_13276;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_45 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_45 <= _GEN_13277;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_46 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_46 <= _GEN_13278;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_47 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_47 <= _GEN_13279;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_48 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_48 <= _GEN_13280;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_49 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_49 <= _GEN_13281;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_50 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_50 <= _GEN_13282;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_51 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_51 <= _GEN_13283;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_52 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_52 <= _GEN_13284;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_53 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_53 <= _GEN_13285;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_54 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_54 <= _GEN_13286;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_55 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_55 <= _GEN_13287;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_56 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_56 <= _GEN_13288;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_57 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_57 <= _GEN_13289;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_58 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_58 <= _GEN_13290;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_59 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_59 <= _GEN_13291;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_60 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_60 <= _GEN_13292;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_61 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_61 <= _GEN_13293;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_62 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_62 <= _GEN_13294;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_63 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_63 <= _GEN_13295;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_64 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_64 <= _GEN_13296;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_65 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_65 <= _GEN_13297;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_66 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_66 <= _GEN_13298;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_67 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_67 <= _GEN_13299;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_68 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_68 <= _GEN_13300;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_69 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_69 <= _GEN_13301;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_70 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_70 <= _GEN_13302;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_71 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_71 <= _GEN_13303;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_72 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_72 <= _GEN_13304;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_73 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_73 <= _GEN_13305;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_74 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_74 <= _GEN_13306;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_75 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_75 <= _GEN_13307;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_76 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_76 <= _GEN_13308;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_77 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_77 <= _GEN_13309;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_78 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_78 <= _GEN_13310;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_79 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_79 <= _GEN_13311;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_80 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_80 <= _GEN_13312;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_81 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_81 <= _GEN_13313;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_82 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_82 <= _GEN_13314;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_83 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_83 <= _GEN_13315;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_84 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_84 <= _GEN_13316;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_85 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_85 <= _GEN_13317;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_86 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_86 <= _GEN_13318;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_87 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_87 <= _GEN_13319;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_88 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_88 <= _GEN_13320;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_89 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_89 <= _GEN_13321;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_90 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_90 <= _GEN_13322;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_91 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_91 <= _GEN_13323;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_92 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_92 <= _GEN_13324;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_93 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_93 <= _GEN_13325;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_94 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_94 <= _GEN_13326;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_95 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_95 <= _GEN_13327;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_96 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_96 <= _GEN_13328;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_97 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_97 <= _GEN_13329;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_98 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_98 <= _GEN_13330;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_99 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_99 <= _GEN_13331;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_100 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_100 <= _GEN_13332;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_101 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_101 <= _GEN_13333;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_102 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_102 <= _GEN_13334;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_103 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_103 <= _GEN_13335;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_104 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_104 <= _GEN_13336;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_105 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_105 <= _GEN_13337;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_106 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_106 <= _GEN_13338;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_107 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_107 <= _GEN_13339;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_108 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_108 <= _GEN_13340;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_109 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_109 <= _GEN_13341;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_110 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_110 <= _GEN_13342;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_111 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_111 <= _GEN_13343;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_112 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_112 <= _GEN_13344;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_113 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_113 <= _GEN_13345;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_114 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_114 <= _GEN_13346;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_115 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_115 <= _GEN_13347;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_116 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_116 <= _GEN_13348;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_117 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_117 <= _GEN_13349;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_118 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_118 <= _GEN_13350;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_119 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_119 <= _GEN_13351;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_120 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_120 <= _GEN_13352;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_121 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_121 <= _GEN_13353;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_122 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_122 <= _GEN_13354;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_123 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_123 <= _GEN_13355;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_124 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_124 <= _GEN_13356;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_125 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_125 <= _GEN_13357;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_126 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_126 <= _GEN_13358;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_127 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_127 <= _GEN_13359;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_0 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_0 <= _GEN_12975;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_1 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_1 <= _GEN_12976;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_2 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_2 <= _GEN_12977;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_3 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_3 <= _GEN_12978;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_4 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_4 <= _GEN_12979;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_5 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_5 <= _GEN_12980;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_6 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_6 <= _GEN_12981;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_7 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_7 <= _GEN_12982;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_8 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_8 <= _GEN_12983;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_9 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_9 <= _GEN_12984;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_10 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_10 <= _GEN_12985;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_11 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_11 <= _GEN_12986;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_12 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_12 <= _GEN_12987;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_13 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_13 <= _GEN_12988;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_14 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_14 <= _GEN_12989;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_15 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_15 <= _GEN_12990;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_16 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_16 <= _GEN_12991;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_17 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_17 <= _GEN_12992;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_18 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_18 <= _GEN_12993;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_19 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_19 <= _GEN_12994;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_20 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_20 <= _GEN_12995;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_21 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_21 <= _GEN_12996;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_22 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_22 <= _GEN_12997;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_23 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_23 <= _GEN_12998;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_24 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_24 <= _GEN_12999;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_25 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_25 <= _GEN_13000;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_26 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_26 <= _GEN_13001;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_27 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_27 <= _GEN_13002;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_28 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_28 <= _GEN_13003;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_29 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_29 <= _GEN_13004;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_30 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_30 <= _GEN_13005;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_31 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_31 <= _GEN_13006;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_32 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_32 <= _GEN_13007;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_33 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_33 <= _GEN_13008;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_34 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_34 <= _GEN_13009;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_35 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_35 <= _GEN_13010;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_36 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_36 <= _GEN_13011;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_37 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_37 <= _GEN_13012;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_38 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_38 <= _GEN_13013;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_39 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_39 <= _GEN_13014;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_40 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_40 <= _GEN_13015;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_41 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_41 <= _GEN_13016;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_42 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_42 <= _GEN_13017;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_43 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_43 <= _GEN_13018;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_44 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_44 <= _GEN_13019;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_45 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_45 <= _GEN_13020;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_46 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_46 <= _GEN_13021;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_47 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_47 <= _GEN_13022;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_48 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_48 <= _GEN_13023;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_49 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_49 <= _GEN_13024;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_50 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_50 <= _GEN_13025;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_51 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_51 <= _GEN_13026;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_52 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_52 <= _GEN_13027;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_53 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_53 <= _GEN_13028;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_54 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_54 <= _GEN_13029;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_55 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_55 <= _GEN_13030;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_56 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_56 <= _GEN_13031;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_57 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_57 <= _GEN_13032;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_58 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_58 <= _GEN_13033;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_59 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_59 <= _GEN_13034;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_60 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_60 <= _GEN_13035;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_61 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_61 <= _GEN_13036;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_62 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_62 <= _GEN_13037;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_63 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_63 <= _GEN_13038;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_64 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_64 <= _GEN_13039;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_65 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_65 <= _GEN_13040;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_66 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_66 <= _GEN_13041;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_67 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_67 <= _GEN_13042;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_68 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_68 <= _GEN_13043;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_69 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_69 <= _GEN_13044;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_70 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_70 <= _GEN_13045;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_71 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_71 <= _GEN_13046;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_72 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_72 <= _GEN_13047;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_73 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_73 <= _GEN_13048;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_74 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_74 <= _GEN_13049;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_75 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_75 <= _GEN_13050;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_76 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_76 <= _GEN_13051;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_77 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_77 <= _GEN_13052;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_78 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_78 <= _GEN_13053;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_79 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_79 <= _GEN_13054;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_80 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_80 <= _GEN_13055;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_81 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_81 <= _GEN_13056;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_82 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_82 <= _GEN_13057;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_83 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_83 <= _GEN_13058;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_84 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_84 <= _GEN_13059;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_85 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_85 <= _GEN_13060;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_86 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_86 <= _GEN_13061;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_87 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_87 <= _GEN_13062;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_88 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_88 <= _GEN_13063;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_89 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_89 <= _GEN_13064;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_90 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_90 <= _GEN_13065;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_91 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_91 <= _GEN_13066;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_92 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_92 <= _GEN_13067;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_93 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_93 <= _GEN_13068;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_94 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_94 <= _GEN_13069;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_95 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_95 <= _GEN_13070;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_96 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_96 <= _GEN_13071;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_97 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_97 <= _GEN_13072;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_98 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_98 <= _GEN_13073;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_99 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_99 <= _GEN_13074;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_100 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_100 <= _GEN_13075;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_101 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_101 <= _GEN_13076;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_102 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_102 <= _GEN_13077;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_103 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_103 <= _GEN_13078;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_104 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_104 <= _GEN_13079;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_105 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_105 <= _GEN_13080;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_106 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_106 <= _GEN_13081;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_107 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_107 <= _GEN_13082;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_108 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_108 <= _GEN_13083;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_109 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_109 <= _GEN_13084;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_110 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_110 <= _GEN_13085;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_111 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_111 <= _GEN_13086;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_112 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_112 <= _GEN_13087;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_113 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_113 <= _GEN_13088;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_114 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_114 <= _GEN_13089;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_115 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_115 <= _GEN_13090;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_116 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_116 <= _GEN_13091;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_117 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_117 <= _GEN_13092;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_118 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_118 <= _GEN_13093;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_119 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_119 <= _GEN_13094;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_120 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_120 <= _GEN_13095;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_121 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_121 <= _GEN_13096;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_122 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_122 <= _GEN_13097;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_123 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_123 <= _GEN_13098;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_124 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_124 <= _GEN_13099;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_125 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_125 <= _GEN_13100;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_126 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_126 <= _GEN_13101;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_127 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_0_127 <= _GEN_13102;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_0 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_0 <= _GEN_13360;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_1 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_1 <= _GEN_13361;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_2 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_2 <= _GEN_13362;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_3 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_3 <= _GEN_13363;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_4 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_4 <= _GEN_13364;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_5 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_5 <= _GEN_13365;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_6 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_6 <= _GEN_13366;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_7 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_7 <= _GEN_13367;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_8 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_8 <= _GEN_13368;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_9 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_9 <= _GEN_13369;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_10 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_10 <= _GEN_13370;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_11 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_11 <= _GEN_13371;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_12 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_12 <= _GEN_13372;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_13 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_13 <= _GEN_13373;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_14 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_14 <= _GEN_13374;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_15 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_15 <= _GEN_13375;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_16 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_16 <= _GEN_13376;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_17 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_17 <= _GEN_13377;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_18 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_18 <= _GEN_13378;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_19 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_19 <= _GEN_13379;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_20 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_20 <= _GEN_13380;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_21 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_21 <= _GEN_13381;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_22 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_22 <= _GEN_13382;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_23 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_23 <= _GEN_13383;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_24 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_24 <= _GEN_13384;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_25 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_25 <= _GEN_13385;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_26 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_26 <= _GEN_13386;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_27 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_27 <= _GEN_13387;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_28 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_28 <= _GEN_13388;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_29 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_29 <= _GEN_13389;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_30 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_30 <= _GEN_13390;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_31 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_31 <= _GEN_13391;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_32 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_32 <= _GEN_13392;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_33 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_33 <= _GEN_13393;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_34 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_34 <= _GEN_13394;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_35 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_35 <= _GEN_13395;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_36 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_36 <= _GEN_13396;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_37 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_37 <= _GEN_13397;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_38 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_38 <= _GEN_13398;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_39 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_39 <= _GEN_13399;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_40 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_40 <= _GEN_13400;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_41 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_41 <= _GEN_13401;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_42 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_42 <= _GEN_13402;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_43 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_43 <= _GEN_13403;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_44 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_44 <= _GEN_13404;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_45 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_45 <= _GEN_13405;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_46 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_46 <= _GEN_13406;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_47 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_47 <= _GEN_13407;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_48 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_48 <= _GEN_13408;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_49 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_49 <= _GEN_13409;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_50 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_50 <= _GEN_13410;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_51 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_51 <= _GEN_13411;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_52 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_52 <= _GEN_13412;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_53 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_53 <= _GEN_13413;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_54 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_54 <= _GEN_13414;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_55 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_55 <= _GEN_13415;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_56 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_56 <= _GEN_13416;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_57 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_57 <= _GEN_13417;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_58 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_58 <= _GEN_13418;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_59 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_59 <= _GEN_13419;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_60 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_60 <= _GEN_13420;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_61 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_61 <= _GEN_13421;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_62 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_62 <= _GEN_13422;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_63 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_63 <= _GEN_13423;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_64 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_64 <= _GEN_13424;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_65 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_65 <= _GEN_13425;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_66 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_66 <= _GEN_13426;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_67 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_67 <= _GEN_13427;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_68 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_68 <= _GEN_13428;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_69 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_69 <= _GEN_13429;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_70 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_70 <= _GEN_13430;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_71 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_71 <= _GEN_13431;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_72 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_72 <= _GEN_13432;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_73 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_73 <= _GEN_13433;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_74 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_74 <= _GEN_13434;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_75 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_75 <= _GEN_13435;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_76 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_76 <= _GEN_13436;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_77 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_77 <= _GEN_13437;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_78 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_78 <= _GEN_13438;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_79 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_79 <= _GEN_13439;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_80 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_80 <= _GEN_13440;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_81 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_81 <= _GEN_13441;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_82 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_82 <= _GEN_13442;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_83 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_83 <= _GEN_13443;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_84 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_84 <= _GEN_13444;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_85 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_85 <= _GEN_13445;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_86 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_86 <= _GEN_13446;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_87 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_87 <= _GEN_13447;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_88 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_88 <= _GEN_13448;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_89 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_89 <= _GEN_13449;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_90 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_90 <= _GEN_13450;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_91 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_91 <= _GEN_13451;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_92 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_92 <= _GEN_13452;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_93 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_93 <= _GEN_13453;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_94 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_94 <= _GEN_13454;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_95 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_95 <= _GEN_13455;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_96 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_96 <= _GEN_13456;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_97 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_97 <= _GEN_13457;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_98 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_98 <= _GEN_13458;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_99 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_99 <= _GEN_13459;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_100 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_100 <= _GEN_13460;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_101 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_101 <= _GEN_13461;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_102 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_102 <= _GEN_13462;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_103 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_103 <= _GEN_13463;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_104 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_104 <= _GEN_13464;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_105 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_105 <= _GEN_13465;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_106 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_106 <= _GEN_13466;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_107 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_107 <= _GEN_13467;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_108 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_108 <= _GEN_13468;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_109 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_109 <= _GEN_13469;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_110 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_110 <= _GEN_13470;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_111 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_111 <= _GEN_13471;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_112 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_112 <= _GEN_13472;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_113 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_113 <= _GEN_13473;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_114 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_114 <= _GEN_13474;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_115 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_115 <= _GEN_13475;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_116 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_116 <= _GEN_13476;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_117 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_117 <= _GEN_13477;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_118 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_118 <= _GEN_13478;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_119 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_119 <= _GEN_13479;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_120 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_120 <= _GEN_13480;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_121 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_121 <= _GEN_13481;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_122 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_122 <= _GEN_13482;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_123 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_123 <= _GEN_13483;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_124 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_124 <= _GEN_13484;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_125 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_125 <= _GEN_13485;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_126 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_126 <= _GEN_13486;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_127 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          valid_1_127 <= _GEN_13487;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_0 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_0 <= _GEN_2699;
        end else begin
          dirty_0_0 <= _GEN_13490;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_1 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_1 <= _GEN_2700;
        end else begin
          dirty_0_1 <= _GEN_13491;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_2 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_2 <= _GEN_2701;
        end else begin
          dirty_0_2 <= _GEN_13492;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_3 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_3 <= _GEN_2702;
        end else begin
          dirty_0_3 <= _GEN_13493;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_4 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_4 <= _GEN_2703;
        end else begin
          dirty_0_4 <= _GEN_13494;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_5 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_5 <= _GEN_2704;
        end else begin
          dirty_0_5 <= _GEN_13495;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_6 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_6 <= _GEN_2705;
        end else begin
          dirty_0_6 <= _GEN_13496;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_7 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_7 <= _GEN_2706;
        end else begin
          dirty_0_7 <= _GEN_13497;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_8 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_8 <= _GEN_2707;
        end else begin
          dirty_0_8 <= _GEN_13498;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_9 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_9 <= _GEN_2708;
        end else begin
          dirty_0_9 <= _GEN_13499;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_10 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_10 <= _GEN_2709;
        end else begin
          dirty_0_10 <= _GEN_13500;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_11 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_11 <= _GEN_2710;
        end else begin
          dirty_0_11 <= _GEN_13501;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_12 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_12 <= _GEN_2711;
        end else begin
          dirty_0_12 <= _GEN_13502;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_13 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_13 <= _GEN_2712;
        end else begin
          dirty_0_13 <= _GEN_13503;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_14 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_14 <= _GEN_2713;
        end else begin
          dirty_0_14 <= _GEN_13504;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_15 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_15 <= _GEN_2714;
        end else begin
          dirty_0_15 <= _GEN_13505;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_16 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_16 <= _GEN_2715;
        end else begin
          dirty_0_16 <= _GEN_13506;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_17 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_17 <= _GEN_2716;
        end else begin
          dirty_0_17 <= _GEN_13507;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_18 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_18 <= _GEN_2717;
        end else begin
          dirty_0_18 <= _GEN_13508;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_19 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_19 <= _GEN_2718;
        end else begin
          dirty_0_19 <= _GEN_13509;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_20 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_20 <= _GEN_2719;
        end else begin
          dirty_0_20 <= _GEN_13510;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_21 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_21 <= _GEN_2720;
        end else begin
          dirty_0_21 <= _GEN_13511;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_22 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_22 <= _GEN_2721;
        end else begin
          dirty_0_22 <= _GEN_13512;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_23 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_23 <= _GEN_2722;
        end else begin
          dirty_0_23 <= _GEN_13513;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_24 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_24 <= _GEN_2723;
        end else begin
          dirty_0_24 <= _GEN_13514;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_25 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_25 <= _GEN_2724;
        end else begin
          dirty_0_25 <= _GEN_13515;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_26 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_26 <= _GEN_2725;
        end else begin
          dirty_0_26 <= _GEN_13516;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_27 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_27 <= _GEN_2726;
        end else begin
          dirty_0_27 <= _GEN_13517;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_28 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_28 <= _GEN_2727;
        end else begin
          dirty_0_28 <= _GEN_13518;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_29 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_29 <= _GEN_2728;
        end else begin
          dirty_0_29 <= _GEN_13519;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_30 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_30 <= _GEN_2729;
        end else begin
          dirty_0_30 <= _GEN_13520;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_31 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_31 <= _GEN_2730;
        end else begin
          dirty_0_31 <= _GEN_13521;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_32 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_32 <= _GEN_2731;
        end else begin
          dirty_0_32 <= _GEN_13522;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_33 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_33 <= _GEN_2732;
        end else begin
          dirty_0_33 <= _GEN_13523;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_34 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_34 <= _GEN_2733;
        end else begin
          dirty_0_34 <= _GEN_13524;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_35 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_35 <= _GEN_2734;
        end else begin
          dirty_0_35 <= _GEN_13525;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_36 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_36 <= _GEN_2735;
        end else begin
          dirty_0_36 <= _GEN_13526;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_37 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_37 <= _GEN_2736;
        end else begin
          dirty_0_37 <= _GEN_13527;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_38 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_38 <= _GEN_2737;
        end else begin
          dirty_0_38 <= _GEN_13528;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_39 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_39 <= _GEN_2738;
        end else begin
          dirty_0_39 <= _GEN_13529;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_40 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_40 <= _GEN_2739;
        end else begin
          dirty_0_40 <= _GEN_13530;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_41 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_41 <= _GEN_2740;
        end else begin
          dirty_0_41 <= _GEN_13531;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_42 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_42 <= _GEN_2741;
        end else begin
          dirty_0_42 <= _GEN_13532;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_43 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_43 <= _GEN_2742;
        end else begin
          dirty_0_43 <= _GEN_13533;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_44 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_44 <= _GEN_2743;
        end else begin
          dirty_0_44 <= _GEN_13534;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_45 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_45 <= _GEN_2744;
        end else begin
          dirty_0_45 <= _GEN_13535;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_46 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_46 <= _GEN_2745;
        end else begin
          dirty_0_46 <= _GEN_13536;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_47 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_47 <= _GEN_2746;
        end else begin
          dirty_0_47 <= _GEN_13537;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_48 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_48 <= _GEN_2747;
        end else begin
          dirty_0_48 <= _GEN_13538;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_49 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_49 <= _GEN_2748;
        end else begin
          dirty_0_49 <= _GEN_13539;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_50 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_50 <= _GEN_2749;
        end else begin
          dirty_0_50 <= _GEN_13540;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_51 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_51 <= _GEN_2750;
        end else begin
          dirty_0_51 <= _GEN_13541;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_52 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_52 <= _GEN_2751;
        end else begin
          dirty_0_52 <= _GEN_13542;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_53 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_53 <= _GEN_2752;
        end else begin
          dirty_0_53 <= _GEN_13543;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_54 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_54 <= _GEN_2753;
        end else begin
          dirty_0_54 <= _GEN_13544;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_55 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_55 <= _GEN_2754;
        end else begin
          dirty_0_55 <= _GEN_13545;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_56 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_56 <= _GEN_2755;
        end else begin
          dirty_0_56 <= _GEN_13546;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_57 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_57 <= _GEN_2756;
        end else begin
          dirty_0_57 <= _GEN_13547;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_58 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_58 <= _GEN_2757;
        end else begin
          dirty_0_58 <= _GEN_13548;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_59 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_59 <= _GEN_2758;
        end else begin
          dirty_0_59 <= _GEN_13549;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_60 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_60 <= _GEN_2759;
        end else begin
          dirty_0_60 <= _GEN_13550;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_61 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_61 <= _GEN_2760;
        end else begin
          dirty_0_61 <= _GEN_13551;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_62 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_62 <= _GEN_2761;
        end else begin
          dirty_0_62 <= _GEN_13552;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_63 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_63 <= _GEN_2762;
        end else begin
          dirty_0_63 <= _GEN_13553;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_64 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_64 <= _GEN_2763;
        end else begin
          dirty_0_64 <= _GEN_13554;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_65 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_65 <= _GEN_2764;
        end else begin
          dirty_0_65 <= _GEN_13555;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_66 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_66 <= _GEN_2765;
        end else begin
          dirty_0_66 <= _GEN_13556;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_67 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_67 <= _GEN_2766;
        end else begin
          dirty_0_67 <= _GEN_13557;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_68 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_68 <= _GEN_2767;
        end else begin
          dirty_0_68 <= _GEN_13558;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_69 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_69 <= _GEN_2768;
        end else begin
          dirty_0_69 <= _GEN_13559;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_70 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_70 <= _GEN_2769;
        end else begin
          dirty_0_70 <= _GEN_13560;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_71 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_71 <= _GEN_2770;
        end else begin
          dirty_0_71 <= _GEN_13561;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_72 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_72 <= _GEN_2771;
        end else begin
          dirty_0_72 <= _GEN_13562;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_73 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_73 <= _GEN_2772;
        end else begin
          dirty_0_73 <= _GEN_13563;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_74 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_74 <= _GEN_2773;
        end else begin
          dirty_0_74 <= _GEN_13564;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_75 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_75 <= _GEN_2774;
        end else begin
          dirty_0_75 <= _GEN_13565;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_76 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_76 <= _GEN_2775;
        end else begin
          dirty_0_76 <= _GEN_13566;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_77 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_77 <= _GEN_2776;
        end else begin
          dirty_0_77 <= _GEN_13567;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_78 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_78 <= _GEN_2777;
        end else begin
          dirty_0_78 <= _GEN_13568;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_79 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_79 <= _GEN_2778;
        end else begin
          dirty_0_79 <= _GEN_13569;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_80 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_80 <= _GEN_2779;
        end else begin
          dirty_0_80 <= _GEN_13570;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_81 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_81 <= _GEN_2780;
        end else begin
          dirty_0_81 <= _GEN_13571;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_82 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_82 <= _GEN_2781;
        end else begin
          dirty_0_82 <= _GEN_13572;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_83 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_83 <= _GEN_2782;
        end else begin
          dirty_0_83 <= _GEN_13573;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_84 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_84 <= _GEN_2783;
        end else begin
          dirty_0_84 <= _GEN_13574;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_85 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_85 <= _GEN_2784;
        end else begin
          dirty_0_85 <= _GEN_13575;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_86 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_86 <= _GEN_2785;
        end else begin
          dirty_0_86 <= _GEN_13576;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_87 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_87 <= _GEN_2786;
        end else begin
          dirty_0_87 <= _GEN_13577;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_88 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_88 <= _GEN_2787;
        end else begin
          dirty_0_88 <= _GEN_13578;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_89 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_89 <= _GEN_2788;
        end else begin
          dirty_0_89 <= _GEN_13579;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_90 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_90 <= _GEN_2789;
        end else begin
          dirty_0_90 <= _GEN_13580;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_91 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_91 <= _GEN_2790;
        end else begin
          dirty_0_91 <= _GEN_13581;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_92 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_92 <= _GEN_2791;
        end else begin
          dirty_0_92 <= _GEN_13582;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_93 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_93 <= _GEN_2792;
        end else begin
          dirty_0_93 <= _GEN_13583;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_94 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_94 <= _GEN_2793;
        end else begin
          dirty_0_94 <= _GEN_13584;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_95 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_95 <= _GEN_2794;
        end else begin
          dirty_0_95 <= _GEN_13585;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_96 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_96 <= _GEN_2795;
        end else begin
          dirty_0_96 <= _GEN_13586;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_97 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_97 <= _GEN_2796;
        end else begin
          dirty_0_97 <= _GEN_13587;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_98 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_98 <= _GEN_2797;
        end else begin
          dirty_0_98 <= _GEN_13588;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_99 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_99 <= _GEN_2798;
        end else begin
          dirty_0_99 <= _GEN_13589;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_100 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_100 <= _GEN_2799;
        end else begin
          dirty_0_100 <= _GEN_13590;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_101 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_101 <= _GEN_2800;
        end else begin
          dirty_0_101 <= _GEN_13591;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_102 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_102 <= _GEN_2801;
        end else begin
          dirty_0_102 <= _GEN_13592;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_103 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_103 <= _GEN_2802;
        end else begin
          dirty_0_103 <= _GEN_13593;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_104 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_104 <= _GEN_2803;
        end else begin
          dirty_0_104 <= _GEN_13594;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_105 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_105 <= _GEN_2804;
        end else begin
          dirty_0_105 <= _GEN_13595;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_106 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_106 <= _GEN_2805;
        end else begin
          dirty_0_106 <= _GEN_13596;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_107 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_107 <= _GEN_2806;
        end else begin
          dirty_0_107 <= _GEN_13597;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_108 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_108 <= _GEN_2807;
        end else begin
          dirty_0_108 <= _GEN_13598;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_109 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_109 <= _GEN_2808;
        end else begin
          dirty_0_109 <= _GEN_13599;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_110 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_110 <= _GEN_2809;
        end else begin
          dirty_0_110 <= _GEN_13600;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_111 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_111 <= _GEN_2810;
        end else begin
          dirty_0_111 <= _GEN_13601;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_112 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_112 <= _GEN_2811;
        end else begin
          dirty_0_112 <= _GEN_13602;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_113 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_113 <= _GEN_2812;
        end else begin
          dirty_0_113 <= _GEN_13603;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_114 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_114 <= _GEN_2813;
        end else begin
          dirty_0_114 <= _GEN_13604;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_115 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_115 <= _GEN_2814;
        end else begin
          dirty_0_115 <= _GEN_13605;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_116 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_116 <= _GEN_2815;
        end else begin
          dirty_0_116 <= _GEN_13606;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_117 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_117 <= _GEN_2816;
        end else begin
          dirty_0_117 <= _GEN_13607;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_118 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_118 <= _GEN_2817;
        end else begin
          dirty_0_118 <= _GEN_13608;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_119 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_119 <= _GEN_2818;
        end else begin
          dirty_0_119 <= _GEN_13609;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_120 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_120 <= _GEN_2819;
        end else begin
          dirty_0_120 <= _GEN_13610;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_121 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_121 <= _GEN_2820;
        end else begin
          dirty_0_121 <= _GEN_13611;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_122 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_122 <= _GEN_2821;
        end else begin
          dirty_0_122 <= _GEN_13612;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_123 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_123 <= _GEN_2822;
        end else begin
          dirty_0_123 <= _GEN_13613;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_124 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_124 <= _GEN_2823;
        end else begin
          dirty_0_124 <= _GEN_13614;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_125 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_125 <= _GEN_2824;
        end else begin
          dirty_0_125 <= _GEN_13615;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_126 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_126 <= _GEN_2825;
        end else begin
          dirty_0_126 <= _GEN_13616;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_127 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_127 <= _GEN_2826;
        end else begin
          dirty_0_127 <= _GEN_13617;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_0 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_0 <= _GEN_3083;
        end else begin
          dirty_1_0 <= _GEN_13618;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_1 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_1 <= _GEN_3084;
        end else begin
          dirty_1_1 <= _GEN_13619;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_2 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_2 <= _GEN_3085;
        end else begin
          dirty_1_2 <= _GEN_13620;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_3 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_3 <= _GEN_3086;
        end else begin
          dirty_1_3 <= _GEN_13621;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_4 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_4 <= _GEN_3087;
        end else begin
          dirty_1_4 <= _GEN_13622;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_5 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_5 <= _GEN_3088;
        end else begin
          dirty_1_5 <= _GEN_13623;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_6 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_6 <= _GEN_3089;
        end else begin
          dirty_1_6 <= _GEN_13624;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_7 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_7 <= _GEN_3090;
        end else begin
          dirty_1_7 <= _GEN_13625;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_8 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_8 <= _GEN_3091;
        end else begin
          dirty_1_8 <= _GEN_13626;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_9 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_9 <= _GEN_3092;
        end else begin
          dirty_1_9 <= _GEN_13627;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_10 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_10 <= _GEN_3093;
        end else begin
          dirty_1_10 <= _GEN_13628;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_11 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_11 <= _GEN_3094;
        end else begin
          dirty_1_11 <= _GEN_13629;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_12 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_12 <= _GEN_3095;
        end else begin
          dirty_1_12 <= _GEN_13630;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_13 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_13 <= _GEN_3096;
        end else begin
          dirty_1_13 <= _GEN_13631;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_14 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_14 <= _GEN_3097;
        end else begin
          dirty_1_14 <= _GEN_13632;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_15 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_15 <= _GEN_3098;
        end else begin
          dirty_1_15 <= _GEN_13633;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_16 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_16 <= _GEN_3099;
        end else begin
          dirty_1_16 <= _GEN_13634;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_17 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_17 <= _GEN_3100;
        end else begin
          dirty_1_17 <= _GEN_13635;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_18 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_18 <= _GEN_3101;
        end else begin
          dirty_1_18 <= _GEN_13636;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_19 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_19 <= _GEN_3102;
        end else begin
          dirty_1_19 <= _GEN_13637;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_20 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_20 <= _GEN_3103;
        end else begin
          dirty_1_20 <= _GEN_13638;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_21 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_21 <= _GEN_3104;
        end else begin
          dirty_1_21 <= _GEN_13639;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_22 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_22 <= _GEN_3105;
        end else begin
          dirty_1_22 <= _GEN_13640;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_23 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_23 <= _GEN_3106;
        end else begin
          dirty_1_23 <= _GEN_13641;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_24 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_24 <= _GEN_3107;
        end else begin
          dirty_1_24 <= _GEN_13642;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_25 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_25 <= _GEN_3108;
        end else begin
          dirty_1_25 <= _GEN_13643;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_26 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_26 <= _GEN_3109;
        end else begin
          dirty_1_26 <= _GEN_13644;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_27 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_27 <= _GEN_3110;
        end else begin
          dirty_1_27 <= _GEN_13645;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_28 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_28 <= _GEN_3111;
        end else begin
          dirty_1_28 <= _GEN_13646;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_29 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_29 <= _GEN_3112;
        end else begin
          dirty_1_29 <= _GEN_13647;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_30 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_30 <= _GEN_3113;
        end else begin
          dirty_1_30 <= _GEN_13648;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_31 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_31 <= _GEN_3114;
        end else begin
          dirty_1_31 <= _GEN_13649;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_32 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_32 <= _GEN_3115;
        end else begin
          dirty_1_32 <= _GEN_13650;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_33 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_33 <= _GEN_3116;
        end else begin
          dirty_1_33 <= _GEN_13651;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_34 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_34 <= _GEN_3117;
        end else begin
          dirty_1_34 <= _GEN_13652;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_35 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_35 <= _GEN_3118;
        end else begin
          dirty_1_35 <= _GEN_13653;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_36 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_36 <= _GEN_3119;
        end else begin
          dirty_1_36 <= _GEN_13654;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_37 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_37 <= _GEN_3120;
        end else begin
          dirty_1_37 <= _GEN_13655;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_38 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_38 <= _GEN_3121;
        end else begin
          dirty_1_38 <= _GEN_13656;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_39 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_39 <= _GEN_3122;
        end else begin
          dirty_1_39 <= _GEN_13657;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_40 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_40 <= _GEN_3123;
        end else begin
          dirty_1_40 <= _GEN_13658;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_41 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_41 <= _GEN_3124;
        end else begin
          dirty_1_41 <= _GEN_13659;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_42 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_42 <= _GEN_3125;
        end else begin
          dirty_1_42 <= _GEN_13660;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_43 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_43 <= _GEN_3126;
        end else begin
          dirty_1_43 <= _GEN_13661;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_44 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_44 <= _GEN_3127;
        end else begin
          dirty_1_44 <= _GEN_13662;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_45 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_45 <= _GEN_3128;
        end else begin
          dirty_1_45 <= _GEN_13663;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_46 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_46 <= _GEN_3129;
        end else begin
          dirty_1_46 <= _GEN_13664;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_47 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_47 <= _GEN_3130;
        end else begin
          dirty_1_47 <= _GEN_13665;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_48 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_48 <= _GEN_3131;
        end else begin
          dirty_1_48 <= _GEN_13666;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_49 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_49 <= _GEN_3132;
        end else begin
          dirty_1_49 <= _GEN_13667;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_50 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_50 <= _GEN_3133;
        end else begin
          dirty_1_50 <= _GEN_13668;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_51 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_51 <= _GEN_3134;
        end else begin
          dirty_1_51 <= _GEN_13669;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_52 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_52 <= _GEN_3135;
        end else begin
          dirty_1_52 <= _GEN_13670;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_53 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_53 <= _GEN_3136;
        end else begin
          dirty_1_53 <= _GEN_13671;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_54 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_54 <= _GEN_3137;
        end else begin
          dirty_1_54 <= _GEN_13672;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_55 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_55 <= _GEN_3138;
        end else begin
          dirty_1_55 <= _GEN_13673;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_56 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_56 <= _GEN_3139;
        end else begin
          dirty_1_56 <= _GEN_13674;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_57 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_57 <= _GEN_3140;
        end else begin
          dirty_1_57 <= _GEN_13675;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_58 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_58 <= _GEN_3141;
        end else begin
          dirty_1_58 <= _GEN_13676;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_59 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_59 <= _GEN_3142;
        end else begin
          dirty_1_59 <= _GEN_13677;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_60 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_60 <= _GEN_3143;
        end else begin
          dirty_1_60 <= _GEN_13678;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_61 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_61 <= _GEN_3144;
        end else begin
          dirty_1_61 <= _GEN_13679;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_62 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_62 <= _GEN_3145;
        end else begin
          dirty_1_62 <= _GEN_13680;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_63 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_63 <= _GEN_3146;
        end else begin
          dirty_1_63 <= _GEN_13681;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_64 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_64 <= _GEN_3147;
        end else begin
          dirty_1_64 <= _GEN_13682;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_65 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_65 <= _GEN_3148;
        end else begin
          dirty_1_65 <= _GEN_13683;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_66 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_66 <= _GEN_3149;
        end else begin
          dirty_1_66 <= _GEN_13684;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_67 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_67 <= _GEN_3150;
        end else begin
          dirty_1_67 <= _GEN_13685;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_68 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_68 <= _GEN_3151;
        end else begin
          dirty_1_68 <= _GEN_13686;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_69 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_69 <= _GEN_3152;
        end else begin
          dirty_1_69 <= _GEN_13687;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_70 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_70 <= _GEN_3153;
        end else begin
          dirty_1_70 <= _GEN_13688;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_71 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_71 <= _GEN_3154;
        end else begin
          dirty_1_71 <= _GEN_13689;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_72 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_72 <= _GEN_3155;
        end else begin
          dirty_1_72 <= _GEN_13690;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_73 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_73 <= _GEN_3156;
        end else begin
          dirty_1_73 <= _GEN_13691;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_74 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_74 <= _GEN_3157;
        end else begin
          dirty_1_74 <= _GEN_13692;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_75 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_75 <= _GEN_3158;
        end else begin
          dirty_1_75 <= _GEN_13693;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_76 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_76 <= _GEN_3159;
        end else begin
          dirty_1_76 <= _GEN_13694;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_77 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_77 <= _GEN_3160;
        end else begin
          dirty_1_77 <= _GEN_13695;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_78 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_78 <= _GEN_3161;
        end else begin
          dirty_1_78 <= _GEN_13696;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_79 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_79 <= _GEN_3162;
        end else begin
          dirty_1_79 <= _GEN_13697;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_80 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_80 <= _GEN_3163;
        end else begin
          dirty_1_80 <= _GEN_13698;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_81 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_81 <= _GEN_3164;
        end else begin
          dirty_1_81 <= _GEN_13699;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_82 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_82 <= _GEN_3165;
        end else begin
          dirty_1_82 <= _GEN_13700;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_83 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_83 <= _GEN_3166;
        end else begin
          dirty_1_83 <= _GEN_13701;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_84 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_84 <= _GEN_3167;
        end else begin
          dirty_1_84 <= _GEN_13702;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_85 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_85 <= _GEN_3168;
        end else begin
          dirty_1_85 <= _GEN_13703;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_86 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_86 <= _GEN_3169;
        end else begin
          dirty_1_86 <= _GEN_13704;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_87 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_87 <= _GEN_3170;
        end else begin
          dirty_1_87 <= _GEN_13705;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_88 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_88 <= _GEN_3171;
        end else begin
          dirty_1_88 <= _GEN_13706;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_89 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_89 <= _GEN_3172;
        end else begin
          dirty_1_89 <= _GEN_13707;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_90 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_90 <= _GEN_3173;
        end else begin
          dirty_1_90 <= _GEN_13708;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_91 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_91 <= _GEN_3174;
        end else begin
          dirty_1_91 <= _GEN_13709;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_92 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_92 <= _GEN_3175;
        end else begin
          dirty_1_92 <= _GEN_13710;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_93 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_93 <= _GEN_3176;
        end else begin
          dirty_1_93 <= _GEN_13711;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_94 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_94 <= _GEN_3177;
        end else begin
          dirty_1_94 <= _GEN_13712;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_95 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_95 <= _GEN_3178;
        end else begin
          dirty_1_95 <= _GEN_13713;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_96 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_96 <= _GEN_3179;
        end else begin
          dirty_1_96 <= _GEN_13714;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_97 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_97 <= _GEN_3180;
        end else begin
          dirty_1_97 <= _GEN_13715;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_98 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_98 <= _GEN_3181;
        end else begin
          dirty_1_98 <= _GEN_13716;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_99 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_99 <= _GEN_3182;
        end else begin
          dirty_1_99 <= _GEN_13717;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_100 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_100 <= _GEN_3183;
        end else begin
          dirty_1_100 <= _GEN_13718;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_101 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_101 <= _GEN_3184;
        end else begin
          dirty_1_101 <= _GEN_13719;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_102 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_102 <= _GEN_3185;
        end else begin
          dirty_1_102 <= _GEN_13720;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_103 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_103 <= _GEN_3186;
        end else begin
          dirty_1_103 <= _GEN_13721;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_104 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_104 <= _GEN_3187;
        end else begin
          dirty_1_104 <= _GEN_13722;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_105 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_105 <= _GEN_3188;
        end else begin
          dirty_1_105 <= _GEN_13723;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_106 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_106 <= _GEN_3189;
        end else begin
          dirty_1_106 <= _GEN_13724;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_107 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_107 <= _GEN_3190;
        end else begin
          dirty_1_107 <= _GEN_13725;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_108 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_108 <= _GEN_3191;
        end else begin
          dirty_1_108 <= _GEN_13726;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_109 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_109 <= _GEN_3192;
        end else begin
          dirty_1_109 <= _GEN_13727;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_110 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_110 <= _GEN_3193;
        end else begin
          dirty_1_110 <= _GEN_13728;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_111 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_111 <= _GEN_3194;
        end else begin
          dirty_1_111 <= _GEN_13729;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_112 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_112 <= _GEN_3195;
        end else begin
          dirty_1_112 <= _GEN_13730;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_113 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_113 <= _GEN_3196;
        end else begin
          dirty_1_113 <= _GEN_13731;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_114 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_114 <= _GEN_3197;
        end else begin
          dirty_1_114 <= _GEN_13732;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_115 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_115 <= _GEN_3198;
        end else begin
          dirty_1_115 <= _GEN_13733;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_116 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_116 <= _GEN_3199;
        end else begin
          dirty_1_116 <= _GEN_13734;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_117 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_117 <= _GEN_3200;
        end else begin
          dirty_1_117 <= _GEN_13735;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_118 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_118 <= _GEN_3201;
        end else begin
          dirty_1_118 <= _GEN_13736;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_119 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_119 <= _GEN_3202;
        end else begin
          dirty_1_119 <= _GEN_13737;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_120 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_120 <= _GEN_3203;
        end else begin
          dirty_1_120 <= _GEN_13738;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_121 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_121 <= _GEN_3204;
        end else begin
          dirty_1_121 <= _GEN_13739;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_122 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_122 <= _GEN_3205;
        end else begin
          dirty_1_122 <= _GEN_13740;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_123 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_123 <= _GEN_3206;
        end else begin
          dirty_1_123 <= _GEN_13741;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_124 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_124 <= _GEN_3207;
        end else begin
          dirty_1_124 <= _GEN_13742;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_125 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_125 <= _GEN_3208;
        end else begin
          dirty_1_125 <= _GEN_13743;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_126 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_126 <= _GEN_3209;
        end else begin
          dirty_1_126 <= _GEN_13744;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_127 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_127 <= _GEN_3210;
        end else begin
          dirty_1_127 <= _GEN_13745;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:27]
      way0_hit <= 1'h0; // @[d_cache.scala 28:27]
    end else begin
      way0_hit <= _T_6;
    end
    if (reset) begin // @[d_cache.scala 29:27]
      way1_hit <= 1'h0; // @[d_cache.scala 29:27]
    end else begin
      way1_hit <= _T_11;
    end
    if (reset) begin // @[d_cache.scala 31:34]
      write_back_data <= 64'h0; // @[d_cache.scala 31:34]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          write_back_data <= _GEN_13488;
        end
      end
    end
    write_back_addr <= _GEN_19500[31:0]; // @[d_cache.scala 32:{34,34}]
    if (reset) begin // @[d_cache.scala 35:28]
      unuse_way <= 2'h0; // @[d_cache.scala 35:28]
    end else if (~_GEN_255) begin // @[d_cache.scala 68:31]
      unuse_way <= 2'h1; // @[d_cache.scala 69:19]
    end else if (~_GEN_512) begin // @[d_cache.scala 70:37]
      unuse_way <= 2'h2; // @[d_cache.scala 71:19]
    end else begin
      unuse_way <= 2'h0; // @[d_cache.scala 73:19]
    end
    if (reset) begin // @[d_cache.scala 36:31]
      receive_data <= 64'h0; // @[d_cache.scala 36:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          receive_data <= _GEN_12718;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:24]
      quene <= 1'h0; // @[d_cache.scala 37:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          quene <= _GEN_13103;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 76:24]
      state <= 3'h0; // @[d_cache.scala 76:24]
    end else if (3'h0 == state) begin // @[d_cache.scala 81:18]
      if (io_from_lsu_arvalid) begin // @[d_cache.scala 83:38]
        state <= 3'h1; // @[d_cache.scala 84:23]
      end else if (io_from_lsu_awvalid) begin // @[d_cache.scala 85:44]
        state <= 3'h2; // @[d_cache.scala 86:23]
      end
    end else if (3'h1 == state) begin // @[d_cache.scala 81:18]
      if (way0_hit) begin // @[d_cache.scala 91:27]
        state <= _GEN_902;
      end else begin
        state <= _GEN_1031;
      end
    end else if (3'h2 == state) begin // @[d_cache.scala 81:18]
      state <= _GEN_2442;
    end else begin
      state <= _GEN_12717;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"read addr : %x  write addr : %x\n",io_from_lsu_araddr,io_from_lsu_awaddr); // @[d_cache.scala 15:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"d_cache state:%d\n",state); // @[d_cache.scala 77:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"receive data:%x\n",receive_data); // @[d_cache.scala 79:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_20 & _T_21 & way0_hit & io_from_lsu_rready & _T_1) begin
          $fwrite(32'h80000002,"dirty_0:%d\n",7'h7f == index[6:0] ? dirty_0_127 : _GEN_900); // @[d_cache.scala 93:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19502 & ~way0_hit & way1_hit & io_from_lsu_rready & _T_1) begin
          $fwrite(32'h80000002,"dirty_1:%d\n",7'h7f == index[6:0] ? dirty_1_127 : _GEN_1029); // @[d_cache.scala 99:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"cacheline0:%x   cacheline1:%x\n",_GEN_1160,_GEN_1672); // @[d_cache.scala 362:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"recent_wdata0:%x  recent_wdata1:%x\n",7'h7f == index[6:0] ? recent_wdata0_127 :
            _GEN_18335,7'h7f == index[6:0] ? recent_wdata1_127 : _GEN_18463); // @[d_cache.scala 363:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ram_0_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ram_0_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ram_0_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ram_0_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ram_0_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ram_0_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ram_0_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ram_0_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  ram_0_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  ram_0_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  ram_0_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  ram_0_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  ram_0_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  ram_0_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  ram_0_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  ram_0_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  ram_0_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  ram_0_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  ram_0_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  ram_0_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  ram_0_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  ram_0_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  ram_0_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  ram_0_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  ram_0_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  ram_0_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  ram_0_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  ram_0_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  ram_0_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  ram_0_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  ram_0_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  ram_0_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  ram_0_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  ram_0_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  ram_0_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  ram_0_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  ram_0_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  ram_0_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  ram_0_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  ram_0_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  ram_0_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  ram_0_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  ram_0_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  ram_0_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  ram_0_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  ram_0_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  ram_0_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  ram_0_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  ram_0_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  ram_0_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  ram_0_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  ram_0_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  ram_0_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  ram_0_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  ram_0_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  ram_0_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  ram_0_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  ram_0_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  ram_0_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  ram_0_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  ram_0_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  ram_0_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  ram_0_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  ram_0_63 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  ram_0_64 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  ram_0_65 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  ram_0_66 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  ram_0_67 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  ram_0_68 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  ram_0_69 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  ram_0_70 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  ram_0_71 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  ram_0_72 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  ram_0_73 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  ram_0_74 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  ram_0_75 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  ram_0_76 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  ram_0_77 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  ram_0_78 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  ram_0_79 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  ram_0_80 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  ram_0_81 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  ram_0_82 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  ram_0_83 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  ram_0_84 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  ram_0_85 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  ram_0_86 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  ram_0_87 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  ram_0_88 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  ram_0_89 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  ram_0_90 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  ram_0_91 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  ram_0_92 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  ram_0_93 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  ram_0_94 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  ram_0_95 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  ram_0_96 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  ram_0_97 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  ram_0_98 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  ram_0_99 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  ram_0_100 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  ram_0_101 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  ram_0_102 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  ram_0_103 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  ram_0_104 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  ram_0_105 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  ram_0_106 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  ram_0_107 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  ram_0_108 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  ram_0_109 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  ram_0_110 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  ram_0_111 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  ram_0_112 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  ram_0_113 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  ram_0_114 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  ram_0_115 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  ram_0_116 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  ram_0_117 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  ram_0_118 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  ram_0_119 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  ram_0_120 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  ram_0_121 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  ram_0_122 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  ram_0_123 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  ram_0_124 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  ram_0_125 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  ram_0_126 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  ram_0_127 = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  ram_1_0 = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  ram_1_1 = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  ram_1_2 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  ram_1_3 = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  ram_1_4 = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  ram_1_5 = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  ram_1_6 = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  ram_1_7 = _RAND_135[63:0];
  _RAND_136 = {2{`RANDOM}};
  ram_1_8 = _RAND_136[63:0];
  _RAND_137 = {2{`RANDOM}};
  ram_1_9 = _RAND_137[63:0];
  _RAND_138 = {2{`RANDOM}};
  ram_1_10 = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  ram_1_11 = _RAND_139[63:0];
  _RAND_140 = {2{`RANDOM}};
  ram_1_12 = _RAND_140[63:0];
  _RAND_141 = {2{`RANDOM}};
  ram_1_13 = _RAND_141[63:0];
  _RAND_142 = {2{`RANDOM}};
  ram_1_14 = _RAND_142[63:0];
  _RAND_143 = {2{`RANDOM}};
  ram_1_15 = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  ram_1_16 = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  ram_1_17 = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  ram_1_18 = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  ram_1_19 = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  ram_1_20 = _RAND_148[63:0];
  _RAND_149 = {2{`RANDOM}};
  ram_1_21 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  ram_1_22 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  ram_1_23 = _RAND_151[63:0];
  _RAND_152 = {2{`RANDOM}};
  ram_1_24 = _RAND_152[63:0];
  _RAND_153 = {2{`RANDOM}};
  ram_1_25 = _RAND_153[63:0];
  _RAND_154 = {2{`RANDOM}};
  ram_1_26 = _RAND_154[63:0];
  _RAND_155 = {2{`RANDOM}};
  ram_1_27 = _RAND_155[63:0];
  _RAND_156 = {2{`RANDOM}};
  ram_1_28 = _RAND_156[63:0];
  _RAND_157 = {2{`RANDOM}};
  ram_1_29 = _RAND_157[63:0];
  _RAND_158 = {2{`RANDOM}};
  ram_1_30 = _RAND_158[63:0];
  _RAND_159 = {2{`RANDOM}};
  ram_1_31 = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  ram_1_32 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  ram_1_33 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  ram_1_34 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  ram_1_35 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  ram_1_36 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  ram_1_37 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  ram_1_38 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  ram_1_39 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  ram_1_40 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  ram_1_41 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  ram_1_42 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  ram_1_43 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  ram_1_44 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  ram_1_45 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  ram_1_46 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  ram_1_47 = _RAND_175[63:0];
  _RAND_176 = {2{`RANDOM}};
  ram_1_48 = _RAND_176[63:0];
  _RAND_177 = {2{`RANDOM}};
  ram_1_49 = _RAND_177[63:0];
  _RAND_178 = {2{`RANDOM}};
  ram_1_50 = _RAND_178[63:0];
  _RAND_179 = {2{`RANDOM}};
  ram_1_51 = _RAND_179[63:0];
  _RAND_180 = {2{`RANDOM}};
  ram_1_52 = _RAND_180[63:0];
  _RAND_181 = {2{`RANDOM}};
  ram_1_53 = _RAND_181[63:0];
  _RAND_182 = {2{`RANDOM}};
  ram_1_54 = _RAND_182[63:0];
  _RAND_183 = {2{`RANDOM}};
  ram_1_55 = _RAND_183[63:0];
  _RAND_184 = {2{`RANDOM}};
  ram_1_56 = _RAND_184[63:0];
  _RAND_185 = {2{`RANDOM}};
  ram_1_57 = _RAND_185[63:0];
  _RAND_186 = {2{`RANDOM}};
  ram_1_58 = _RAND_186[63:0];
  _RAND_187 = {2{`RANDOM}};
  ram_1_59 = _RAND_187[63:0];
  _RAND_188 = {2{`RANDOM}};
  ram_1_60 = _RAND_188[63:0];
  _RAND_189 = {2{`RANDOM}};
  ram_1_61 = _RAND_189[63:0];
  _RAND_190 = {2{`RANDOM}};
  ram_1_62 = _RAND_190[63:0];
  _RAND_191 = {2{`RANDOM}};
  ram_1_63 = _RAND_191[63:0];
  _RAND_192 = {2{`RANDOM}};
  ram_1_64 = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  ram_1_65 = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  ram_1_66 = _RAND_194[63:0];
  _RAND_195 = {2{`RANDOM}};
  ram_1_67 = _RAND_195[63:0];
  _RAND_196 = {2{`RANDOM}};
  ram_1_68 = _RAND_196[63:0];
  _RAND_197 = {2{`RANDOM}};
  ram_1_69 = _RAND_197[63:0];
  _RAND_198 = {2{`RANDOM}};
  ram_1_70 = _RAND_198[63:0];
  _RAND_199 = {2{`RANDOM}};
  ram_1_71 = _RAND_199[63:0];
  _RAND_200 = {2{`RANDOM}};
  ram_1_72 = _RAND_200[63:0];
  _RAND_201 = {2{`RANDOM}};
  ram_1_73 = _RAND_201[63:0];
  _RAND_202 = {2{`RANDOM}};
  ram_1_74 = _RAND_202[63:0];
  _RAND_203 = {2{`RANDOM}};
  ram_1_75 = _RAND_203[63:0];
  _RAND_204 = {2{`RANDOM}};
  ram_1_76 = _RAND_204[63:0];
  _RAND_205 = {2{`RANDOM}};
  ram_1_77 = _RAND_205[63:0];
  _RAND_206 = {2{`RANDOM}};
  ram_1_78 = _RAND_206[63:0];
  _RAND_207 = {2{`RANDOM}};
  ram_1_79 = _RAND_207[63:0];
  _RAND_208 = {2{`RANDOM}};
  ram_1_80 = _RAND_208[63:0];
  _RAND_209 = {2{`RANDOM}};
  ram_1_81 = _RAND_209[63:0];
  _RAND_210 = {2{`RANDOM}};
  ram_1_82 = _RAND_210[63:0];
  _RAND_211 = {2{`RANDOM}};
  ram_1_83 = _RAND_211[63:0];
  _RAND_212 = {2{`RANDOM}};
  ram_1_84 = _RAND_212[63:0];
  _RAND_213 = {2{`RANDOM}};
  ram_1_85 = _RAND_213[63:0];
  _RAND_214 = {2{`RANDOM}};
  ram_1_86 = _RAND_214[63:0];
  _RAND_215 = {2{`RANDOM}};
  ram_1_87 = _RAND_215[63:0];
  _RAND_216 = {2{`RANDOM}};
  ram_1_88 = _RAND_216[63:0];
  _RAND_217 = {2{`RANDOM}};
  ram_1_89 = _RAND_217[63:0];
  _RAND_218 = {2{`RANDOM}};
  ram_1_90 = _RAND_218[63:0];
  _RAND_219 = {2{`RANDOM}};
  ram_1_91 = _RAND_219[63:0];
  _RAND_220 = {2{`RANDOM}};
  ram_1_92 = _RAND_220[63:0];
  _RAND_221 = {2{`RANDOM}};
  ram_1_93 = _RAND_221[63:0];
  _RAND_222 = {2{`RANDOM}};
  ram_1_94 = _RAND_222[63:0];
  _RAND_223 = {2{`RANDOM}};
  ram_1_95 = _RAND_223[63:0];
  _RAND_224 = {2{`RANDOM}};
  ram_1_96 = _RAND_224[63:0];
  _RAND_225 = {2{`RANDOM}};
  ram_1_97 = _RAND_225[63:0];
  _RAND_226 = {2{`RANDOM}};
  ram_1_98 = _RAND_226[63:0];
  _RAND_227 = {2{`RANDOM}};
  ram_1_99 = _RAND_227[63:0];
  _RAND_228 = {2{`RANDOM}};
  ram_1_100 = _RAND_228[63:0];
  _RAND_229 = {2{`RANDOM}};
  ram_1_101 = _RAND_229[63:0];
  _RAND_230 = {2{`RANDOM}};
  ram_1_102 = _RAND_230[63:0];
  _RAND_231 = {2{`RANDOM}};
  ram_1_103 = _RAND_231[63:0];
  _RAND_232 = {2{`RANDOM}};
  ram_1_104 = _RAND_232[63:0];
  _RAND_233 = {2{`RANDOM}};
  ram_1_105 = _RAND_233[63:0];
  _RAND_234 = {2{`RANDOM}};
  ram_1_106 = _RAND_234[63:0];
  _RAND_235 = {2{`RANDOM}};
  ram_1_107 = _RAND_235[63:0];
  _RAND_236 = {2{`RANDOM}};
  ram_1_108 = _RAND_236[63:0];
  _RAND_237 = {2{`RANDOM}};
  ram_1_109 = _RAND_237[63:0];
  _RAND_238 = {2{`RANDOM}};
  ram_1_110 = _RAND_238[63:0];
  _RAND_239 = {2{`RANDOM}};
  ram_1_111 = _RAND_239[63:0];
  _RAND_240 = {2{`RANDOM}};
  ram_1_112 = _RAND_240[63:0];
  _RAND_241 = {2{`RANDOM}};
  ram_1_113 = _RAND_241[63:0];
  _RAND_242 = {2{`RANDOM}};
  ram_1_114 = _RAND_242[63:0];
  _RAND_243 = {2{`RANDOM}};
  ram_1_115 = _RAND_243[63:0];
  _RAND_244 = {2{`RANDOM}};
  ram_1_116 = _RAND_244[63:0];
  _RAND_245 = {2{`RANDOM}};
  ram_1_117 = _RAND_245[63:0];
  _RAND_246 = {2{`RANDOM}};
  ram_1_118 = _RAND_246[63:0];
  _RAND_247 = {2{`RANDOM}};
  ram_1_119 = _RAND_247[63:0];
  _RAND_248 = {2{`RANDOM}};
  ram_1_120 = _RAND_248[63:0];
  _RAND_249 = {2{`RANDOM}};
  ram_1_121 = _RAND_249[63:0];
  _RAND_250 = {2{`RANDOM}};
  ram_1_122 = _RAND_250[63:0];
  _RAND_251 = {2{`RANDOM}};
  ram_1_123 = _RAND_251[63:0];
  _RAND_252 = {2{`RANDOM}};
  ram_1_124 = _RAND_252[63:0];
  _RAND_253 = {2{`RANDOM}};
  ram_1_125 = _RAND_253[63:0];
  _RAND_254 = {2{`RANDOM}};
  ram_1_126 = _RAND_254[63:0];
  _RAND_255 = {2{`RANDOM}};
  ram_1_127 = _RAND_255[63:0];
  _RAND_256 = {2{`RANDOM}};
  recent_wdata0_0 = _RAND_256[63:0];
  _RAND_257 = {2{`RANDOM}};
  recent_wdata0_1 = _RAND_257[63:0];
  _RAND_258 = {2{`RANDOM}};
  recent_wdata0_2 = _RAND_258[63:0];
  _RAND_259 = {2{`RANDOM}};
  recent_wdata0_3 = _RAND_259[63:0];
  _RAND_260 = {2{`RANDOM}};
  recent_wdata0_4 = _RAND_260[63:0];
  _RAND_261 = {2{`RANDOM}};
  recent_wdata0_5 = _RAND_261[63:0];
  _RAND_262 = {2{`RANDOM}};
  recent_wdata0_6 = _RAND_262[63:0];
  _RAND_263 = {2{`RANDOM}};
  recent_wdata0_7 = _RAND_263[63:0];
  _RAND_264 = {2{`RANDOM}};
  recent_wdata0_8 = _RAND_264[63:0];
  _RAND_265 = {2{`RANDOM}};
  recent_wdata0_9 = _RAND_265[63:0];
  _RAND_266 = {2{`RANDOM}};
  recent_wdata0_10 = _RAND_266[63:0];
  _RAND_267 = {2{`RANDOM}};
  recent_wdata0_11 = _RAND_267[63:0];
  _RAND_268 = {2{`RANDOM}};
  recent_wdata0_12 = _RAND_268[63:0];
  _RAND_269 = {2{`RANDOM}};
  recent_wdata0_13 = _RAND_269[63:0];
  _RAND_270 = {2{`RANDOM}};
  recent_wdata0_14 = _RAND_270[63:0];
  _RAND_271 = {2{`RANDOM}};
  recent_wdata0_15 = _RAND_271[63:0];
  _RAND_272 = {2{`RANDOM}};
  recent_wdata0_16 = _RAND_272[63:0];
  _RAND_273 = {2{`RANDOM}};
  recent_wdata0_17 = _RAND_273[63:0];
  _RAND_274 = {2{`RANDOM}};
  recent_wdata0_18 = _RAND_274[63:0];
  _RAND_275 = {2{`RANDOM}};
  recent_wdata0_19 = _RAND_275[63:0];
  _RAND_276 = {2{`RANDOM}};
  recent_wdata0_20 = _RAND_276[63:0];
  _RAND_277 = {2{`RANDOM}};
  recent_wdata0_21 = _RAND_277[63:0];
  _RAND_278 = {2{`RANDOM}};
  recent_wdata0_22 = _RAND_278[63:0];
  _RAND_279 = {2{`RANDOM}};
  recent_wdata0_23 = _RAND_279[63:0];
  _RAND_280 = {2{`RANDOM}};
  recent_wdata0_24 = _RAND_280[63:0];
  _RAND_281 = {2{`RANDOM}};
  recent_wdata0_25 = _RAND_281[63:0];
  _RAND_282 = {2{`RANDOM}};
  recent_wdata0_26 = _RAND_282[63:0];
  _RAND_283 = {2{`RANDOM}};
  recent_wdata0_27 = _RAND_283[63:0];
  _RAND_284 = {2{`RANDOM}};
  recent_wdata0_28 = _RAND_284[63:0];
  _RAND_285 = {2{`RANDOM}};
  recent_wdata0_29 = _RAND_285[63:0];
  _RAND_286 = {2{`RANDOM}};
  recent_wdata0_30 = _RAND_286[63:0];
  _RAND_287 = {2{`RANDOM}};
  recent_wdata0_31 = _RAND_287[63:0];
  _RAND_288 = {2{`RANDOM}};
  recent_wdata0_32 = _RAND_288[63:0];
  _RAND_289 = {2{`RANDOM}};
  recent_wdata0_33 = _RAND_289[63:0];
  _RAND_290 = {2{`RANDOM}};
  recent_wdata0_34 = _RAND_290[63:0];
  _RAND_291 = {2{`RANDOM}};
  recent_wdata0_35 = _RAND_291[63:0];
  _RAND_292 = {2{`RANDOM}};
  recent_wdata0_36 = _RAND_292[63:0];
  _RAND_293 = {2{`RANDOM}};
  recent_wdata0_37 = _RAND_293[63:0];
  _RAND_294 = {2{`RANDOM}};
  recent_wdata0_38 = _RAND_294[63:0];
  _RAND_295 = {2{`RANDOM}};
  recent_wdata0_39 = _RAND_295[63:0];
  _RAND_296 = {2{`RANDOM}};
  recent_wdata0_40 = _RAND_296[63:0];
  _RAND_297 = {2{`RANDOM}};
  recent_wdata0_41 = _RAND_297[63:0];
  _RAND_298 = {2{`RANDOM}};
  recent_wdata0_42 = _RAND_298[63:0];
  _RAND_299 = {2{`RANDOM}};
  recent_wdata0_43 = _RAND_299[63:0];
  _RAND_300 = {2{`RANDOM}};
  recent_wdata0_44 = _RAND_300[63:0];
  _RAND_301 = {2{`RANDOM}};
  recent_wdata0_45 = _RAND_301[63:0];
  _RAND_302 = {2{`RANDOM}};
  recent_wdata0_46 = _RAND_302[63:0];
  _RAND_303 = {2{`RANDOM}};
  recent_wdata0_47 = _RAND_303[63:0];
  _RAND_304 = {2{`RANDOM}};
  recent_wdata0_48 = _RAND_304[63:0];
  _RAND_305 = {2{`RANDOM}};
  recent_wdata0_49 = _RAND_305[63:0];
  _RAND_306 = {2{`RANDOM}};
  recent_wdata0_50 = _RAND_306[63:0];
  _RAND_307 = {2{`RANDOM}};
  recent_wdata0_51 = _RAND_307[63:0];
  _RAND_308 = {2{`RANDOM}};
  recent_wdata0_52 = _RAND_308[63:0];
  _RAND_309 = {2{`RANDOM}};
  recent_wdata0_53 = _RAND_309[63:0];
  _RAND_310 = {2{`RANDOM}};
  recent_wdata0_54 = _RAND_310[63:0];
  _RAND_311 = {2{`RANDOM}};
  recent_wdata0_55 = _RAND_311[63:0];
  _RAND_312 = {2{`RANDOM}};
  recent_wdata0_56 = _RAND_312[63:0];
  _RAND_313 = {2{`RANDOM}};
  recent_wdata0_57 = _RAND_313[63:0];
  _RAND_314 = {2{`RANDOM}};
  recent_wdata0_58 = _RAND_314[63:0];
  _RAND_315 = {2{`RANDOM}};
  recent_wdata0_59 = _RAND_315[63:0];
  _RAND_316 = {2{`RANDOM}};
  recent_wdata0_60 = _RAND_316[63:0];
  _RAND_317 = {2{`RANDOM}};
  recent_wdata0_61 = _RAND_317[63:0];
  _RAND_318 = {2{`RANDOM}};
  recent_wdata0_62 = _RAND_318[63:0];
  _RAND_319 = {2{`RANDOM}};
  recent_wdata0_63 = _RAND_319[63:0];
  _RAND_320 = {2{`RANDOM}};
  recent_wdata0_64 = _RAND_320[63:0];
  _RAND_321 = {2{`RANDOM}};
  recent_wdata0_65 = _RAND_321[63:0];
  _RAND_322 = {2{`RANDOM}};
  recent_wdata0_66 = _RAND_322[63:0];
  _RAND_323 = {2{`RANDOM}};
  recent_wdata0_67 = _RAND_323[63:0];
  _RAND_324 = {2{`RANDOM}};
  recent_wdata0_68 = _RAND_324[63:0];
  _RAND_325 = {2{`RANDOM}};
  recent_wdata0_69 = _RAND_325[63:0];
  _RAND_326 = {2{`RANDOM}};
  recent_wdata0_70 = _RAND_326[63:0];
  _RAND_327 = {2{`RANDOM}};
  recent_wdata0_71 = _RAND_327[63:0];
  _RAND_328 = {2{`RANDOM}};
  recent_wdata0_72 = _RAND_328[63:0];
  _RAND_329 = {2{`RANDOM}};
  recent_wdata0_73 = _RAND_329[63:0];
  _RAND_330 = {2{`RANDOM}};
  recent_wdata0_74 = _RAND_330[63:0];
  _RAND_331 = {2{`RANDOM}};
  recent_wdata0_75 = _RAND_331[63:0];
  _RAND_332 = {2{`RANDOM}};
  recent_wdata0_76 = _RAND_332[63:0];
  _RAND_333 = {2{`RANDOM}};
  recent_wdata0_77 = _RAND_333[63:0];
  _RAND_334 = {2{`RANDOM}};
  recent_wdata0_78 = _RAND_334[63:0];
  _RAND_335 = {2{`RANDOM}};
  recent_wdata0_79 = _RAND_335[63:0];
  _RAND_336 = {2{`RANDOM}};
  recent_wdata0_80 = _RAND_336[63:0];
  _RAND_337 = {2{`RANDOM}};
  recent_wdata0_81 = _RAND_337[63:0];
  _RAND_338 = {2{`RANDOM}};
  recent_wdata0_82 = _RAND_338[63:0];
  _RAND_339 = {2{`RANDOM}};
  recent_wdata0_83 = _RAND_339[63:0];
  _RAND_340 = {2{`RANDOM}};
  recent_wdata0_84 = _RAND_340[63:0];
  _RAND_341 = {2{`RANDOM}};
  recent_wdata0_85 = _RAND_341[63:0];
  _RAND_342 = {2{`RANDOM}};
  recent_wdata0_86 = _RAND_342[63:0];
  _RAND_343 = {2{`RANDOM}};
  recent_wdata0_87 = _RAND_343[63:0];
  _RAND_344 = {2{`RANDOM}};
  recent_wdata0_88 = _RAND_344[63:0];
  _RAND_345 = {2{`RANDOM}};
  recent_wdata0_89 = _RAND_345[63:0];
  _RAND_346 = {2{`RANDOM}};
  recent_wdata0_90 = _RAND_346[63:0];
  _RAND_347 = {2{`RANDOM}};
  recent_wdata0_91 = _RAND_347[63:0];
  _RAND_348 = {2{`RANDOM}};
  recent_wdata0_92 = _RAND_348[63:0];
  _RAND_349 = {2{`RANDOM}};
  recent_wdata0_93 = _RAND_349[63:0];
  _RAND_350 = {2{`RANDOM}};
  recent_wdata0_94 = _RAND_350[63:0];
  _RAND_351 = {2{`RANDOM}};
  recent_wdata0_95 = _RAND_351[63:0];
  _RAND_352 = {2{`RANDOM}};
  recent_wdata0_96 = _RAND_352[63:0];
  _RAND_353 = {2{`RANDOM}};
  recent_wdata0_97 = _RAND_353[63:0];
  _RAND_354 = {2{`RANDOM}};
  recent_wdata0_98 = _RAND_354[63:0];
  _RAND_355 = {2{`RANDOM}};
  recent_wdata0_99 = _RAND_355[63:0];
  _RAND_356 = {2{`RANDOM}};
  recent_wdata0_100 = _RAND_356[63:0];
  _RAND_357 = {2{`RANDOM}};
  recent_wdata0_101 = _RAND_357[63:0];
  _RAND_358 = {2{`RANDOM}};
  recent_wdata0_102 = _RAND_358[63:0];
  _RAND_359 = {2{`RANDOM}};
  recent_wdata0_103 = _RAND_359[63:0];
  _RAND_360 = {2{`RANDOM}};
  recent_wdata0_104 = _RAND_360[63:0];
  _RAND_361 = {2{`RANDOM}};
  recent_wdata0_105 = _RAND_361[63:0];
  _RAND_362 = {2{`RANDOM}};
  recent_wdata0_106 = _RAND_362[63:0];
  _RAND_363 = {2{`RANDOM}};
  recent_wdata0_107 = _RAND_363[63:0];
  _RAND_364 = {2{`RANDOM}};
  recent_wdata0_108 = _RAND_364[63:0];
  _RAND_365 = {2{`RANDOM}};
  recent_wdata0_109 = _RAND_365[63:0];
  _RAND_366 = {2{`RANDOM}};
  recent_wdata0_110 = _RAND_366[63:0];
  _RAND_367 = {2{`RANDOM}};
  recent_wdata0_111 = _RAND_367[63:0];
  _RAND_368 = {2{`RANDOM}};
  recent_wdata0_112 = _RAND_368[63:0];
  _RAND_369 = {2{`RANDOM}};
  recent_wdata0_113 = _RAND_369[63:0];
  _RAND_370 = {2{`RANDOM}};
  recent_wdata0_114 = _RAND_370[63:0];
  _RAND_371 = {2{`RANDOM}};
  recent_wdata0_115 = _RAND_371[63:0];
  _RAND_372 = {2{`RANDOM}};
  recent_wdata0_116 = _RAND_372[63:0];
  _RAND_373 = {2{`RANDOM}};
  recent_wdata0_117 = _RAND_373[63:0];
  _RAND_374 = {2{`RANDOM}};
  recent_wdata0_118 = _RAND_374[63:0];
  _RAND_375 = {2{`RANDOM}};
  recent_wdata0_119 = _RAND_375[63:0];
  _RAND_376 = {2{`RANDOM}};
  recent_wdata0_120 = _RAND_376[63:0];
  _RAND_377 = {2{`RANDOM}};
  recent_wdata0_121 = _RAND_377[63:0];
  _RAND_378 = {2{`RANDOM}};
  recent_wdata0_122 = _RAND_378[63:0];
  _RAND_379 = {2{`RANDOM}};
  recent_wdata0_123 = _RAND_379[63:0];
  _RAND_380 = {2{`RANDOM}};
  recent_wdata0_124 = _RAND_380[63:0];
  _RAND_381 = {2{`RANDOM}};
  recent_wdata0_125 = _RAND_381[63:0];
  _RAND_382 = {2{`RANDOM}};
  recent_wdata0_126 = _RAND_382[63:0];
  _RAND_383 = {2{`RANDOM}};
  recent_wdata0_127 = _RAND_383[63:0];
  _RAND_384 = {2{`RANDOM}};
  recent_wdata1_0 = _RAND_384[63:0];
  _RAND_385 = {2{`RANDOM}};
  recent_wdata1_1 = _RAND_385[63:0];
  _RAND_386 = {2{`RANDOM}};
  recent_wdata1_2 = _RAND_386[63:0];
  _RAND_387 = {2{`RANDOM}};
  recent_wdata1_3 = _RAND_387[63:0];
  _RAND_388 = {2{`RANDOM}};
  recent_wdata1_4 = _RAND_388[63:0];
  _RAND_389 = {2{`RANDOM}};
  recent_wdata1_5 = _RAND_389[63:0];
  _RAND_390 = {2{`RANDOM}};
  recent_wdata1_6 = _RAND_390[63:0];
  _RAND_391 = {2{`RANDOM}};
  recent_wdata1_7 = _RAND_391[63:0];
  _RAND_392 = {2{`RANDOM}};
  recent_wdata1_8 = _RAND_392[63:0];
  _RAND_393 = {2{`RANDOM}};
  recent_wdata1_9 = _RAND_393[63:0];
  _RAND_394 = {2{`RANDOM}};
  recent_wdata1_10 = _RAND_394[63:0];
  _RAND_395 = {2{`RANDOM}};
  recent_wdata1_11 = _RAND_395[63:0];
  _RAND_396 = {2{`RANDOM}};
  recent_wdata1_12 = _RAND_396[63:0];
  _RAND_397 = {2{`RANDOM}};
  recent_wdata1_13 = _RAND_397[63:0];
  _RAND_398 = {2{`RANDOM}};
  recent_wdata1_14 = _RAND_398[63:0];
  _RAND_399 = {2{`RANDOM}};
  recent_wdata1_15 = _RAND_399[63:0];
  _RAND_400 = {2{`RANDOM}};
  recent_wdata1_16 = _RAND_400[63:0];
  _RAND_401 = {2{`RANDOM}};
  recent_wdata1_17 = _RAND_401[63:0];
  _RAND_402 = {2{`RANDOM}};
  recent_wdata1_18 = _RAND_402[63:0];
  _RAND_403 = {2{`RANDOM}};
  recent_wdata1_19 = _RAND_403[63:0];
  _RAND_404 = {2{`RANDOM}};
  recent_wdata1_20 = _RAND_404[63:0];
  _RAND_405 = {2{`RANDOM}};
  recent_wdata1_21 = _RAND_405[63:0];
  _RAND_406 = {2{`RANDOM}};
  recent_wdata1_22 = _RAND_406[63:0];
  _RAND_407 = {2{`RANDOM}};
  recent_wdata1_23 = _RAND_407[63:0];
  _RAND_408 = {2{`RANDOM}};
  recent_wdata1_24 = _RAND_408[63:0];
  _RAND_409 = {2{`RANDOM}};
  recent_wdata1_25 = _RAND_409[63:0];
  _RAND_410 = {2{`RANDOM}};
  recent_wdata1_26 = _RAND_410[63:0];
  _RAND_411 = {2{`RANDOM}};
  recent_wdata1_27 = _RAND_411[63:0];
  _RAND_412 = {2{`RANDOM}};
  recent_wdata1_28 = _RAND_412[63:0];
  _RAND_413 = {2{`RANDOM}};
  recent_wdata1_29 = _RAND_413[63:0];
  _RAND_414 = {2{`RANDOM}};
  recent_wdata1_30 = _RAND_414[63:0];
  _RAND_415 = {2{`RANDOM}};
  recent_wdata1_31 = _RAND_415[63:0];
  _RAND_416 = {2{`RANDOM}};
  recent_wdata1_32 = _RAND_416[63:0];
  _RAND_417 = {2{`RANDOM}};
  recent_wdata1_33 = _RAND_417[63:0];
  _RAND_418 = {2{`RANDOM}};
  recent_wdata1_34 = _RAND_418[63:0];
  _RAND_419 = {2{`RANDOM}};
  recent_wdata1_35 = _RAND_419[63:0];
  _RAND_420 = {2{`RANDOM}};
  recent_wdata1_36 = _RAND_420[63:0];
  _RAND_421 = {2{`RANDOM}};
  recent_wdata1_37 = _RAND_421[63:0];
  _RAND_422 = {2{`RANDOM}};
  recent_wdata1_38 = _RAND_422[63:0];
  _RAND_423 = {2{`RANDOM}};
  recent_wdata1_39 = _RAND_423[63:0];
  _RAND_424 = {2{`RANDOM}};
  recent_wdata1_40 = _RAND_424[63:0];
  _RAND_425 = {2{`RANDOM}};
  recent_wdata1_41 = _RAND_425[63:0];
  _RAND_426 = {2{`RANDOM}};
  recent_wdata1_42 = _RAND_426[63:0];
  _RAND_427 = {2{`RANDOM}};
  recent_wdata1_43 = _RAND_427[63:0];
  _RAND_428 = {2{`RANDOM}};
  recent_wdata1_44 = _RAND_428[63:0];
  _RAND_429 = {2{`RANDOM}};
  recent_wdata1_45 = _RAND_429[63:0];
  _RAND_430 = {2{`RANDOM}};
  recent_wdata1_46 = _RAND_430[63:0];
  _RAND_431 = {2{`RANDOM}};
  recent_wdata1_47 = _RAND_431[63:0];
  _RAND_432 = {2{`RANDOM}};
  recent_wdata1_48 = _RAND_432[63:0];
  _RAND_433 = {2{`RANDOM}};
  recent_wdata1_49 = _RAND_433[63:0];
  _RAND_434 = {2{`RANDOM}};
  recent_wdata1_50 = _RAND_434[63:0];
  _RAND_435 = {2{`RANDOM}};
  recent_wdata1_51 = _RAND_435[63:0];
  _RAND_436 = {2{`RANDOM}};
  recent_wdata1_52 = _RAND_436[63:0];
  _RAND_437 = {2{`RANDOM}};
  recent_wdata1_53 = _RAND_437[63:0];
  _RAND_438 = {2{`RANDOM}};
  recent_wdata1_54 = _RAND_438[63:0];
  _RAND_439 = {2{`RANDOM}};
  recent_wdata1_55 = _RAND_439[63:0];
  _RAND_440 = {2{`RANDOM}};
  recent_wdata1_56 = _RAND_440[63:0];
  _RAND_441 = {2{`RANDOM}};
  recent_wdata1_57 = _RAND_441[63:0];
  _RAND_442 = {2{`RANDOM}};
  recent_wdata1_58 = _RAND_442[63:0];
  _RAND_443 = {2{`RANDOM}};
  recent_wdata1_59 = _RAND_443[63:0];
  _RAND_444 = {2{`RANDOM}};
  recent_wdata1_60 = _RAND_444[63:0];
  _RAND_445 = {2{`RANDOM}};
  recent_wdata1_61 = _RAND_445[63:0];
  _RAND_446 = {2{`RANDOM}};
  recent_wdata1_62 = _RAND_446[63:0];
  _RAND_447 = {2{`RANDOM}};
  recent_wdata1_63 = _RAND_447[63:0];
  _RAND_448 = {2{`RANDOM}};
  recent_wdata1_64 = _RAND_448[63:0];
  _RAND_449 = {2{`RANDOM}};
  recent_wdata1_65 = _RAND_449[63:0];
  _RAND_450 = {2{`RANDOM}};
  recent_wdata1_66 = _RAND_450[63:0];
  _RAND_451 = {2{`RANDOM}};
  recent_wdata1_67 = _RAND_451[63:0];
  _RAND_452 = {2{`RANDOM}};
  recent_wdata1_68 = _RAND_452[63:0];
  _RAND_453 = {2{`RANDOM}};
  recent_wdata1_69 = _RAND_453[63:0];
  _RAND_454 = {2{`RANDOM}};
  recent_wdata1_70 = _RAND_454[63:0];
  _RAND_455 = {2{`RANDOM}};
  recent_wdata1_71 = _RAND_455[63:0];
  _RAND_456 = {2{`RANDOM}};
  recent_wdata1_72 = _RAND_456[63:0];
  _RAND_457 = {2{`RANDOM}};
  recent_wdata1_73 = _RAND_457[63:0];
  _RAND_458 = {2{`RANDOM}};
  recent_wdata1_74 = _RAND_458[63:0];
  _RAND_459 = {2{`RANDOM}};
  recent_wdata1_75 = _RAND_459[63:0];
  _RAND_460 = {2{`RANDOM}};
  recent_wdata1_76 = _RAND_460[63:0];
  _RAND_461 = {2{`RANDOM}};
  recent_wdata1_77 = _RAND_461[63:0];
  _RAND_462 = {2{`RANDOM}};
  recent_wdata1_78 = _RAND_462[63:0];
  _RAND_463 = {2{`RANDOM}};
  recent_wdata1_79 = _RAND_463[63:0];
  _RAND_464 = {2{`RANDOM}};
  recent_wdata1_80 = _RAND_464[63:0];
  _RAND_465 = {2{`RANDOM}};
  recent_wdata1_81 = _RAND_465[63:0];
  _RAND_466 = {2{`RANDOM}};
  recent_wdata1_82 = _RAND_466[63:0];
  _RAND_467 = {2{`RANDOM}};
  recent_wdata1_83 = _RAND_467[63:0];
  _RAND_468 = {2{`RANDOM}};
  recent_wdata1_84 = _RAND_468[63:0];
  _RAND_469 = {2{`RANDOM}};
  recent_wdata1_85 = _RAND_469[63:0];
  _RAND_470 = {2{`RANDOM}};
  recent_wdata1_86 = _RAND_470[63:0];
  _RAND_471 = {2{`RANDOM}};
  recent_wdata1_87 = _RAND_471[63:0];
  _RAND_472 = {2{`RANDOM}};
  recent_wdata1_88 = _RAND_472[63:0];
  _RAND_473 = {2{`RANDOM}};
  recent_wdata1_89 = _RAND_473[63:0];
  _RAND_474 = {2{`RANDOM}};
  recent_wdata1_90 = _RAND_474[63:0];
  _RAND_475 = {2{`RANDOM}};
  recent_wdata1_91 = _RAND_475[63:0];
  _RAND_476 = {2{`RANDOM}};
  recent_wdata1_92 = _RAND_476[63:0];
  _RAND_477 = {2{`RANDOM}};
  recent_wdata1_93 = _RAND_477[63:0];
  _RAND_478 = {2{`RANDOM}};
  recent_wdata1_94 = _RAND_478[63:0];
  _RAND_479 = {2{`RANDOM}};
  recent_wdata1_95 = _RAND_479[63:0];
  _RAND_480 = {2{`RANDOM}};
  recent_wdata1_96 = _RAND_480[63:0];
  _RAND_481 = {2{`RANDOM}};
  recent_wdata1_97 = _RAND_481[63:0];
  _RAND_482 = {2{`RANDOM}};
  recent_wdata1_98 = _RAND_482[63:0];
  _RAND_483 = {2{`RANDOM}};
  recent_wdata1_99 = _RAND_483[63:0];
  _RAND_484 = {2{`RANDOM}};
  recent_wdata1_100 = _RAND_484[63:0];
  _RAND_485 = {2{`RANDOM}};
  recent_wdata1_101 = _RAND_485[63:0];
  _RAND_486 = {2{`RANDOM}};
  recent_wdata1_102 = _RAND_486[63:0];
  _RAND_487 = {2{`RANDOM}};
  recent_wdata1_103 = _RAND_487[63:0];
  _RAND_488 = {2{`RANDOM}};
  recent_wdata1_104 = _RAND_488[63:0];
  _RAND_489 = {2{`RANDOM}};
  recent_wdata1_105 = _RAND_489[63:0];
  _RAND_490 = {2{`RANDOM}};
  recent_wdata1_106 = _RAND_490[63:0];
  _RAND_491 = {2{`RANDOM}};
  recent_wdata1_107 = _RAND_491[63:0];
  _RAND_492 = {2{`RANDOM}};
  recent_wdata1_108 = _RAND_492[63:0];
  _RAND_493 = {2{`RANDOM}};
  recent_wdata1_109 = _RAND_493[63:0];
  _RAND_494 = {2{`RANDOM}};
  recent_wdata1_110 = _RAND_494[63:0];
  _RAND_495 = {2{`RANDOM}};
  recent_wdata1_111 = _RAND_495[63:0];
  _RAND_496 = {2{`RANDOM}};
  recent_wdata1_112 = _RAND_496[63:0];
  _RAND_497 = {2{`RANDOM}};
  recent_wdata1_113 = _RAND_497[63:0];
  _RAND_498 = {2{`RANDOM}};
  recent_wdata1_114 = _RAND_498[63:0];
  _RAND_499 = {2{`RANDOM}};
  recent_wdata1_115 = _RAND_499[63:0];
  _RAND_500 = {2{`RANDOM}};
  recent_wdata1_116 = _RAND_500[63:0];
  _RAND_501 = {2{`RANDOM}};
  recent_wdata1_117 = _RAND_501[63:0];
  _RAND_502 = {2{`RANDOM}};
  recent_wdata1_118 = _RAND_502[63:0];
  _RAND_503 = {2{`RANDOM}};
  recent_wdata1_119 = _RAND_503[63:0];
  _RAND_504 = {2{`RANDOM}};
  recent_wdata1_120 = _RAND_504[63:0];
  _RAND_505 = {2{`RANDOM}};
  recent_wdata1_121 = _RAND_505[63:0];
  _RAND_506 = {2{`RANDOM}};
  recent_wdata1_122 = _RAND_506[63:0];
  _RAND_507 = {2{`RANDOM}};
  recent_wdata1_123 = _RAND_507[63:0];
  _RAND_508 = {2{`RANDOM}};
  recent_wdata1_124 = _RAND_508[63:0];
  _RAND_509 = {2{`RANDOM}};
  recent_wdata1_125 = _RAND_509[63:0];
  _RAND_510 = {2{`RANDOM}};
  recent_wdata1_126 = _RAND_510[63:0];
  _RAND_511 = {2{`RANDOM}};
  recent_wdata1_127 = _RAND_511[63:0];
  _RAND_512 = {1{`RANDOM}};
  tag_0_0 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  tag_0_1 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  tag_0_2 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  tag_0_3 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  tag_0_4 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  tag_0_5 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  tag_0_6 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  tag_0_7 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  tag_0_8 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  tag_0_9 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  tag_0_10 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  tag_0_11 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  tag_0_12 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  tag_0_13 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  tag_0_14 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  tag_0_15 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  tag_0_16 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  tag_0_17 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  tag_0_18 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  tag_0_19 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  tag_0_20 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  tag_0_21 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  tag_0_22 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  tag_0_23 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  tag_0_24 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  tag_0_25 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  tag_0_26 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  tag_0_27 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  tag_0_28 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  tag_0_29 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  tag_0_30 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  tag_0_31 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  tag_0_32 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  tag_0_33 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  tag_0_34 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  tag_0_35 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  tag_0_36 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  tag_0_37 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  tag_0_38 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  tag_0_39 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  tag_0_40 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  tag_0_41 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  tag_0_42 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  tag_0_43 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  tag_0_44 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  tag_0_45 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  tag_0_46 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  tag_0_47 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  tag_0_48 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  tag_0_49 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  tag_0_50 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  tag_0_51 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  tag_0_52 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  tag_0_53 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  tag_0_54 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  tag_0_55 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  tag_0_56 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  tag_0_57 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  tag_0_58 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  tag_0_59 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  tag_0_60 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  tag_0_61 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  tag_0_62 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  tag_0_63 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  tag_0_64 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  tag_0_65 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  tag_0_66 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  tag_0_67 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  tag_0_68 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  tag_0_69 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  tag_0_70 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  tag_0_71 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  tag_0_72 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  tag_0_73 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  tag_0_74 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  tag_0_75 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  tag_0_76 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  tag_0_77 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  tag_0_78 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  tag_0_79 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  tag_0_80 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  tag_0_81 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  tag_0_82 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  tag_0_83 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  tag_0_84 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  tag_0_85 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  tag_0_86 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  tag_0_87 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  tag_0_88 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  tag_0_89 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  tag_0_90 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  tag_0_91 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  tag_0_92 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  tag_0_93 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  tag_0_94 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  tag_0_95 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  tag_0_96 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  tag_0_97 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  tag_0_98 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  tag_0_99 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  tag_0_100 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  tag_0_101 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  tag_0_102 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  tag_0_103 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  tag_0_104 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  tag_0_105 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  tag_0_106 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  tag_0_107 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  tag_0_108 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  tag_0_109 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  tag_0_110 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  tag_0_111 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  tag_0_112 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  tag_0_113 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  tag_0_114 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  tag_0_115 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  tag_0_116 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  tag_0_117 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  tag_0_118 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  tag_0_119 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  tag_0_120 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  tag_0_121 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  tag_0_122 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  tag_0_123 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  tag_0_124 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  tag_0_125 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  tag_0_126 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  tag_0_127 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  tag_1_0 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  tag_1_1 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  tag_1_2 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  tag_1_3 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  tag_1_4 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  tag_1_5 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  tag_1_6 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  tag_1_7 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  tag_1_8 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  tag_1_9 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  tag_1_10 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  tag_1_11 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  tag_1_12 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  tag_1_13 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  tag_1_14 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  tag_1_15 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  tag_1_16 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  tag_1_17 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  tag_1_18 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  tag_1_19 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  tag_1_20 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  tag_1_21 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  tag_1_22 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  tag_1_23 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  tag_1_24 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  tag_1_25 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  tag_1_26 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  tag_1_27 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  tag_1_28 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  tag_1_29 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  tag_1_30 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  tag_1_31 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  tag_1_32 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  tag_1_33 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  tag_1_34 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  tag_1_35 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  tag_1_36 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  tag_1_37 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  tag_1_38 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  tag_1_39 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  tag_1_40 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  tag_1_41 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  tag_1_42 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  tag_1_43 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  tag_1_44 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  tag_1_45 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  tag_1_46 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  tag_1_47 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  tag_1_48 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  tag_1_49 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  tag_1_50 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  tag_1_51 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  tag_1_52 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  tag_1_53 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  tag_1_54 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  tag_1_55 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  tag_1_56 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  tag_1_57 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  tag_1_58 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  tag_1_59 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  tag_1_60 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  tag_1_61 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  tag_1_62 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  tag_1_63 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  tag_1_64 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  tag_1_65 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  tag_1_66 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  tag_1_67 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  tag_1_68 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  tag_1_69 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  tag_1_70 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  tag_1_71 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  tag_1_72 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  tag_1_73 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  tag_1_74 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  tag_1_75 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  tag_1_76 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  tag_1_77 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  tag_1_78 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  tag_1_79 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  tag_1_80 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  tag_1_81 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  tag_1_82 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  tag_1_83 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  tag_1_84 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  tag_1_85 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  tag_1_86 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  tag_1_87 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  tag_1_88 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  tag_1_89 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  tag_1_90 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  tag_1_91 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  tag_1_92 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  tag_1_93 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  tag_1_94 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  tag_1_95 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  tag_1_96 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  tag_1_97 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  tag_1_98 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  tag_1_99 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  tag_1_100 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  tag_1_101 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  tag_1_102 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  tag_1_103 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  tag_1_104 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  tag_1_105 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  tag_1_106 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  tag_1_107 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  tag_1_108 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  tag_1_109 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  tag_1_110 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  tag_1_111 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  tag_1_112 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  tag_1_113 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  tag_1_114 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  tag_1_115 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  tag_1_116 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  tag_1_117 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  tag_1_118 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  tag_1_119 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  tag_1_120 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  tag_1_121 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  tag_1_122 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  tag_1_123 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  tag_1_124 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  tag_1_125 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  tag_1_126 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  tag_1_127 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  valid_0_0 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  valid_0_1 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  valid_0_2 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  valid_0_3 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  valid_0_4 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  valid_0_5 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  valid_0_6 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  valid_0_7 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  valid_0_8 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  valid_0_9 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  valid_0_10 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  valid_0_11 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  valid_0_12 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  valid_0_13 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  valid_0_14 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  valid_0_15 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  valid_0_16 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  valid_0_17 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  valid_0_18 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  valid_0_19 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  valid_0_20 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  valid_0_21 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  valid_0_22 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  valid_0_23 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  valid_0_24 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  valid_0_25 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  valid_0_26 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  valid_0_27 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  valid_0_28 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  valid_0_29 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  valid_0_30 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  valid_0_31 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  valid_0_32 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  valid_0_33 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  valid_0_34 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  valid_0_35 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  valid_0_36 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  valid_0_37 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  valid_0_38 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  valid_0_39 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  valid_0_40 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  valid_0_41 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  valid_0_42 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  valid_0_43 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  valid_0_44 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  valid_0_45 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  valid_0_46 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  valid_0_47 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  valid_0_48 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  valid_0_49 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  valid_0_50 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  valid_0_51 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  valid_0_52 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  valid_0_53 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  valid_0_54 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  valid_0_55 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  valid_0_56 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  valid_0_57 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  valid_0_58 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  valid_0_59 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  valid_0_60 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  valid_0_61 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  valid_0_62 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  valid_0_63 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  valid_0_64 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  valid_0_65 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  valid_0_66 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  valid_0_67 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  valid_0_68 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  valid_0_69 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  valid_0_70 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  valid_0_71 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  valid_0_72 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  valid_0_73 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  valid_0_74 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  valid_0_75 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  valid_0_76 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  valid_0_77 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  valid_0_78 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  valid_0_79 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  valid_0_80 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  valid_0_81 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  valid_0_82 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  valid_0_83 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  valid_0_84 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  valid_0_85 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  valid_0_86 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  valid_0_87 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  valid_0_88 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  valid_0_89 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  valid_0_90 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  valid_0_91 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  valid_0_92 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  valid_0_93 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  valid_0_94 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  valid_0_95 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  valid_0_96 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  valid_0_97 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  valid_0_98 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  valid_0_99 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  valid_0_100 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  valid_0_101 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  valid_0_102 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  valid_0_103 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  valid_0_104 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  valid_0_105 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  valid_0_106 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  valid_0_107 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  valid_0_108 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  valid_0_109 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  valid_0_110 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  valid_0_111 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  valid_0_112 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  valid_0_113 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  valid_0_114 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  valid_0_115 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  valid_0_116 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  valid_0_117 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  valid_0_118 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  valid_0_119 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  valid_0_120 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  valid_0_121 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  valid_0_122 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  valid_0_123 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  valid_0_124 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  valid_0_125 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  valid_0_126 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  valid_0_127 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  valid_1_0 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  valid_1_1 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  valid_1_2 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  valid_1_3 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  valid_1_4 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  valid_1_5 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  valid_1_6 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  valid_1_7 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  valid_1_8 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  valid_1_9 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  valid_1_10 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  valid_1_11 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  valid_1_12 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  valid_1_13 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  valid_1_14 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  valid_1_15 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  valid_1_16 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  valid_1_17 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  valid_1_18 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  valid_1_19 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  valid_1_20 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  valid_1_21 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  valid_1_22 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  valid_1_23 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  valid_1_24 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  valid_1_25 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  valid_1_26 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  valid_1_27 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  valid_1_28 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  valid_1_29 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  valid_1_30 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  valid_1_31 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  valid_1_32 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  valid_1_33 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  valid_1_34 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  valid_1_35 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  valid_1_36 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  valid_1_37 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  valid_1_38 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  valid_1_39 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  valid_1_40 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  valid_1_41 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  valid_1_42 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  valid_1_43 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  valid_1_44 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  valid_1_45 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  valid_1_46 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  valid_1_47 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  valid_1_48 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  valid_1_49 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  valid_1_50 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  valid_1_51 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  valid_1_52 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  valid_1_53 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  valid_1_54 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  valid_1_55 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  valid_1_56 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  valid_1_57 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  valid_1_58 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  valid_1_59 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  valid_1_60 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  valid_1_61 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  valid_1_62 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  valid_1_63 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  valid_1_64 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  valid_1_65 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  valid_1_66 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  valid_1_67 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  valid_1_68 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  valid_1_69 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  valid_1_70 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  valid_1_71 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  valid_1_72 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  valid_1_73 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  valid_1_74 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  valid_1_75 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  valid_1_76 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  valid_1_77 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  valid_1_78 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  valid_1_79 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  valid_1_80 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  valid_1_81 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  valid_1_82 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  valid_1_83 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  valid_1_84 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  valid_1_85 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  valid_1_86 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  valid_1_87 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  valid_1_88 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  valid_1_89 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  valid_1_90 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  valid_1_91 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  valid_1_92 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  valid_1_93 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  valid_1_94 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  valid_1_95 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  valid_1_96 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  valid_1_97 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  valid_1_98 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  valid_1_99 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  valid_1_100 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  valid_1_101 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  valid_1_102 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  valid_1_103 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  valid_1_104 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  valid_1_105 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  valid_1_106 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  valid_1_107 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  valid_1_108 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  valid_1_109 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  valid_1_110 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  valid_1_111 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  valid_1_112 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  valid_1_113 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  valid_1_114 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  valid_1_115 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  valid_1_116 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  valid_1_117 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  valid_1_118 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  valid_1_119 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  valid_1_120 = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  valid_1_121 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  valid_1_122 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  valid_1_123 = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  valid_1_124 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  valid_1_125 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  valid_1_126 = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  valid_1_127 = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  dirty_0_0 = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  dirty_0_1 = _RAND_1025[0:0];
  _RAND_1026 = {1{`RANDOM}};
  dirty_0_2 = _RAND_1026[0:0];
  _RAND_1027 = {1{`RANDOM}};
  dirty_0_3 = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  dirty_0_4 = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  dirty_0_5 = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  dirty_0_6 = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  dirty_0_7 = _RAND_1031[0:0];
  _RAND_1032 = {1{`RANDOM}};
  dirty_0_8 = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  dirty_0_9 = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  dirty_0_10 = _RAND_1034[0:0];
  _RAND_1035 = {1{`RANDOM}};
  dirty_0_11 = _RAND_1035[0:0];
  _RAND_1036 = {1{`RANDOM}};
  dirty_0_12 = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  dirty_0_13 = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  dirty_0_14 = _RAND_1038[0:0];
  _RAND_1039 = {1{`RANDOM}};
  dirty_0_15 = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  dirty_0_16 = _RAND_1040[0:0];
  _RAND_1041 = {1{`RANDOM}};
  dirty_0_17 = _RAND_1041[0:0];
  _RAND_1042 = {1{`RANDOM}};
  dirty_0_18 = _RAND_1042[0:0];
  _RAND_1043 = {1{`RANDOM}};
  dirty_0_19 = _RAND_1043[0:0];
  _RAND_1044 = {1{`RANDOM}};
  dirty_0_20 = _RAND_1044[0:0];
  _RAND_1045 = {1{`RANDOM}};
  dirty_0_21 = _RAND_1045[0:0];
  _RAND_1046 = {1{`RANDOM}};
  dirty_0_22 = _RAND_1046[0:0];
  _RAND_1047 = {1{`RANDOM}};
  dirty_0_23 = _RAND_1047[0:0];
  _RAND_1048 = {1{`RANDOM}};
  dirty_0_24 = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  dirty_0_25 = _RAND_1049[0:0];
  _RAND_1050 = {1{`RANDOM}};
  dirty_0_26 = _RAND_1050[0:0];
  _RAND_1051 = {1{`RANDOM}};
  dirty_0_27 = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  dirty_0_28 = _RAND_1052[0:0];
  _RAND_1053 = {1{`RANDOM}};
  dirty_0_29 = _RAND_1053[0:0];
  _RAND_1054 = {1{`RANDOM}};
  dirty_0_30 = _RAND_1054[0:0];
  _RAND_1055 = {1{`RANDOM}};
  dirty_0_31 = _RAND_1055[0:0];
  _RAND_1056 = {1{`RANDOM}};
  dirty_0_32 = _RAND_1056[0:0];
  _RAND_1057 = {1{`RANDOM}};
  dirty_0_33 = _RAND_1057[0:0];
  _RAND_1058 = {1{`RANDOM}};
  dirty_0_34 = _RAND_1058[0:0];
  _RAND_1059 = {1{`RANDOM}};
  dirty_0_35 = _RAND_1059[0:0];
  _RAND_1060 = {1{`RANDOM}};
  dirty_0_36 = _RAND_1060[0:0];
  _RAND_1061 = {1{`RANDOM}};
  dirty_0_37 = _RAND_1061[0:0];
  _RAND_1062 = {1{`RANDOM}};
  dirty_0_38 = _RAND_1062[0:0];
  _RAND_1063 = {1{`RANDOM}};
  dirty_0_39 = _RAND_1063[0:0];
  _RAND_1064 = {1{`RANDOM}};
  dirty_0_40 = _RAND_1064[0:0];
  _RAND_1065 = {1{`RANDOM}};
  dirty_0_41 = _RAND_1065[0:0];
  _RAND_1066 = {1{`RANDOM}};
  dirty_0_42 = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  dirty_0_43 = _RAND_1067[0:0];
  _RAND_1068 = {1{`RANDOM}};
  dirty_0_44 = _RAND_1068[0:0];
  _RAND_1069 = {1{`RANDOM}};
  dirty_0_45 = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  dirty_0_46 = _RAND_1070[0:0];
  _RAND_1071 = {1{`RANDOM}};
  dirty_0_47 = _RAND_1071[0:0];
  _RAND_1072 = {1{`RANDOM}};
  dirty_0_48 = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  dirty_0_49 = _RAND_1073[0:0];
  _RAND_1074 = {1{`RANDOM}};
  dirty_0_50 = _RAND_1074[0:0];
  _RAND_1075 = {1{`RANDOM}};
  dirty_0_51 = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  dirty_0_52 = _RAND_1076[0:0];
  _RAND_1077 = {1{`RANDOM}};
  dirty_0_53 = _RAND_1077[0:0];
  _RAND_1078 = {1{`RANDOM}};
  dirty_0_54 = _RAND_1078[0:0];
  _RAND_1079 = {1{`RANDOM}};
  dirty_0_55 = _RAND_1079[0:0];
  _RAND_1080 = {1{`RANDOM}};
  dirty_0_56 = _RAND_1080[0:0];
  _RAND_1081 = {1{`RANDOM}};
  dirty_0_57 = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  dirty_0_58 = _RAND_1082[0:0];
  _RAND_1083 = {1{`RANDOM}};
  dirty_0_59 = _RAND_1083[0:0];
  _RAND_1084 = {1{`RANDOM}};
  dirty_0_60 = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  dirty_0_61 = _RAND_1085[0:0];
  _RAND_1086 = {1{`RANDOM}};
  dirty_0_62 = _RAND_1086[0:0];
  _RAND_1087 = {1{`RANDOM}};
  dirty_0_63 = _RAND_1087[0:0];
  _RAND_1088 = {1{`RANDOM}};
  dirty_0_64 = _RAND_1088[0:0];
  _RAND_1089 = {1{`RANDOM}};
  dirty_0_65 = _RAND_1089[0:0];
  _RAND_1090 = {1{`RANDOM}};
  dirty_0_66 = _RAND_1090[0:0];
  _RAND_1091 = {1{`RANDOM}};
  dirty_0_67 = _RAND_1091[0:0];
  _RAND_1092 = {1{`RANDOM}};
  dirty_0_68 = _RAND_1092[0:0];
  _RAND_1093 = {1{`RANDOM}};
  dirty_0_69 = _RAND_1093[0:0];
  _RAND_1094 = {1{`RANDOM}};
  dirty_0_70 = _RAND_1094[0:0];
  _RAND_1095 = {1{`RANDOM}};
  dirty_0_71 = _RAND_1095[0:0];
  _RAND_1096 = {1{`RANDOM}};
  dirty_0_72 = _RAND_1096[0:0];
  _RAND_1097 = {1{`RANDOM}};
  dirty_0_73 = _RAND_1097[0:0];
  _RAND_1098 = {1{`RANDOM}};
  dirty_0_74 = _RAND_1098[0:0];
  _RAND_1099 = {1{`RANDOM}};
  dirty_0_75 = _RAND_1099[0:0];
  _RAND_1100 = {1{`RANDOM}};
  dirty_0_76 = _RAND_1100[0:0];
  _RAND_1101 = {1{`RANDOM}};
  dirty_0_77 = _RAND_1101[0:0];
  _RAND_1102 = {1{`RANDOM}};
  dirty_0_78 = _RAND_1102[0:0];
  _RAND_1103 = {1{`RANDOM}};
  dirty_0_79 = _RAND_1103[0:0];
  _RAND_1104 = {1{`RANDOM}};
  dirty_0_80 = _RAND_1104[0:0];
  _RAND_1105 = {1{`RANDOM}};
  dirty_0_81 = _RAND_1105[0:0];
  _RAND_1106 = {1{`RANDOM}};
  dirty_0_82 = _RAND_1106[0:0];
  _RAND_1107 = {1{`RANDOM}};
  dirty_0_83 = _RAND_1107[0:0];
  _RAND_1108 = {1{`RANDOM}};
  dirty_0_84 = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  dirty_0_85 = _RAND_1109[0:0];
  _RAND_1110 = {1{`RANDOM}};
  dirty_0_86 = _RAND_1110[0:0];
  _RAND_1111 = {1{`RANDOM}};
  dirty_0_87 = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  dirty_0_88 = _RAND_1112[0:0];
  _RAND_1113 = {1{`RANDOM}};
  dirty_0_89 = _RAND_1113[0:0];
  _RAND_1114 = {1{`RANDOM}};
  dirty_0_90 = _RAND_1114[0:0];
  _RAND_1115 = {1{`RANDOM}};
  dirty_0_91 = _RAND_1115[0:0];
  _RAND_1116 = {1{`RANDOM}};
  dirty_0_92 = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  dirty_0_93 = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  dirty_0_94 = _RAND_1118[0:0];
  _RAND_1119 = {1{`RANDOM}};
  dirty_0_95 = _RAND_1119[0:0];
  _RAND_1120 = {1{`RANDOM}};
  dirty_0_96 = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  dirty_0_97 = _RAND_1121[0:0];
  _RAND_1122 = {1{`RANDOM}};
  dirty_0_98 = _RAND_1122[0:0];
  _RAND_1123 = {1{`RANDOM}};
  dirty_0_99 = _RAND_1123[0:0];
  _RAND_1124 = {1{`RANDOM}};
  dirty_0_100 = _RAND_1124[0:0];
  _RAND_1125 = {1{`RANDOM}};
  dirty_0_101 = _RAND_1125[0:0];
  _RAND_1126 = {1{`RANDOM}};
  dirty_0_102 = _RAND_1126[0:0];
  _RAND_1127 = {1{`RANDOM}};
  dirty_0_103 = _RAND_1127[0:0];
  _RAND_1128 = {1{`RANDOM}};
  dirty_0_104 = _RAND_1128[0:0];
  _RAND_1129 = {1{`RANDOM}};
  dirty_0_105 = _RAND_1129[0:0];
  _RAND_1130 = {1{`RANDOM}};
  dirty_0_106 = _RAND_1130[0:0];
  _RAND_1131 = {1{`RANDOM}};
  dirty_0_107 = _RAND_1131[0:0];
  _RAND_1132 = {1{`RANDOM}};
  dirty_0_108 = _RAND_1132[0:0];
  _RAND_1133 = {1{`RANDOM}};
  dirty_0_109 = _RAND_1133[0:0];
  _RAND_1134 = {1{`RANDOM}};
  dirty_0_110 = _RAND_1134[0:0];
  _RAND_1135 = {1{`RANDOM}};
  dirty_0_111 = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  dirty_0_112 = _RAND_1136[0:0];
  _RAND_1137 = {1{`RANDOM}};
  dirty_0_113 = _RAND_1137[0:0];
  _RAND_1138 = {1{`RANDOM}};
  dirty_0_114 = _RAND_1138[0:0];
  _RAND_1139 = {1{`RANDOM}};
  dirty_0_115 = _RAND_1139[0:0];
  _RAND_1140 = {1{`RANDOM}};
  dirty_0_116 = _RAND_1140[0:0];
  _RAND_1141 = {1{`RANDOM}};
  dirty_0_117 = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  dirty_0_118 = _RAND_1142[0:0];
  _RAND_1143 = {1{`RANDOM}};
  dirty_0_119 = _RAND_1143[0:0];
  _RAND_1144 = {1{`RANDOM}};
  dirty_0_120 = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  dirty_0_121 = _RAND_1145[0:0];
  _RAND_1146 = {1{`RANDOM}};
  dirty_0_122 = _RAND_1146[0:0];
  _RAND_1147 = {1{`RANDOM}};
  dirty_0_123 = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  dirty_0_124 = _RAND_1148[0:0];
  _RAND_1149 = {1{`RANDOM}};
  dirty_0_125 = _RAND_1149[0:0];
  _RAND_1150 = {1{`RANDOM}};
  dirty_0_126 = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  dirty_0_127 = _RAND_1151[0:0];
  _RAND_1152 = {1{`RANDOM}};
  dirty_1_0 = _RAND_1152[0:0];
  _RAND_1153 = {1{`RANDOM}};
  dirty_1_1 = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  dirty_1_2 = _RAND_1154[0:0];
  _RAND_1155 = {1{`RANDOM}};
  dirty_1_3 = _RAND_1155[0:0];
  _RAND_1156 = {1{`RANDOM}};
  dirty_1_4 = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  dirty_1_5 = _RAND_1157[0:0];
  _RAND_1158 = {1{`RANDOM}};
  dirty_1_6 = _RAND_1158[0:0];
  _RAND_1159 = {1{`RANDOM}};
  dirty_1_7 = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  dirty_1_8 = _RAND_1160[0:0];
  _RAND_1161 = {1{`RANDOM}};
  dirty_1_9 = _RAND_1161[0:0];
  _RAND_1162 = {1{`RANDOM}};
  dirty_1_10 = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  dirty_1_11 = _RAND_1163[0:0];
  _RAND_1164 = {1{`RANDOM}};
  dirty_1_12 = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  dirty_1_13 = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  dirty_1_14 = _RAND_1166[0:0];
  _RAND_1167 = {1{`RANDOM}};
  dirty_1_15 = _RAND_1167[0:0];
  _RAND_1168 = {1{`RANDOM}};
  dirty_1_16 = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  dirty_1_17 = _RAND_1169[0:0];
  _RAND_1170 = {1{`RANDOM}};
  dirty_1_18 = _RAND_1170[0:0];
  _RAND_1171 = {1{`RANDOM}};
  dirty_1_19 = _RAND_1171[0:0];
  _RAND_1172 = {1{`RANDOM}};
  dirty_1_20 = _RAND_1172[0:0];
  _RAND_1173 = {1{`RANDOM}};
  dirty_1_21 = _RAND_1173[0:0];
  _RAND_1174 = {1{`RANDOM}};
  dirty_1_22 = _RAND_1174[0:0];
  _RAND_1175 = {1{`RANDOM}};
  dirty_1_23 = _RAND_1175[0:0];
  _RAND_1176 = {1{`RANDOM}};
  dirty_1_24 = _RAND_1176[0:0];
  _RAND_1177 = {1{`RANDOM}};
  dirty_1_25 = _RAND_1177[0:0];
  _RAND_1178 = {1{`RANDOM}};
  dirty_1_26 = _RAND_1178[0:0];
  _RAND_1179 = {1{`RANDOM}};
  dirty_1_27 = _RAND_1179[0:0];
  _RAND_1180 = {1{`RANDOM}};
  dirty_1_28 = _RAND_1180[0:0];
  _RAND_1181 = {1{`RANDOM}};
  dirty_1_29 = _RAND_1181[0:0];
  _RAND_1182 = {1{`RANDOM}};
  dirty_1_30 = _RAND_1182[0:0];
  _RAND_1183 = {1{`RANDOM}};
  dirty_1_31 = _RAND_1183[0:0];
  _RAND_1184 = {1{`RANDOM}};
  dirty_1_32 = _RAND_1184[0:0];
  _RAND_1185 = {1{`RANDOM}};
  dirty_1_33 = _RAND_1185[0:0];
  _RAND_1186 = {1{`RANDOM}};
  dirty_1_34 = _RAND_1186[0:0];
  _RAND_1187 = {1{`RANDOM}};
  dirty_1_35 = _RAND_1187[0:0];
  _RAND_1188 = {1{`RANDOM}};
  dirty_1_36 = _RAND_1188[0:0];
  _RAND_1189 = {1{`RANDOM}};
  dirty_1_37 = _RAND_1189[0:0];
  _RAND_1190 = {1{`RANDOM}};
  dirty_1_38 = _RAND_1190[0:0];
  _RAND_1191 = {1{`RANDOM}};
  dirty_1_39 = _RAND_1191[0:0];
  _RAND_1192 = {1{`RANDOM}};
  dirty_1_40 = _RAND_1192[0:0];
  _RAND_1193 = {1{`RANDOM}};
  dirty_1_41 = _RAND_1193[0:0];
  _RAND_1194 = {1{`RANDOM}};
  dirty_1_42 = _RAND_1194[0:0];
  _RAND_1195 = {1{`RANDOM}};
  dirty_1_43 = _RAND_1195[0:0];
  _RAND_1196 = {1{`RANDOM}};
  dirty_1_44 = _RAND_1196[0:0];
  _RAND_1197 = {1{`RANDOM}};
  dirty_1_45 = _RAND_1197[0:0];
  _RAND_1198 = {1{`RANDOM}};
  dirty_1_46 = _RAND_1198[0:0];
  _RAND_1199 = {1{`RANDOM}};
  dirty_1_47 = _RAND_1199[0:0];
  _RAND_1200 = {1{`RANDOM}};
  dirty_1_48 = _RAND_1200[0:0];
  _RAND_1201 = {1{`RANDOM}};
  dirty_1_49 = _RAND_1201[0:0];
  _RAND_1202 = {1{`RANDOM}};
  dirty_1_50 = _RAND_1202[0:0];
  _RAND_1203 = {1{`RANDOM}};
  dirty_1_51 = _RAND_1203[0:0];
  _RAND_1204 = {1{`RANDOM}};
  dirty_1_52 = _RAND_1204[0:0];
  _RAND_1205 = {1{`RANDOM}};
  dirty_1_53 = _RAND_1205[0:0];
  _RAND_1206 = {1{`RANDOM}};
  dirty_1_54 = _RAND_1206[0:0];
  _RAND_1207 = {1{`RANDOM}};
  dirty_1_55 = _RAND_1207[0:0];
  _RAND_1208 = {1{`RANDOM}};
  dirty_1_56 = _RAND_1208[0:0];
  _RAND_1209 = {1{`RANDOM}};
  dirty_1_57 = _RAND_1209[0:0];
  _RAND_1210 = {1{`RANDOM}};
  dirty_1_58 = _RAND_1210[0:0];
  _RAND_1211 = {1{`RANDOM}};
  dirty_1_59 = _RAND_1211[0:0];
  _RAND_1212 = {1{`RANDOM}};
  dirty_1_60 = _RAND_1212[0:0];
  _RAND_1213 = {1{`RANDOM}};
  dirty_1_61 = _RAND_1213[0:0];
  _RAND_1214 = {1{`RANDOM}};
  dirty_1_62 = _RAND_1214[0:0];
  _RAND_1215 = {1{`RANDOM}};
  dirty_1_63 = _RAND_1215[0:0];
  _RAND_1216 = {1{`RANDOM}};
  dirty_1_64 = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  dirty_1_65 = _RAND_1217[0:0];
  _RAND_1218 = {1{`RANDOM}};
  dirty_1_66 = _RAND_1218[0:0];
  _RAND_1219 = {1{`RANDOM}};
  dirty_1_67 = _RAND_1219[0:0];
  _RAND_1220 = {1{`RANDOM}};
  dirty_1_68 = _RAND_1220[0:0];
  _RAND_1221 = {1{`RANDOM}};
  dirty_1_69 = _RAND_1221[0:0];
  _RAND_1222 = {1{`RANDOM}};
  dirty_1_70 = _RAND_1222[0:0];
  _RAND_1223 = {1{`RANDOM}};
  dirty_1_71 = _RAND_1223[0:0];
  _RAND_1224 = {1{`RANDOM}};
  dirty_1_72 = _RAND_1224[0:0];
  _RAND_1225 = {1{`RANDOM}};
  dirty_1_73 = _RAND_1225[0:0];
  _RAND_1226 = {1{`RANDOM}};
  dirty_1_74 = _RAND_1226[0:0];
  _RAND_1227 = {1{`RANDOM}};
  dirty_1_75 = _RAND_1227[0:0];
  _RAND_1228 = {1{`RANDOM}};
  dirty_1_76 = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  dirty_1_77 = _RAND_1229[0:0];
  _RAND_1230 = {1{`RANDOM}};
  dirty_1_78 = _RAND_1230[0:0];
  _RAND_1231 = {1{`RANDOM}};
  dirty_1_79 = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  dirty_1_80 = _RAND_1232[0:0];
  _RAND_1233 = {1{`RANDOM}};
  dirty_1_81 = _RAND_1233[0:0];
  _RAND_1234 = {1{`RANDOM}};
  dirty_1_82 = _RAND_1234[0:0];
  _RAND_1235 = {1{`RANDOM}};
  dirty_1_83 = _RAND_1235[0:0];
  _RAND_1236 = {1{`RANDOM}};
  dirty_1_84 = _RAND_1236[0:0];
  _RAND_1237 = {1{`RANDOM}};
  dirty_1_85 = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  dirty_1_86 = _RAND_1238[0:0];
  _RAND_1239 = {1{`RANDOM}};
  dirty_1_87 = _RAND_1239[0:0];
  _RAND_1240 = {1{`RANDOM}};
  dirty_1_88 = _RAND_1240[0:0];
  _RAND_1241 = {1{`RANDOM}};
  dirty_1_89 = _RAND_1241[0:0];
  _RAND_1242 = {1{`RANDOM}};
  dirty_1_90 = _RAND_1242[0:0];
  _RAND_1243 = {1{`RANDOM}};
  dirty_1_91 = _RAND_1243[0:0];
  _RAND_1244 = {1{`RANDOM}};
  dirty_1_92 = _RAND_1244[0:0];
  _RAND_1245 = {1{`RANDOM}};
  dirty_1_93 = _RAND_1245[0:0];
  _RAND_1246 = {1{`RANDOM}};
  dirty_1_94 = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  dirty_1_95 = _RAND_1247[0:0];
  _RAND_1248 = {1{`RANDOM}};
  dirty_1_96 = _RAND_1248[0:0];
  _RAND_1249 = {1{`RANDOM}};
  dirty_1_97 = _RAND_1249[0:0];
  _RAND_1250 = {1{`RANDOM}};
  dirty_1_98 = _RAND_1250[0:0];
  _RAND_1251 = {1{`RANDOM}};
  dirty_1_99 = _RAND_1251[0:0];
  _RAND_1252 = {1{`RANDOM}};
  dirty_1_100 = _RAND_1252[0:0];
  _RAND_1253 = {1{`RANDOM}};
  dirty_1_101 = _RAND_1253[0:0];
  _RAND_1254 = {1{`RANDOM}};
  dirty_1_102 = _RAND_1254[0:0];
  _RAND_1255 = {1{`RANDOM}};
  dirty_1_103 = _RAND_1255[0:0];
  _RAND_1256 = {1{`RANDOM}};
  dirty_1_104 = _RAND_1256[0:0];
  _RAND_1257 = {1{`RANDOM}};
  dirty_1_105 = _RAND_1257[0:0];
  _RAND_1258 = {1{`RANDOM}};
  dirty_1_106 = _RAND_1258[0:0];
  _RAND_1259 = {1{`RANDOM}};
  dirty_1_107 = _RAND_1259[0:0];
  _RAND_1260 = {1{`RANDOM}};
  dirty_1_108 = _RAND_1260[0:0];
  _RAND_1261 = {1{`RANDOM}};
  dirty_1_109 = _RAND_1261[0:0];
  _RAND_1262 = {1{`RANDOM}};
  dirty_1_110 = _RAND_1262[0:0];
  _RAND_1263 = {1{`RANDOM}};
  dirty_1_111 = _RAND_1263[0:0];
  _RAND_1264 = {1{`RANDOM}};
  dirty_1_112 = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  dirty_1_113 = _RAND_1265[0:0];
  _RAND_1266 = {1{`RANDOM}};
  dirty_1_114 = _RAND_1266[0:0];
  _RAND_1267 = {1{`RANDOM}};
  dirty_1_115 = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  dirty_1_116 = _RAND_1268[0:0];
  _RAND_1269 = {1{`RANDOM}};
  dirty_1_117 = _RAND_1269[0:0];
  _RAND_1270 = {1{`RANDOM}};
  dirty_1_118 = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  dirty_1_119 = _RAND_1271[0:0];
  _RAND_1272 = {1{`RANDOM}};
  dirty_1_120 = _RAND_1272[0:0];
  _RAND_1273 = {1{`RANDOM}};
  dirty_1_121 = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  dirty_1_122 = _RAND_1274[0:0];
  _RAND_1275 = {1{`RANDOM}};
  dirty_1_123 = _RAND_1275[0:0];
  _RAND_1276 = {1{`RANDOM}};
  dirty_1_124 = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  dirty_1_125 = _RAND_1277[0:0];
  _RAND_1278 = {1{`RANDOM}};
  dirty_1_126 = _RAND_1278[0:0];
  _RAND_1279 = {1{`RANDOM}};
  dirty_1_127 = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  way0_hit = _RAND_1280[0:0];
  _RAND_1281 = {1{`RANDOM}};
  way1_hit = _RAND_1281[0:0];
  _RAND_1282 = {2{`RANDOM}};
  write_back_data = _RAND_1282[63:0];
  _RAND_1283 = {1{`RANDOM}};
  write_back_addr = _RAND_1283[31:0];
  _RAND_1284 = {1{`RANDOM}};
  unuse_way = _RAND_1284[1:0];
  _RAND_1285 = {2{`RANDOM}};
  receive_data = _RAND_1285[63:0];
  _RAND_1286 = {1{`RANDOM}};
  quene = _RAND_1286[0:0];
  _RAND_1287 = {1{`RANDOM}};
  state = _RAND_1287[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IDU(
  input  [31:0] io_inst,
  output [31:0] io_inst_now,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2,
  output [4:0]  io_rd,
  output [63:0] io_imm,
  output        io_ctrl_sign_reg_write,
  output        io_ctrl_sign_csr_write,
  output        io_ctrl_sign_src2_is_imm,
  output        io_ctrl_sign_src1_is_pc,
  output        io_ctrl_sign_Writemem_en,
  output        io_ctrl_sign_Readmem_en,
  output [7:0]  io_ctrl_sign_Wmask
);
  wire [4:0] rd = io_inst[11:7]; // @[IDU.scala 150:15]
  wire [31:0] _inst_type_T = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_1 = 32'h13 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_2 = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_3 = 32'h17 == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_5 = 32'h37 == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_7 = 32'h6f == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_9 = 32'h67 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_11 = 32'h3023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_13 = 32'h3013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_15 = 32'h2003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_16 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_17 = 32'h3b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_19 = 32'h40000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_21 = 32'h1063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_23 = 32'h63 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_25 = 32'h3003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_27 = 32'h1b == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_29 = 32'h33 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_30 = io_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_31 = 32'h40005013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_33 = 32'h4003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_35 = 32'h1023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_37 = 32'h23 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_39 = 32'h6033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_41 = 32'h4013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_43 = 32'h7033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_45 = 32'h7013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_47 = 32'h4000003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_49 = 32'h103b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_51 = 32'h1013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_53 = 32'h5013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_55 = 32'h101b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_57 = 32'h4000501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_59 = 32'h501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_61 = 32'h4000503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_63 = 32'h503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_65 = 32'h3033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_67 = 32'h2033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_69 = 32'h5063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_71 = 32'h4063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_73 = 32'h6063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_75 = 32'h2023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_77 = 32'h1003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_79 = 32'h5003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_81 = 32'h2000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_83 = 32'h200003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_85 = 32'h200403b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_87 = 32'h200603b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_89 = 32'h4033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_91 = 32'h6013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_93 = 32'h2005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_95 = 32'h2004033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_97 = 32'h200503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_99 = 32'h200703b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_101 = 32'h2007033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_103 = 32'h2006033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_105 = 32'h1033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_107 = 32'h5033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_109 = 32'h40005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_111 = 32'h2013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_113 = 32'h6003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_115 = 32'h3 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_117 = 32'h7063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_119 = 32'h73 == io_inst; // @[Lookup.scala 31:38]
  wire  _inst_type_T_121 = 32'h1073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_123 = 32'h2073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_125 = 32'h3073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [6:0] _inst_type_T_126 = _inst_type_T_125 ? 7'h40 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_127 = _inst_type_T_123 ? 7'h40 : _inst_type_T_126; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_128 = _inst_type_T_121 ? 7'h40 : _inst_type_T_127; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_129 = _inst_type_T_119 ? 7'h40 : _inst_type_T_128; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_130 = _inst_type_T_117 ? 7'h45 : _inst_type_T_129; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_131 = _inst_type_T_115 ? 7'h40 : _inst_type_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_132 = _inst_type_T_113 ? 7'h40 : _inst_type_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_133 = _inst_type_T_111 ? 7'h40 : _inst_type_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_134 = _inst_type_T_109 ? 7'h41 : _inst_type_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_135 = _inst_type_T_107 ? 7'h41 : _inst_type_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_136 = _inst_type_T_105 ? 7'h41 : _inst_type_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_137 = _inst_type_T_103 ? 7'h41 : _inst_type_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_138 = _inst_type_T_101 ? 7'h41 : _inst_type_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_139 = _inst_type_T_99 ? 7'h41 : _inst_type_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_140 = _inst_type_T_97 ? 7'h41 : _inst_type_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_141 = _inst_type_T_95 ? 7'h41 : _inst_type_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_142 = _inst_type_T_93 ? 7'h41 : _inst_type_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_143 = _inst_type_T_91 ? 7'h40 : _inst_type_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_144 = _inst_type_T_89 ? 7'h41 : _inst_type_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_145 = _inst_type_T_87 ? 7'h41 : _inst_type_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_146 = _inst_type_T_85 ? 7'h41 : _inst_type_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_147 = _inst_type_T_83 ? 7'h41 : _inst_type_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_148 = _inst_type_T_81 ? 7'h41 : _inst_type_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_149 = _inst_type_T_79 ? 7'h40 : _inst_type_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_150 = _inst_type_T_77 ? 7'h40 : _inst_type_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_151 = _inst_type_T_75 ? 7'h44 : _inst_type_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_152 = _inst_type_T_73 ? 7'h45 : _inst_type_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_153 = _inst_type_T_71 ? 7'h45 : _inst_type_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_154 = _inst_type_T_69 ? 7'h45 : _inst_type_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_155 = _inst_type_T_67 ? 7'h41 : _inst_type_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_156 = _inst_type_T_65 ? 7'h41 : _inst_type_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_157 = _inst_type_T_63 ? 7'h41 : _inst_type_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_158 = _inst_type_T_61 ? 7'h41 : _inst_type_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_159 = _inst_type_T_59 ? 7'h40 : _inst_type_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_160 = _inst_type_T_57 ? 7'h40 : _inst_type_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_161 = _inst_type_T_55 ? 7'h40 : _inst_type_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_162 = _inst_type_T_53 ? 7'h40 : _inst_type_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_163 = _inst_type_T_51 ? 7'h40 : _inst_type_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_164 = _inst_type_T_49 ? 7'h41 : _inst_type_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_165 = _inst_type_T_47 ? 7'h41 : _inst_type_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_166 = _inst_type_T_45 ? 7'h40 : _inst_type_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_167 = _inst_type_T_43 ? 7'h41 : _inst_type_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_168 = _inst_type_T_41 ? 7'h40 : _inst_type_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_169 = _inst_type_T_39 ? 7'h41 : _inst_type_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_170 = _inst_type_T_37 ? 7'h44 : _inst_type_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_171 = _inst_type_T_35 ? 7'h44 : _inst_type_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_172 = _inst_type_T_33 ? 7'h40 : _inst_type_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_173 = _inst_type_T_31 ? 7'h40 : _inst_type_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_174 = _inst_type_T_29 ? 7'h41 : _inst_type_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_175 = _inst_type_T_27 ? 7'h40 : _inst_type_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_176 = _inst_type_T_25 ? 7'h40 : _inst_type_T_175; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_177 = _inst_type_T_23 ? 7'h45 : _inst_type_T_176; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_178 = _inst_type_T_21 ? 7'h45 : _inst_type_T_177; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_179 = _inst_type_T_19 ? 7'h41 : _inst_type_T_178; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_180 = _inst_type_T_17 ? 7'h41 : _inst_type_T_179; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_181 = _inst_type_T_15 ? 7'h40 : _inst_type_T_180; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_182 = _inst_type_T_13 ? 7'h40 : _inst_type_T_181; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_183 = _inst_type_T_11 ? 7'h44 : _inst_type_T_182; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_184 = _inst_type_T_9 ? 7'h40 : _inst_type_T_183; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_185 = _inst_type_T_7 ? 7'h43 : _inst_type_T_184; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_186 = _inst_type_T_5 ? 7'h42 : _inst_type_T_185; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_187 = _inst_type_T_3 ? 7'h42 : _inst_type_T_186; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_188 = _inst_type_T_1 ? 7'h40 : _inst_type_T_187; // @[Lookup.scala 34:39]
  wire [11:0] imm_imm = io_inst[31:20]; // @[IDU.scala 24:23]
  wire [51:0] _imm_T_2 = imm_imm[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_3 = {_imm_T_2,imm_imm}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_1 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21]}; // @[Cat.scala 31:58]
  wire [42:0] _imm_T_6 = imm_imm_1[19] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_7 = {_imm_T_6,io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_2 = io_inst[31:12]; // @[IDU.scala 28:23]
  wire [31:0] _imm_T_10 = imm_imm_2[19] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_12 = {_imm_T_10,imm_imm_2,12'h0}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_3 = {io_inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [51:0] _imm_T_15 = imm_imm_3[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_16 = {_imm_T_15,io_inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_4 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8]}; // @[Cat.scala 31:58]
  wire [50:0] _imm_T_19 = imm_imm_4[11] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_20 = {_imm_T_19,io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] inst_type = {{25'd0}, _inst_type_T_188}; // @[IDU.scala 133:25 152:15]
  wire [63:0] _imm_T_22 = 32'h40 == inst_type ? _imm_T_3 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_24 = 32'h43 == inst_type ? _imm_T_7 : _imm_T_22; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_26 = 32'h42 == inst_type ? _imm_T_12 : _imm_T_24; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_28 = 32'h44 == inst_type ? _imm_T_16 : _imm_T_26; // @[Mux.scala 81:58]
  wire  _inst_now_T_3 = 32'h100073 == io_inst; // @[Lookup.scala 31:38]
  wire  _inst_now_T_123 = 32'h30200073 == io_inst; // @[Lookup.scala 31:38]
  wire [6:0] _inst_now_T_130 = _inst_type_T_125 ? 7'h47 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_131 = _inst_type_T_123 ? 7'h46 : _inst_now_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_132 = _inst_type_T_121 ? 7'h3f : _inst_now_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_133 = _inst_now_T_123 ? 7'h3e : _inst_now_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_134 = _inst_type_T_119 ? 7'h3d : _inst_now_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_135 = _inst_type_T_117 ? 7'h3c : _inst_now_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_136 = _inst_type_T_115 ? 7'h3b : _inst_now_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_137 = _inst_type_T_113 ? 7'h3a : _inst_now_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_138 = _inst_type_T_111 ? 7'h36 : _inst_now_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_139 = _inst_type_T_109 ? 7'h39 : _inst_now_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_140 = _inst_type_T_107 ? 7'h38 : _inst_now_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_141 = _inst_type_T_105 ? 7'h37 : _inst_now_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_142 = _inst_type_T_103 ? 7'h34 : _inst_now_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_143 = _inst_type_T_101 ? 7'h33 : _inst_now_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_144 = _inst_type_T_99 ? 7'h32 : _inst_now_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_145 = _inst_type_T_97 ? 7'h35 : _inst_now_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_146 = _inst_type_T_95 ? 7'h31 : _inst_now_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_147 = _inst_type_T_93 ? 7'h30 : _inst_now_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_148 = _inst_type_T_91 ? 7'h2f : _inst_now_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_149 = _inst_type_T_89 ? 7'h2e : _inst_now_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_150 = _inst_type_T_87 ? 7'h14 : _inst_now_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_151 = _inst_type_T_85 ? 7'h13 : _inst_now_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_152 = _inst_type_T_83 ? 7'h12 : _inst_now_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_153 = _inst_type_T_81 ? 7'h11 : _inst_now_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_154 = _inst_type_T_79 ? 7'h25 : _inst_now_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_155 = _inst_type_T_77 ? 7'h24 : _inst_now_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_156 = _inst_type_T_75 ? 7'h27 : _inst_now_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_157 = _inst_type_T_73 ? 7'h2d : _inst_now_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_158 = _inst_type_T_71 ? 7'h2c : _inst_now_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_159 = _inst_type_T_69 ? 7'h2b : _inst_now_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_160 = _inst_type_T_67 ? 7'h1f : _inst_now_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_161 = _inst_type_T_65 ? 7'h1e : _inst_now_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_162 = _inst_type_T_63 ? 7'h1d : _inst_now_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_163 = _inst_type_T_61 ? 7'h1c : _inst_now_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_164 = _inst_type_T_59 ? 7'h1b : _inst_now_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_165 = _inst_type_T_57 ? 7'h1a : _inst_now_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_166 = _inst_type_T_55 ? 7'h19 : _inst_now_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_167 = _inst_type_T_53 ? 7'h18 : _inst_now_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_168 = _inst_type_T_51 ? 7'h17 : _inst_now_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_169 = _inst_type_T_49 ? 7'h16 : _inst_now_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_170 = _inst_type_T_47 ? 7'hd : _inst_now_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_171 = _inst_type_T_45 ? 7'h9 : _inst_now_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_172 = _inst_type_T_43 ? 7'h8 : _inst_now_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_173 = _inst_type_T_41 ? 7'ha : _inst_now_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_174 = _inst_type_T_39 ? 7'hb : _inst_now_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_175 = _inst_type_T_37 ? 7'h28 : _inst_now_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_176 = _inst_type_T_35 ? 7'h26 : _inst_now_T_175; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_177 = _inst_type_T_33 ? 7'h23 : _inst_now_T_176; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_178 = _inst_type_T_31 ? 7'h15 : _inst_now_T_177; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_179 = _inst_type_T_29 ? 7'hf : _inst_now_T_178; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_180 = _inst_type_T_27 ? 7'h10 : _inst_now_T_179; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_181 = _inst_type_T_25 ? 7'h22 : _inst_now_T_180; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_182 = _inst_type_T_23 ? 7'h29 : _inst_now_T_181; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_183 = _inst_type_T_21 ? 7'h2a : _inst_now_T_182; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_184 = _inst_type_T_19 ? 7'he : _inst_now_T_183; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_185 = _inst_type_T_17 ? 7'hc : _inst_now_T_184; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_186 = _inst_type_T_15 ? 7'h21 : _inst_now_T_185; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_187 = _inst_type_T_13 ? 7'h20 : _inst_now_T_186; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_188 = _inst_type_T_11 ? 7'h7 : _inst_now_T_187; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_189 = _inst_type_T_9 ? 7'h6 : _inst_now_T_188; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_190 = _inst_type_T_7 ? 7'h5 : _inst_now_T_189; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_191 = _inst_type_T_5 ? 7'h4 : _inst_now_T_190; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_192 = _inst_type_T_3 ? 7'h3 : _inst_now_T_191; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_193 = _inst_now_T_3 ? 7'h2 : _inst_now_T_192; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_194 = _inst_type_T_1 ? 7'h1 : _inst_now_T_193; // @[Lookup.scala 34:39]
  wire  _reg_write_T_26 = _inst_now_T_123 ? 1'h0 : 1'h1; // @[Lookup.scala 34:39]
  wire  _reg_write_T_27 = _inst_type_T_119 ? 1'h0 : _reg_write_T_26; // @[Lookup.scala 34:39]
  wire  _reg_write_T_28 = _inst_type_T_117 ? 1'h0 : _reg_write_T_27; // @[Lookup.scala 34:39]
  wire  _reg_write_T_29 = _inst_type_T_73 ? 1'h0 : _reg_write_T_28; // @[Lookup.scala 34:39]
  wire  _reg_write_T_30 = _inst_type_T_71 ? 1'h0 : _reg_write_T_29; // @[Lookup.scala 34:39]
  wire  _reg_write_T_31 = _inst_type_T_69 ? 1'h0 : _reg_write_T_30; // @[Lookup.scala 34:39]
  wire  _reg_write_T_32 = _inst_type_T_23 ? 1'h0 : _reg_write_T_31; // @[Lookup.scala 34:39]
  wire  _reg_write_T_33 = _inst_type_T_21 ? 1'h0 : _reg_write_T_32; // @[Lookup.scala 34:39]
  wire  _reg_write_T_34 = _inst_type_T_75 ? 1'h0 : _reg_write_T_33; // @[Lookup.scala 34:39]
  wire  _reg_write_T_35 = _inst_type_T_37 ? 1'h0 : _reg_write_T_34; // @[Lookup.scala 34:39]
  wire  _reg_write_T_36 = _inst_type_T_35 ? 1'h0 : _reg_write_T_35; // @[Lookup.scala 34:39]
  wire  _reg_write_T_37 = _inst_type_T_11 ? 1'h0 : _reg_write_T_36; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_8 = _inst_type_T_75 ? 4'hf : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_9 = _inst_type_T_37 ? 4'h1 : _Wmask_T_8; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_10 = _inst_type_T_35 ? 4'h3 : _Wmask_T_9; // @[Lookup.scala 34:39]
  assign io_inst_now = {{25'd0}, _inst_now_T_194}; // @[IDU.scala 132:24 226:14]
  assign io_rs1 = io_inst[19:15]; // @[IDU.scala 149:16]
  assign io_rs2 = io_inst[24:20]; // @[IDU.scala 148:16]
  assign io_rd = io_inst[11:7]; // @[IDU.scala 150:15]
  assign io_imm = 32'h45 == inst_type ? _imm_T_20 : _imm_T_28; // @[Mux.scala 81:58]
  assign io_ctrl_sign_reg_write = _inst_now_T_3 ? 1'h0 : _reg_write_T_37; // @[Lookup.scala 34:39]
  assign io_ctrl_sign_csr_write = _inst_type_T_121 | (_inst_type_T_123 | _inst_type_T_125); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_src2_is_imm = 32'h45 == inst_type | (32'h43 == inst_type | (32'h44 == inst_type | (32'h42 ==
    inst_type | 32'h40 == inst_type))); // @[Mux.scala 81:58]
  assign io_ctrl_sign_src1_is_pc = _inst_type_T_7 | (_inst_type_T_3 | (_inst_type_T_21 | (_inst_type_T_23 | (
    _inst_type_T_69 | (_inst_type_T_71 | (_inst_type_T_73 | _inst_type_T_117)))))); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Writemem_en = 32'h44 == inst_type; // @[Mux.scala 81:61]
  assign io_ctrl_sign_Readmem_en = _inst_type_T_25 | (_inst_type_T_15 | (_inst_type_T_113 | (_inst_type_T_77 | (
    _inst_type_T_79 | (_inst_type_T_115 | _inst_type_T_33))))); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Wmask = _inst_type_T_11 ? 8'hff : {{4'd0}, _Wmask_T_10}; // @[Lookup.scala 34:39]
endmodule
module EXU_AXI(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  output [63:0] io_pc_next,
  input  [31:0] io_inst_now,
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [4:0]  io_rd,
  input  [63:0] io_imm,
  input         io_ctrl_sign_reg_write,
  input         io_ctrl_sign_csr_write,
  input         io_ctrl_sign_src2_is_imm,
  input         io_ctrl_sign_src1_is_pc,
  input         io_ctrl_sign_Writemem_en,
  input         io_ctrl_sign_Readmem_en,
  input  [7:0]  io_ctrl_sign_Wmask,
  output [63:0] io_res2rd,
  input         io_inst_valid,
  output        io_inst_store,
  output        io_inst_load,
  output [31:0] io_Mem_addr,
  input  [63:0] io_Mem_rdata,
  output [63:0] io_Mem_wdata,
  output [7:0]  io_Mem_wstrb,
  input         io_rdata_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] Regfile [0:31]; // @[EXU_AXI.scala 37:22]
  wire  Regfile_src1_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_src1_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_src1_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_src2_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_src2_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_src2_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_4_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_MPORT_4_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_MPORT_4_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_1_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_1_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_1_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_2_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_2_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_2_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_3_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_3_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_3_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_4_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_4_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_4_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_5_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_5_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_5_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_6_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_6_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_6_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_7_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_7_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_7_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_8_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_8_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_8_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_9_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_9_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_9_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_10_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_10_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_10_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_11_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_11_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_11_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_0_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_0_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_0_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_1_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_1_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_1_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_2_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_2_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_2_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_3_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_3_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_3_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_4_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_4_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_4_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_5_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_5_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_5_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_6_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_6_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_6_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_7_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_7_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_7_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_8_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_8_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_8_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_9_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_9_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_9_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_10_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_10_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_10_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_11_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_11_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_11_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_12_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_12_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_12_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_13_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_13_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_13_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_14_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_14_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_14_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_15_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_15_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_15_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_16_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_16_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_16_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_17_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_17_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_17_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_18_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_18_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_18_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_19_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_19_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_19_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_20_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_20_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_20_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_21_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_21_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_21_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_22_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_22_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_22_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_23_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_23_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_23_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_24_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_24_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_24_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_25_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_25_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_25_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_26_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_26_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_26_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_27_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_27_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_27_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_28_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_28_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_28_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_29_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_29_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_29_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_30_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_30_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_30_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_31_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_31_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_31_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_1_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_1_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_1_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_2_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_2_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_2_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_3_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_3_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_3_data; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_mask; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_en; // @[EXU_AXI.scala 37:22]
  reg [63:0] CSR_Reg [0:3]; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_2_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_2_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_2_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_csr_wdata_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_csr_wdata_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_csr_wdata_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_csr_wdata_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_csr_wdata_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_csr_wdata_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_2_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_2_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_2_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_5_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_5_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_5_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_7_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_7_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_7_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_j_pc_MPORT_12_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_j_pc_MPORT_12_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_j_pc_MPORT_12_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_j_pc_MPORT_13_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_j_pc_MPORT_13_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_j_pc_MPORT_13_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_0_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_1_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_2_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_1_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_3_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_3_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_3_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_3_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_6_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_6_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_6_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_6_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] reg_trace_input_reg_0; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_1; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_2; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_3; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_4; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_5; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_6; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_7; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_8; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_9; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_10; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_11; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_12; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_13; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_14; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_15; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_16; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_17; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_18; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_19; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_20; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_21; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_22; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_23; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_24; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_25; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_26; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_27; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_28; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_29; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_30; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_31; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_0; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_1; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_2; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_3; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_pc; // @[EXU_AXI.scala 163:27]
  wire [11:0] csr_addr = io_imm[11:0]; // @[EXU_AXI.scala 39:26]
  wire [1:0] _csr_index_T_5 = 12'h300 == csr_addr ? 2'h2 : {{1'd0}, 12'h341 == csr_addr}; // @[Mux.scala 81:58]
  wire  _csr_index_T_6 = 12'h342 == csr_addr; // @[Mux.scala 81:61]
  wire [63:0] _src1_value_T_1 = io_rs1 == 5'h0 ? 64'h0 : Regfile_src1_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] src1_value = io_ctrl_sign_src1_is_pc ? io_pc : _src1_value_T_1; // @[EXU_AXI.scala 49:25]
  wire [63:0] _src2_value_T_1 = io_rs2 == 5'h0 ? 64'h0 : Regfile_src2_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] src2_value = io_ctrl_sign_src2_is_imm ? io_imm : _src2_value_T_1; // @[EXU_AXI.scala 50:25]
  wire [63:0] add_res = src1_value + src2_value; // @[EXU_AXI.scala 51:30]
  wire [63:0] sub_res = src1_value - src2_value; // @[EXU_AXI.scala 52:30]
  wire [63:0] _sra_res_T = io_ctrl_sign_src1_is_pc ? io_pc : _src1_value_T_1; // @[EXU_AXI.scala 53:37]
  wire [63:0] sra_res = $signed(_sra_res_T) >>> src2_value[5:0]; // @[EXU_AXI.scala 53:60]
  wire [63:0] srl_res = src1_value >> src2_value[5:0]; // @[EXU_AXI.scala 54:30]
  wire [126:0] _GEN_1 = {{63'd0}, src1_value}; // @[EXU_AXI.scala 55:30]
  wire [126:0] sll_res = _GEN_1 << src2_value[5:0]; // @[EXU_AXI.scala 55:30]
  wire [31:0] _sraw_res_T_1 = src1_value[31:0]; // @[EXU_AXI.scala 56:43]
  wire [31:0] sraw_res = $signed(_sraw_res_T_1) >>> src2_value[4:0]; // @[EXU_AXI.scala 56:46]
  wire [31:0] srlw_res = src1_value[31:0] >> src2_value[4:0]; // @[EXU_AXI.scala 57:37]
  wire [62:0] _GEN_2 = {{31'd0}, src1_value[31:0]}; // @[EXU_AXI.scala 58:37]
  wire [62:0] sllw_res = _GEN_2 << src2_value[4:0]; // @[EXU_AXI.scala 58:37]
  wire [63:0] or_res = src1_value | src2_value; // @[EXU_AXI.scala 59:29]
  wire [63:0] xor_res = src1_value ^ src2_value; // @[EXU_AXI.scala 60:30]
  wire [63:0] and_res = src1_value & src2_value; // @[EXU_AXI.scala 61:30]
  wire [127:0] _mlu_res_T = src1_value * src2_value; // @[EXU_AXI.scala 62:31]
  wire [63:0] mlu_res = _mlu_res_T[63:0]; // @[EXU_AXI.scala 62:44]
  wire [63:0] _mluw_res_T_2 = src1_value[31:0] * src2_value[31:0]; // @[EXU_AXI.scala 63:38]
  wire [31:0] mluw_res = _mluw_res_T_2[31:0]; // @[EXU_AXI.scala 63:57]
  wire [31:0] _divw_res_T_3 = src2_value[31:0]; // @[EXU_AXI.scala 64:64]
  wire [32:0] _divw_res_T_4 = $signed(_sraw_res_T_1) / $signed(_divw_res_T_3); // @[EXU_AXI.scala 64:45]
  wire [31:0] divw_res = _divw_res_T_4[31:0]; // @[EXU_AXI.scala 64:71]
  wire [31:0] divuw_res = src1_value[31:0] / src2_value[31:0]; // @[EXU_AXI.scala 65:39]
  wire [31:0] remw_res = $signed(_sraw_res_T_1) % $signed(_divw_res_T_3); // @[EXU_AXI.scala 66:71]
  wire [31:0] remuw_res = src1_value[31:0] % src2_value[31:0]; // @[EXU_AXI.scala 67:39]
  wire [63:0] _div_res_T_1 = io_ctrl_sign_src2_is_imm ? io_imm : _src2_value_T_1; // @[EXU_AXI.scala 68:51]
  wire [64:0] div_res = $signed(_sra_res_T) / $signed(_div_res_T_1); // @[EXU_AXI.scala 68:59]
  wire [63:0] divu_res = src1_value / src2_value; // @[EXU_AXI.scala 69:31]
  wire [63:0] rem_res = $signed(_sra_res_T) % $signed(_div_res_T_1); // @[EXU_AXI.scala 70:59]
  wire [63:0] remu_res = src1_value % src2_value; // @[EXU_AXI.scala 71:31]
  wire [63:0] _io_res2rd_T_1 = io_pc + 64'h4; // @[EXU_AXI.scala 76:24]
  wire  _io_res2rd_T_4 = src1_value < src2_value; // @[EXU_AXI.scala 78:34]
  wire  _io_res2rd_T_10 = $signed(_sra_res_T) < $signed(_div_res_T_1); // @[EXU_AXI.scala 80:42]
  wire [31:0] _io_res2rd_T_18 = io_Mem_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_20 = {_io_res2rd_T_18,io_Mem_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_23 = {56'h0,io_Mem_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_26 = {32'h0,io_Mem_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [47:0] _io_res2rd_T_29 = io_Mem_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_31 = {_io_res2rd_T_29,io_Mem_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [55:0] _io_res2rd_T_34 = io_Mem_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_36 = {_io_res2rd_T_34,io_Mem_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_39 = {48'h0,io_Mem_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_42 = add_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_44 = {_io_res2rd_T_42,add_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_52 = sub_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_54 = {_io_res2rd_T_52,sub_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_57 = sllw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_59 = {_io_res2rd_T_57,sllw_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_67 = sraw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _io_res2rd_T_68 = $signed(_sraw_res_T_1) >>> src2_value[4:0]; // @[EXU_AXI.scala 105:56]
  wire [63:0] _io_res2rd_T_69 = {_io_res2rd_T_67,_io_res2rd_T_68}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_72 = srlw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_74 = {_io_res2rd_T_72,srlw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_87 = mluw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_88 = {_io_res2rd_T_87,mluw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_91 = divw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_92 = {_io_res2rd_T_91,divw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_95 = divuw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_96 = {_io_res2rd_T_95,divuw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_99 = remw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_100 = {_io_res2rd_T_99,remw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_103 = remuw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_104 = {_io_res2rd_T_103,remuw_res}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_106 = 32'h1 == io_inst_now ? add_res : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_108 = 32'h3 == io_inst_now ? add_res : _io_res2rd_T_106; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_110 = 32'h4 == io_inst_now ? io_imm : _io_res2rd_T_108; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_112 = 32'h5 == io_inst_now ? _io_res2rd_T_1 : _io_res2rd_T_110; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_114 = 32'h6 == io_inst_now ? _io_res2rd_T_1 : _io_res2rd_T_112; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_116 = 32'h20 == io_inst_now ? {{63'd0}, _io_res2rd_T_4} : _io_res2rd_T_114; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_118 = 32'h1e == io_inst_now ? {{63'd0}, _io_res2rd_T_4} : _io_res2rd_T_116; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_120 = 32'h36 == io_inst_now ? {{63'd0}, _io_res2rd_T_10} : _io_res2rd_T_118; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_122 = 32'h1f == io_inst_now ? {{63'd0}, _io_res2rd_T_10} : _io_res2rd_T_120; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_124 = 32'h21 == io_inst_now ? _io_res2rd_T_20 : _io_res2rd_T_122; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_126 = 32'h22 == io_inst_now ? io_Mem_rdata : _io_res2rd_T_124; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_128 = 32'h23 == io_inst_now ? _io_res2rd_T_23 : _io_res2rd_T_126; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_130 = 32'h3a == io_inst_now ? _io_res2rd_T_26 : _io_res2rd_T_128; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_132 = 32'h24 == io_inst_now ? _io_res2rd_T_31 : _io_res2rd_T_130; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_134 = 32'h3b == io_inst_now ? _io_res2rd_T_36 : _io_res2rd_T_132; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_136 = 32'h25 == io_inst_now ? _io_res2rd_T_39 : _io_res2rd_T_134; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_138 = 32'hc == io_inst_now ? _io_res2rd_T_44 : _io_res2rd_T_136; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_140 = 32'he == io_inst_now ? sub_res : _io_res2rd_T_138; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_142 = 32'h10 == io_inst_now ? _io_res2rd_T_44 : _io_res2rd_T_140; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_144 = 32'hf == io_inst_now ? add_res : _io_res2rd_T_142; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_146 = 32'h15 == io_inst_now ? sra_res : _io_res2rd_T_144; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_148 = 32'hb == io_inst_now ? or_res : _io_res2rd_T_146; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_150 = 32'h2f == io_inst_now ? or_res : _io_res2rd_T_148; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_152 = 32'h2e == io_inst_now ? xor_res : _io_res2rd_T_150; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_154 = 32'ha == io_inst_now ? xor_res : _io_res2rd_T_152; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_156 = 32'h8 == io_inst_now ? and_res : _io_res2rd_T_154; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_158 = 32'h9 == io_inst_now ? and_res : _io_res2rd_T_156; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_160 = 32'hd == io_inst_now ? _io_res2rd_T_54 : _io_res2rd_T_158; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_162 = 32'h16 == io_inst_now ? _io_res2rd_T_59 : _io_res2rd_T_160; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_164 = 32'h17 == io_inst_now ? sll_res : {{63'd0}, _io_res2rd_T_162}; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_166 = 32'h18 == io_inst_now ? {{63'd0}, srl_res} : _io_res2rd_T_164; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_168 = 32'h19 == io_inst_now ? {{63'd0}, _io_res2rd_T_59} : _io_res2rd_T_166; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_170 = 32'h1a == io_inst_now ? {{63'd0}, _io_res2rd_T_69} : _io_res2rd_T_168; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_172 = 32'h1b == io_inst_now ? {{63'd0}, _io_res2rd_T_74} : _io_res2rd_T_170; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_174 = 32'h1c == io_inst_now ? {{63'd0}, _io_res2rd_T_69} : _io_res2rd_T_172; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_176 = 32'h1d == io_inst_now ? {{63'd0}, _io_res2rd_T_74} : _io_res2rd_T_174; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_178 = 32'h11 == io_inst_now ? {{63'd0}, mlu_res} : _io_res2rd_T_176; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_180 = 32'h12 == io_inst_now ? {{63'd0}, _io_res2rd_T_88} : _io_res2rd_T_178; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_182 = 32'h13 == io_inst_now ? {{63'd0}, _io_res2rd_T_92} : _io_res2rd_T_180; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_184 = 32'h30 == io_inst_now ? {{63'd0}, divu_res} : _io_res2rd_T_182; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_186 = 32'h31 == io_inst_now ? {{62'd0}, div_res} : _io_res2rd_T_184; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_188 = 32'h35 == io_inst_now ? {{63'd0}, _io_res2rd_T_96} : _io_res2rd_T_186; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_190 = 32'h14 == io_inst_now ? {{63'd0}, _io_res2rd_T_100} : _io_res2rd_T_188; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_192 = 32'h32 == io_inst_now ? {{63'd0}, _io_res2rd_T_104} : _io_res2rd_T_190; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_194 = 32'h33 == io_inst_now ? {{63'd0}, remu_res} : _io_res2rd_T_192; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_196 = 32'h34 == io_inst_now ? {{63'd0}, rem_res} : _io_res2rd_T_194; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_198 = 32'h37 == io_inst_now ? sll_res : _io_res2rd_T_196; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_200 = 32'h39 == io_inst_now ? {{63'd0}, sra_res} : _io_res2rd_T_198; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_202 = 32'h38 == io_inst_now ? {{63'd0}, srl_res} : _io_res2rd_T_200; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_204 = 32'h3f == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_data} : _io_res2rd_T_202; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_206 = 32'h46 == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_1_data} : _io_res2rd_T_204; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_208 = 32'h47 == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_2_data} : _io_res2rd_T_206; // @[Mux.scala 81:58]
  wire [63:0] reg_value = io_rd == 5'h0 ? 64'h0 : Regfile_reg_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire  _T_6 = io_ctrl_sign_reg_write & io_rd != 5'h0 & (io_inst_valid & ~io_ctrl_sign_Readmem_en |
    io_ctrl_sign_Readmem_en & io_rdata_valid); // @[EXU_AXI.scala 129:63]
  wire [63:0] _csr_wdata_T = src1_value | CSR_Reg_csr_wdata_MPORT_data; // @[EXU_AXI.scala 134:32]
  wire [63:0] _csr_wdata_T_1 = ~CSR_Reg_csr_wdata_MPORT_1_data; // @[EXU_AXI.scala 135:35]
  wire [63:0] _csr_wdata_T_2 = src1_value & _csr_wdata_T_1; // @[EXU_AXI.scala 135:32]
  wire [63:0] _csr_wdata_T_4 = 32'h3f == io_inst_now ? src1_value : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _csr_wdata_T_6 = 32'h46 == io_inst_now ? _csr_wdata_T : _csr_wdata_T_4; // @[Mux.scala 81:58]
  wire [63:0] csr_wdata = 32'h47 == io_inst_now ? _csr_wdata_T_2 : _csr_wdata_T_6; // @[Mux.scala 81:58]
  wire  _T_9 = io_inst_now == 32'h3d & io_inst_valid; // @[EXU_AXI.scala 138:48]
  wire  _T_14 = io_ctrl_sign_csr_write & io_inst_valid; // @[EXU_AXI.scala 141:53]
  wire [63:0] _j_pc_T = add_res & 64'hfffffffffffffffe; // @[EXU_AXI.scala 148:28]
  wire [63:0] _j_pc_T_3 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_data; // @[EXU_AXI.scala 149:39]
  wire [63:0] _j_pc_T_6 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_1_data; // @[EXU_AXI.scala 149:67]
  wire [63:0] _j_pc_T_8 = $signed(_j_pc_T_3) != $signed(_j_pc_T_6) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 149:21]
  wire [63:0] _j_pc_T_11 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_2_data; // @[EXU_AXI.scala 150:39]
  wire [63:0] _j_pc_T_14 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_3_data; // @[EXU_AXI.scala 150:67]
  wire [63:0] _j_pc_T_16 = $signed(_j_pc_T_11) == $signed(_j_pc_T_14) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 150:21]
  wire [63:0] _j_pc_T_19 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_4_data; // @[EXU_AXI.scala 151:39]
  wire [63:0] _j_pc_T_22 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_5_data; // @[EXU_AXI.scala 151:66]
  wire [63:0] _j_pc_T_24 = $signed(_j_pc_T_19) >= $signed(_j_pc_T_22) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 151:21]
  wire [63:0] _j_pc_T_27 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_6_data; // @[EXU_AXI.scala 152:39]
  wire [63:0] _j_pc_T_30 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_7_data; // @[EXU_AXI.scala 152:65]
  wire [63:0] _j_pc_T_32 = $signed(_j_pc_T_27) < $signed(_j_pc_T_30) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 152:21]
  wire [63:0] _j_pc_T_34 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_8_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_36 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_9_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_38 = _j_pc_T_34 < _j_pc_T_36 ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 153:22]
  wire [63:0] _j_pc_T_40 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_10_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_42 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_11_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_44 = _j_pc_T_40 >= _j_pc_T_42 ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 154:22]
  wire [63:0] _j_pc_T_46 = CSR_Reg_j_pc_MPORT_13_data + 64'h4; // @[EXU_AXI.scala 156:33]
  wire [63:0] _j_pc_T_48 = 32'h5 == io_inst_now ? add_res : _io_res2rd_T_1; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_50 = 32'h6 == io_inst_now ? _j_pc_T : _j_pc_T_48; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_52 = 32'h2a == io_inst_now ? _j_pc_T_8 : _j_pc_T_50; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_54 = 32'h29 == io_inst_now ? _j_pc_T_16 : _j_pc_T_52; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_56 = 32'h2b == io_inst_now ? _j_pc_T_24 : _j_pc_T_54; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_58 = 32'h2c == io_inst_now ? _j_pc_T_32 : _j_pc_T_56; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_60 = 32'h2d == io_inst_now ? _j_pc_T_38 : _j_pc_T_58; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_62 = 32'h3c == io_inst_now ? _j_pc_T_44 : _j_pc_T_60; // @[Mux.scala 81:58]
  reg [63:0] pc_next; // @[EXU_AXI.scala 158:26]
  wire [63:0] _mem_wdata_T_1 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_3 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_1_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_6 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_2_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_9 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_3_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_12 = 32'h7 == io_inst_now ? _mem_wdata_T_1 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _mem_wdata_T_14 = 32'h26 == io_inst_now ? {{48'd0}, _mem_wdata_T_3[15:0]} : _mem_wdata_T_12; // @[Mux.scala 81:58]
  wire [63:0] _mem_wdata_T_16 = 32'h28 == io_inst_now ? {{56'd0}, _mem_wdata_T_6[7:0]} : _mem_wdata_T_14; // @[Mux.scala 81:58]
  traceregs reg_trace ( // @[EXU_AXI.scala 163:27]
    .input_reg_0(reg_trace_input_reg_0),
    .input_reg_1(reg_trace_input_reg_1),
    .input_reg_2(reg_trace_input_reg_2),
    .input_reg_3(reg_trace_input_reg_3),
    .input_reg_4(reg_trace_input_reg_4),
    .input_reg_5(reg_trace_input_reg_5),
    .input_reg_6(reg_trace_input_reg_6),
    .input_reg_7(reg_trace_input_reg_7),
    .input_reg_8(reg_trace_input_reg_8),
    .input_reg_9(reg_trace_input_reg_9),
    .input_reg_10(reg_trace_input_reg_10),
    .input_reg_11(reg_trace_input_reg_11),
    .input_reg_12(reg_trace_input_reg_12),
    .input_reg_13(reg_trace_input_reg_13),
    .input_reg_14(reg_trace_input_reg_14),
    .input_reg_15(reg_trace_input_reg_15),
    .input_reg_16(reg_trace_input_reg_16),
    .input_reg_17(reg_trace_input_reg_17),
    .input_reg_18(reg_trace_input_reg_18),
    .input_reg_19(reg_trace_input_reg_19),
    .input_reg_20(reg_trace_input_reg_20),
    .input_reg_21(reg_trace_input_reg_21),
    .input_reg_22(reg_trace_input_reg_22),
    .input_reg_23(reg_trace_input_reg_23),
    .input_reg_24(reg_trace_input_reg_24),
    .input_reg_25(reg_trace_input_reg_25),
    .input_reg_26(reg_trace_input_reg_26),
    .input_reg_27(reg_trace_input_reg_27),
    .input_reg_28(reg_trace_input_reg_28),
    .input_reg_29(reg_trace_input_reg_29),
    .input_reg_30(reg_trace_input_reg_30),
    .input_reg_31(reg_trace_input_reg_31),
    .csr_reg_0(reg_trace_csr_reg_0),
    .csr_reg_1(reg_trace_csr_reg_1),
    .csr_reg_2(reg_trace_csr_reg_2),
    .csr_reg_3(reg_trace_csr_reg_3),
    .pc(reg_trace_pc)
  );
  assign Regfile_src1_value_MPORT_en = 1'h1;
  assign Regfile_src1_value_MPORT_addr = io_rs1;
  assign Regfile_src1_value_MPORT_data = Regfile[Regfile_src1_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_src2_value_MPORT_en = 1'h1;
  assign Regfile_src2_value_MPORT_addr = io_rs2;
  assign Regfile_src2_value_MPORT_data = Regfile[Regfile_src2_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_value_MPORT_en = 1'h1;
  assign Regfile_reg_value_MPORT_addr = io_rd;
  assign Regfile_reg_value_MPORT_data = Regfile[Regfile_reg_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_MPORT_4_en = 1'h1;
  assign Regfile_MPORT_4_addr = 5'h11;
  assign Regfile_MPORT_4_data = Regfile[Regfile_MPORT_4_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_en = 1'h1;
  assign Regfile_j_pc_MPORT_addr = io_rs1;
  assign Regfile_j_pc_MPORT_data = Regfile[Regfile_j_pc_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_1_en = 1'h1;
  assign Regfile_j_pc_MPORT_1_addr = io_rs2;
  assign Regfile_j_pc_MPORT_1_data = Regfile[Regfile_j_pc_MPORT_1_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_2_en = 1'h1;
  assign Regfile_j_pc_MPORT_2_addr = io_rs1;
  assign Regfile_j_pc_MPORT_2_data = Regfile[Regfile_j_pc_MPORT_2_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_3_en = 1'h1;
  assign Regfile_j_pc_MPORT_3_addr = io_rs2;
  assign Regfile_j_pc_MPORT_3_data = Regfile[Regfile_j_pc_MPORT_3_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_4_en = 1'h1;
  assign Regfile_j_pc_MPORT_4_addr = io_rs1;
  assign Regfile_j_pc_MPORT_4_data = Regfile[Regfile_j_pc_MPORT_4_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_5_en = 1'h1;
  assign Regfile_j_pc_MPORT_5_addr = io_rs2;
  assign Regfile_j_pc_MPORT_5_data = Regfile[Regfile_j_pc_MPORT_5_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_6_en = 1'h1;
  assign Regfile_j_pc_MPORT_6_addr = io_rs1;
  assign Regfile_j_pc_MPORT_6_data = Regfile[Regfile_j_pc_MPORT_6_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_7_en = 1'h1;
  assign Regfile_j_pc_MPORT_7_addr = io_rs2;
  assign Regfile_j_pc_MPORT_7_data = Regfile[Regfile_j_pc_MPORT_7_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_8_en = 1'h1;
  assign Regfile_j_pc_MPORT_8_addr = io_rs1;
  assign Regfile_j_pc_MPORT_8_data = Regfile[Regfile_j_pc_MPORT_8_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_9_en = 1'h1;
  assign Regfile_j_pc_MPORT_9_addr = io_rs2;
  assign Regfile_j_pc_MPORT_9_data = Regfile[Regfile_j_pc_MPORT_9_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_10_en = 1'h1;
  assign Regfile_j_pc_MPORT_10_addr = io_rs1;
  assign Regfile_j_pc_MPORT_10_data = Regfile[Regfile_j_pc_MPORT_10_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_11_en = 1'h1;
  assign Regfile_j_pc_MPORT_11_addr = io_rs2;
  assign Regfile_j_pc_MPORT_11_data = Regfile[Regfile_j_pc_MPORT_11_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_0_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_0_MPORT_addr = 5'h0;
  assign Regfile_reg_trace_io_input_reg_0_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_0_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_1_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_1_MPORT_addr = 5'h1;
  assign Regfile_reg_trace_io_input_reg_1_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_1_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_2_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_2_MPORT_addr = 5'h2;
  assign Regfile_reg_trace_io_input_reg_2_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_2_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_3_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_3_MPORT_addr = 5'h3;
  assign Regfile_reg_trace_io_input_reg_3_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_3_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_4_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_4_MPORT_addr = 5'h4;
  assign Regfile_reg_trace_io_input_reg_4_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_4_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_5_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_5_MPORT_addr = 5'h5;
  assign Regfile_reg_trace_io_input_reg_5_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_5_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_6_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_6_MPORT_addr = 5'h6;
  assign Regfile_reg_trace_io_input_reg_6_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_6_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_7_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_7_MPORT_addr = 5'h7;
  assign Regfile_reg_trace_io_input_reg_7_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_7_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_8_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_8_MPORT_addr = 5'h8;
  assign Regfile_reg_trace_io_input_reg_8_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_8_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_9_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_9_MPORT_addr = 5'h9;
  assign Regfile_reg_trace_io_input_reg_9_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_9_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_10_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_10_MPORT_addr = 5'ha;
  assign Regfile_reg_trace_io_input_reg_10_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_10_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_11_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_11_MPORT_addr = 5'hb;
  assign Regfile_reg_trace_io_input_reg_11_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_11_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_12_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_12_MPORT_addr = 5'hc;
  assign Regfile_reg_trace_io_input_reg_12_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_12_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_13_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_13_MPORT_addr = 5'hd;
  assign Regfile_reg_trace_io_input_reg_13_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_13_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_14_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_14_MPORT_addr = 5'he;
  assign Regfile_reg_trace_io_input_reg_14_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_14_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_15_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_15_MPORT_addr = 5'hf;
  assign Regfile_reg_trace_io_input_reg_15_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_15_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_16_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_16_MPORT_addr = 5'h10;
  assign Regfile_reg_trace_io_input_reg_16_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_16_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_17_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_17_MPORT_addr = 5'h11;
  assign Regfile_reg_trace_io_input_reg_17_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_17_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_18_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_18_MPORT_addr = 5'h12;
  assign Regfile_reg_trace_io_input_reg_18_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_18_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_19_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_19_MPORT_addr = 5'h13;
  assign Regfile_reg_trace_io_input_reg_19_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_19_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_20_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_20_MPORT_addr = 5'h14;
  assign Regfile_reg_trace_io_input_reg_20_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_20_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_21_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_21_MPORT_addr = 5'h15;
  assign Regfile_reg_trace_io_input_reg_21_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_21_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_22_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_22_MPORT_addr = 5'h16;
  assign Regfile_reg_trace_io_input_reg_22_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_22_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_23_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_23_MPORT_addr = 5'h17;
  assign Regfile_reg_trace_io_input_reg_23_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_23_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_24_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_24_MPORT_addr = 5'h18;
  assign Regfile_reg_trace_io_input_reg_24_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_24_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_25_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_25_MPORT_addr = 5'h19;
  assign Regfile_reg_trace_io_input_reg_25_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_25_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_26_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_26_MPORT_addr = 5'h1a;
  assign Regfile_reg_trace_io_input_reg_26_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_26_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_27_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_27_MPORT_addr = 5'h1b;
  assign Regfile_reg_trace_io_input_reg_27_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_27_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_28_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_28_MPORT_addr = 5'h1c;
  assign Regfile_reg_trace_io_input_reg_28_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_28_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_29_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_29_MPORT_addr = 5'h1d;
  assign Regfile_reg_trace_io_input_reg_29_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_29_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_30_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_30_MPORT_addr = 5'h1e;
  assign Regfile_reg_trace_io_input_reg_30_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_30_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_31_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_31_MPORT_addr = 5'h1f;
  assign Regfile_reg_trace_io_input_reg_31_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_31_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_data = Regfile[Regfile_mem_wdata_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_1_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_1_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_1_data = Regfile[Regfile_mem_wdata_MPORT_1_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_2_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_2_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_2_data = Regfile[Regfile_mem_wdata_MPORT_2_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_3_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_3_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_3_data = Regfile[Regfile_mem_wdata_MPORT_3_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_MPORT_data = _T_6 ? io_res2rd : reg_value;
  assign Regfile_MPORT_addr = io_rd;
  assign Regfile_MPORT_mask = 1'h1;
  assign Regfile_MPORT_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_io_res2rd_MPORT_1_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_1_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_1_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_1_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_io_res2rd_MPORT_2_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_2_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_2_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_2_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_csr_wdata_MPORT_en = 1'h1;
  assign CSR_Reg_csr_wdata_MPORT_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_csr_wdata_MPORT_data = CSR_Reg[CSR_Reg_csr_wdata_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_csr_wdata_MPORT_1_en = 1'h1;
  assign CSR_Reg_csr_wdata_MPORT_1_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_csr_wdata_MPORT_1_data = CSR_Reg[CSR_Reg_csr_wdata_MPORT_1_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_2_en = 1'h1;
  assign CSR_Reg_MPORT_2_addr = 2'h1;
  assign CSR_Reg_MPORT_2_data = CSR_Reg[CSR_Reg_MPORT_2_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_5_en = 1'h1;
  assign CSR_Reg_MPORT_5_addr = 2'h3;
  assign CSR_Reg_MPORT_5_data = CSR_Reg[CSR_Reg_MPORT_5_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_7_en = 1'h1;
  assign CSR_Reg_MPORT_7_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_MPORT_7_data = CSR_Reg[CSR_Reg_MPORT_7_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_j_pc_MPORT_12_en = 1'h1;
  assign CSR_Reg_j_pc_MPORT_12_addr = 2'h0;
  assign CSR_Reg_j_pc_MPORT_12_data = CSR_Reg[CSR_Reg_j_pc_MPORT_12_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_j_pc_MPORT_13_en = 1'h1;
  assign CSR_Reg_j_pc_MPORT_13_addr = 2'h1;
  assign CSR_Reg_j_pc_MPORT_13_data = CSR_Reg[CSR_Reg_j_pc_MPORT_13_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr = 2'h0;
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr = 2'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr = 2'h2;
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_1_data = _T_9 ? io_pc : CSR_Reg_MPORT_2_data;
  assign CSR_Reg_MPORT_1_addr = 2'h1;
  assign CSR_Reg_MPORT_1_mask = 1'h1;
  assign CSR_Reg_MPORT_1_en = 1'h1;
  assign CSR_Reg_MPORT_3_data = _T_9 ? Regfile_MPORT_4_data : CSR_Reg_MPORT_5_data;
  assign CSR_Reg_MPORT_3_addr = 2'h3;
  assign CSR_Reg_MPORT_3_mask = 1'h1;
  assign CSR_Reg_MPORT_3_en = 1'h1;
  assign CSR_Reg_MPORT_6_data = _T_14 ? csr_wdata : CSR_Reg_MPORT_7_data;
  assign CSR_Reg_MPORT_6_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_MPORT_6_mask = 1'h1;
  assign CSR_Reg_MPORT_6_en = 1'h1;
  assign io_pc_next = pc_next; // @[EXU_AXI.scala 162:16]
  assign io_res2rd = _io_res2rd_T_208[63:0]; // @[EXU_AXI.scala 72:15]
  assign io_inst_store = io_ctrl_sign_Writemem_en; // @[EXU_AXI.scala 188:19]
  assign io_inst_load = io_ctrl_sign_Readmem_en; // @[EXU_AXI.scala 189:18]
  assign io_Mem_addr = add_res[31:0]; // @[EXU_AXI.scala 190:17]
  assign io_Mem_wdata = 32'h27 == io_inst_now ? {{32'd0}, _mem_wdata_T_9[31:0]} : _mem_wdata_T_16; // @[Mux.scala 81:58]
  assign io_Mem_wstrb = io_ctrl_sign_Wmask; // @[EXU_AXI.scala 192:18]
  assign reg_trace_input_reg_0 = Regfile_reg_trace_io_input_reg_0_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_1 = Regfile_reg_trace_io_input_reg_1_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_2 = Regfile_reg_trace_io_input_reg_2_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_3 = Regfile_reg_trace_io_input_reg_3_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_4 = Regfile_reg_trace_io_input_reg_4_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_5 = Regfile_reg_trace_io_input_reg_5_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_6 = Regfile_reg_trace_io_input_reg_6_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_7 = Regfile_reg_trace_io_input_reg_7_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_8 = Regfile_reg_trace_io_input_reg_8_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_9 = Regfile_reg_trace_io_input_reg_9_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_10 = Regfile_reg_trace_io_input_reg_10_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_11 = Regfile_reg_trace_io_input_reg_11_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_12 = Regfile_reg_trace_io_input_reg_12_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_13 = Regfile_reg_trace_io_input_reg_13_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_14 = Regfile_reg_trace_io_input_reg_14_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_15 = Regfile_reg_trace_io_input_reg_15_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_16 = Regfile_reg_trace_io_input_reg_16_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_17 = Regfile_reg_trace_io_input_reg_17_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_18 = Regfile_reg_trace_io_input_reg_18_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_19 = Regfile_reg_trace_io_input_reg_19_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_20 = Regfile_reg_trace_io_input_reg_20_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_21 = Regfile_reg_trace_io_input_reg_21_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_22 = Regfile_reg_trace_io_input_reg_22_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_23 = Regfile_reg_trace_io_input_reg_23_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_24 = Regfile_reg_trace_io_input_reg_24_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_25 = Regfile_reg_trace_io_input_reg_25_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_26 = Regfile_reg_trace_io_input_reg_26_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_27 = Regfile_reg_trace_io_input_reg_27_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_28 = Regfile_reg_trace_io_input_reg_28_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_29 = Regfile_reg_trace_io_input_reg_29_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_30 = Regfile_reg_trace_io_input_reg_30_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_31 = Regfile_reg_trace_io_input_reg_31_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_csr_reg_0 = CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_1 = CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_2 = CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_3 = 64'h0; // @[EXU_AXI.scala 167:{36,36}]
  assign reg_trace_pc = io_pc; // @[EXU_AXI.scala 166:21]
  always @(posedge clock) begin
    if (Regfile_MPORT_en & Regfile_MPORT_mask) begin
      Regfile[Regfile_MPORT_addr] <= Regfile_MPORT_data; // @[EXU_AXI.scala 37:22]
    end
    if (CSR_Reg_MPORT_1_en & CSR_Reg_MPORT_1_mask) begin
      CSR_Reg[CSR_Reg_MPORT_1_addr] <= CSR_Reg_MPORT_1_data; // @[EXU_AXI.scala 38:22]
    end
    if (CSR_Reg_MPORT_3_en & CSR_Reg_MPORT_3_mask) begin
      CSR_Reg[CSR_Reg_MPORT_3_addr] <= CSR_Reg_MPORT_3_data; // @[EXU_AXI.scala 38:22]
    end
    if (CSR_Reg_MPORT_6_en & CSR_Reg_MPORT_6_mask) begin
      CSR_Reg[CSR_Reg_MPORT_6_addr] <= CSR_Reg_MPORT_6_data; // @[EXU_AXI.scala 38:22]
    end
    if (reset) begin // @[EXU_AXI.scala 158:26]
      pc_next <= 64'h0; // @[EXU_AXI.scala 158:26]
    end else if (io_inst_valid) begin // @[EXU_AXI.scala 159:24]
      if (32'h3e == io_inst_now) begin // @[Mux.scala 81:58]
        pc_next <= _j_pc_T_46;
      end else if (32'h3d == io_inst_now) begin // @[Mux.scala 81:58]
        pc_next <= CSR_Reg_j_pc_MPORT_12_data;
      end else begin
        pc_next <= _j_pc_T_62;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    Regfile[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    CSR_Reg[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  pc_next = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top(
  input         clock,
  input         reset,
  output [31:0] io_inst,
  output [63:0] io_pc,
  output [63:0] io_pc_next,
  output [63:0] io_outval,
  output        io_step
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  axi_clock; // @[top.scala 18:21]
  wire  axi_reset; // @[top.scala 18:21]
  wire [31:0] axi_io_axi_in_araddr; // @[top.scala 18:21]
  wire  axi_io_axi_in_arvalid; // @[top.scala 18:21]
  wire  axi_io_axi_in_rready; // @[top.scala 18:21]
  wire [31:0] axi_io_axi_in_awaddr; // @[top.scala 18:21]
  wire  axi_io_axi_in_awvalid; // @[top.scala 18:21]
  wire [31:0] axi_io_axi_in_wdata; // @[top.scala 18:21]
  wire [7:0] axi_io_axi_in_wstrb; // @[top.scala 18:21]
  wire  axi_io_axi_in_wvalid; // @[top.scala 18:21]
  wire  axi_io_axi_in_bready; // @[top.scala 18:21]
  wire  axi_io_axi_out_arready; // @[top.scala 18:21]
  wire [63:0] axi_io_axi_out_rdata; // @[top.scala 18:21]
  wire  axi_io_axi_out_rvalid; // @[top.scala 18:21]
  wire  axi_io_axi_out_awready; // @[top.scala 18:21]
  wire  axi_io_axi_out_wready; // @[top.scala 18:21]
  wire  axi_io_axi_out_bvalid; // @[top.scala 18:21]
  wire  lsu_step_clock; // @[top.scala 19:26]
  wire  lsu_step_reset; // @[top.scala 19:26]
  wire  lsu_step_io_inst_store; // @[top.scala 19:26]
  wire  lsu_step_io_inst_load; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_mem_addr; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_mem_wdata; // @[top.scala 19:26]
  wire [7:0] lsu_step_io_mem_wstrb; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_mem_rdata; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_arready; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_axi_in_rdata; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_rvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_awready; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_wready; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_bvalid; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_axi_out_araddr; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_arvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_rready; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_axi_out_awaddr; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_awvalid; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_axi_out_wdata; // @[top.scala 19:26]
  wire [7:0] lsu_step_io_axi_out_wstrb; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_wvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_bready; // @[top.scala 19:26]
  wire  arbiter_clock; // @[top.scala 20:25]
  wire  arbiter_reset; // @[top.scala 20:25]
  wire [31:0] arbiter_io_ifu_axi_in_araddr; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_in_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_in_rready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_ifu_axi_out_rdata; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_out_rvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_lsu_axi_in_araddr; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_rready; // @[top.scala 20:25]
  wire [31:0] arbiter_io_lsu_axi_in_awaddr; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_awvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_lsu_axi_in_wdata; // @[top.scala 20:25]
  wire [7:0] arbiter_io_lsu_axi_in_wstrb; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_wvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_bready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_arready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_lsu_axi_out_rdata; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_rvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_awready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_wready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_bvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_arready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_axi_in_rdata; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_rvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_awready; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_wready; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_bvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_axi_out_araddr; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_rready; // @[top.scala 20:25]
  wire [31:0] arbiter_io_axi_out_awaddr; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_awvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_axi_out_wdata; // @[top.scala 20:25]
  wire [7:0] arbiter_io_axi_out_wstrb; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_wvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_bready; // @[top.scala 20:25]
  wire  ifu_step_clock; // @[top.scala 21:26]
  wire  ifu_step_reset; // @[top.scala 21:26]
  wire [63:0] ifu_step_io_pc; // @[top.scala 21:26]
  wire  ifu_step_io_pc_valid; // @[top.scala 21:26]
  wire  ifu_step_io_inst_valid; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_inst; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_inst_reg; // @[top.scala 21:26]
  wire [63:0] ifu_step_io_axi_in_rdata; // @[top.scala 21:26]
  wire  ifu_step_io_axi_in_rvalid; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_axi_out_araddr; // @[top.scala 21:26]
  wire  ifu_step_io_axi_out_arvalid; // @[top.scala 21:26]
  wire  ifu_step_io_axi_out_rready; // @[top.scala 21:26]
  wire  i_cache_clock; // @[top.scala 22:25]
  wire  i_cache_reset; // @[top.scala 22:25]
  wire [31:0] i_cache_io_from_ifu_araddr; // @[top.scala 22:25]
  wire  i_cache_io_from_ifu_arvalid; // @[top.scala 22:25]
  wire  i_cache_io_from_ifu_rready; // @[top.scala 22:25]
  wire [63:0] i_cache_io_to_ifu_rdata; // @[top.scala 22:25]
  wire  i_cache_io_to_ifu_rvalid; // @[top.scala 22:25]
  wire [31:0] i_cache_io_to_axi_araddr; // @[top.scala 22:25]
  wire  i_cache_io_to_axi_arvalid; // @[top.scala 22:25]
  wire  i_cache_io_to_axi_rready; // @[top.scala 22:25]
  wire [63:0] i_cache_io_from_axi_rdata; // @[top.scala 22:25]
  wire  i_cache_io_from_axi_rvalid; // @[top.scala 22:25]
  wire  d_cache_clock; // @[top.scala 23:25]
  wire  d_cache_reset; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_araddr; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_arvalid; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_rready; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_awaddr; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_awvalid; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_wdata; // @[top.scala 23:25]
  wire [7:0] d_cache_io_from_lsu_wstrb; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_wvalid; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_bready; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_arready; // @[top.scala 23:25]
  wire [63:0] d_cache_io_to_lsu_rdata; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_rvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_awready; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_wready; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_bvalid; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_araddr; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_arvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_rready; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_awaddr; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_awvalid; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_wdata; // @[top.scala 23:25]
  wire [7:0] d_cache_io_to_axi_wstrb; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_wvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_bready; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_arready; // @[top.scala 23:25]
  wire [63:0] d_cache_io_from_axi_rdata; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_rvalid; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_awready; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_wready; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_bvalid; // @[top.scala 23:25]
  wire [31:0] idu_step_io_inst; // @[top.scala 46:26]
  wire [31:0] idu_step_io_inst_now; // @[top.scala 46:26]
  wire [4:0] idu_step_io_rs1; // @[top.scala 46:26]
  wire [4:0] idu_step_io_rs2; // @[top.scala 46:26]
  wire [4:0] idu_step_io_rd; // @[top.scala 46:26]
  wire [63:0] idu_step_io_imm; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_reg_write; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_csr_write; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_Writemem_en; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_Readmem_en; // @[top.scala 46:26]
  wire [7:0] idu_step_io_ctrl_sign_Wmask; // @[top.scala 46:26]
  wire  exu_step_clock; // @[top.scala 51:26]
  wire  exu_step_reset; // @[top.scala 51:26]
  wire [63:0] exu_step_io_pc; // @[top.scala 51:26]
  wire [63:0] exu_step_io_pc_next; // @[top.scala 51:26]
  wire [31:0] exu_step_io_inst_now; // @[top.scala 51:26]
  wire [4:0] exu_step_io_rs1; // @[top.scala 51:26]
  wire [4:0] exu_step_io_rs2; // @[top.scala 51:26]
  wire [4:0] exu_step_io_rd; // @[top.scala 51:26]
  wire [63:0] exu_step_io_imm; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_reg_write; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_csr_write; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_Writemem_en; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_Readmem_en; // @[top.scala 51:26]
  wire [7:0] exu_step_io_ctrl_sign_Wmask; // @[top.scala 51:26]
  wire [63:0] exu_step_io_res2rd; // @[top.scala 51:26]
  wire  exu_step_io_inst_valid; // @[top.scala 51:26]
  wire  exu_step_io_inst_store; // @[top.scala 51:26]
  wire  exu_step_io_inst_load; // @[top.scala 51:26]
  wire [31:0] exu_step_io_Mem_addr; // @[top.scala 51:26]
  wire [63:0] exu_step_io_Mem_rdata; // @[top.scala 51:26]
  wire [63:0] exu_step_io_Mem_wdata; // @[top.scala 51:26]
  wire [7:0] exu_step_io_Mem_wstrb; // @[top.scala 51:26]
  wire  exu_step_io_rdata_valid; // @[top.scala 51:26]
  wire [31:0] dpi_flag; // @[top.scala 73:21]
  wire [31:0] dpi_ecall_flag; // @[top.scala 73:21]
  reg [63:0] pc_now; // @[top.scala 15:25]
  reg  execute_end; // @[top.scala 17:30]
  reg  pc_valid; // @[top.scala 87:27]
  reg  diff_step; // @[top.scala 90:28]
  AXI axi ( // @[top.scala 18:21]
    .clock(axi_clock),
    .reset(axi_reset),
    .io_axi_in_araddr(axi_io_axi_in_araddr),
    .io_axi_in_arvalid(axi_io_axi_in_arvalid),
    .io_axi_in_rready(axi_io_axi_in_rready),
    .io_axi_in_awaddr(axi_io_axi_in_awaddr),
    .io_axi_in_awvalid(axi_io_axi_in_awvalid),
    .io_axi_in_wdata(axi_io_axi_in_wdata),
    .io_axi_in_wstrb(axi_io_axi_in_wstrb),
    .io_axi_in_wvalid(axi_io_axi_in_wvalid),
    .io_axi_in_bready(axi_io_axi_in_bready),
    .io_axi_out_arready(axi_io_axi_out_arready),
    .io_axi_out_rdata(axi_io_axi_out_rdata),
    .io_axi_out_rvalid(axi_io_axi_out_rvalid),
    .io_axi_out_awready(axi_io_axi_out_awready),
    .io_axi_out_wready(axi_io_axi_out_wready),
    .io_axi_out_bvalid(axi_io_axi_out_bvalid)
  );
  LSU lsu_step ( // @[top.scala 19:26]
    .clock(lsu_step_clock),
    .reset(lsu_step_reset),
    .io_inst_store(lsu_step_io_inst_store),
    .io_inst_load(lsu_step_io_inst_load),
    .io_mem_addr(lsu_step_io_mem_addr),
    .io_mem_wdata(lsu_step_io_mem_wdata),
    .io_mem_wstrb(lsu_step_io_mem_wstrb),
    .io_mem_rdata(lsu_step_io_mem_rdata),
    .io_axi_in_arready(lsu_step_io_axi_in_arready),
    .io_axi_in_rdata(lsu_step_io_axi_in_rdata),
    .io_axi_in_rvalid(lsu_step_io_axi_in_rvalid),
    .io_axi_in_awready(lsu_step_io_axi_in_awready),
    .io_axi_in_wready(lsu_step_io_axi_in_wready),
    .io_axi_in_bvalid(lsu_step_io_axi_in_bvalid),
    .io_axi_out_araddr(lsu_step_io_axi_out_araddr),
    .io_axi_out_arvalid(lsu_step_io_axi_out_arvalid),
    .io_axi_out_rready(lsu_step_io_axi_out_rready),
    .io_axi_out_awaddr(lsu_step_io_axi_out_awaddr),
    .io_axi_out_awvalid(lsu_step_io_axi_out_awvalid),
    .io_axi_out_wdata(lsu_step_io_axi_out_wdata),
    .io_axi_out_wstrb(lsu_step_io_axi_out_wstrb),
    .io_axi_out_wvalid(lsu_step_io_axi_out_wvalid),
    .io_axi_out_bready(lsu_step_io_axi_out_bready)
  );
  AXI_ARBITER arbiter ( // @[top.scala 20:25]
    .clock(arbiter_clock),
    .reset(arbiter_reset),
    .io_ifu_axi_in_araddr(arbiter_io_ifu_axi_in_araddr),
    .io_ifu_axi_in_arvalid(arbiter_io_ifu_axi_in_arvalid),
    .io_ifu_axi_in_rready(arbiter_io_ifu_axi_in_rready),
    .io_ifu_axi_out_rdata(arbiter_io_ifu_axi_out_rdata),
    .io_ifu_axi_out_rvalid(arbiter_io_ifu_axi_out_rvalid),
    .io_lsu_axi_in_araddr(arbiter_io_lsu_axi_in_araddr),
    .io_lsu_axi_in_arvalid(arbiter_io_lsu_axi_in_arvalid),
    .io_lsu_axi_in_rready(arbiter_io_lsu_axi_in_rready),
    .io_lsu_axi_in_awaddr(arbiter_io_lsu_axi_in_awaddr),
    .io_lsu_axi_in_awvalid(arbiter_io_lsu_axi_in_awvalid),
    .io_lsu_axi_in_wdata(arbiter_io_lsu_axi_in_wdata),
    .io_lsu_axi_in_wstrb(arbiter_io_lsu_axi_in_wstrb),
    .io_lsu_axi_in_wvalid(arbiter_io_lsu_axi_in_wvalid),
    .io_lsu_axi_in_bready(arbiter_io_lsu_axi_in_bready),
    .io_lsu_axi_out_arready(arbiter_io_lsu_axi_out_arready),
    .io_lsu_axi_out_rdata(arbiter_io_lsu_axi_out_rdata),
    .io_lsu_axi_out_rvalid(arbiter_io_lsu_axi_out_rvalid),
    .io_lsu_axi_out_awready(arbiter_io_lsu_axi_out_awready),
    .io_lsu_axi_out_wready(arbiter_io_lsu_axi_out_wready),
    .io_lsu_axi_out_bvalid(arbiter_io_lsu_axi_out_bvalid),
    .io_axi_in_arready(arbiter_io_axi_in_arready),
    .io_axi_in_rdata(arbiter_io_axi_in_rdata),
    .io_axi_in_rvalid(arbiter_io_axi_in_rvalid),
    .io_axi_in_awready(arbiter_io_axi_in_awready),
    .io_axi_in_wready(arbiter_io_axi_in_wready),
    .io_axi_in_bvalid(arbiter_io_axi_in_bvalid),
    .io_axi_out_araddr(arbiter_io_axi_out_araddr),
    .io_axi_out_arvalid(arbiter_io_axi_out_arvalid),
    .io_axi_out_rready(arbiter_io_axi_out_rready),
    .io_axi_out_awaddr(arbiter_io_axi_out_awaddr),
    .io_axi_out_awvalid(arbiter_io_axi_out_awvalid),
    .io_axi_out_wdata(arbiter_io_axi_out_wdata),
    .io_axi_out_wstrb(arbiter_io_axi_out_wstrb),
    .io_axi_out_wvalid(arbiter_io_axi_out_wvalid),
    .io_axi_out_bready(arbiter_io_axi_out_bready)
  );
  IFU_AXI ifu_step ( // @[top.scala 21:26]
    .clock(ifu_step_clock),
    .reset(ifu_step_reset),
    .io_pc(ifu_step_io_pc),
    .io_pc_valid(ifu_step_io_pc_valid),
    .io_inst_valid(ifu_step_io_inst_valid),
    .io_inst(ifu_step_io_inst),
    .io_inst_reg(ifu_step_io_inst_reg),
    .io_axi_in_rdata(ifu_step_io_axi_in_rdata),
    .io_axi_in_rvalid(ifu_step_io_axi_in_rvalid),
    .io_axi_out_araddr(ifu_step_io_axi_out_araddr),
    .io_axi_out_arvalid(ifu_step_io_axi_out_arvalid),
    .io_axi_out_rready(ifu_step_io_axi_out_rready)
  );
  I_CACHE i_cache ( // @[top.scala 22:25]
    .clock(i_cache_clock),
    .reset(i_cache_reset),
    .io_from_ifu_araddr(i_cache_io_from_ifu_araddr),
    .io_from_ifu_arvalid(i_cache_io_from_ifu_arvalid),
    .io_from_ifu_rready(i_cache_io_from_ifu_rready),
    .io_to_ifu_rdata(i_cache_io_to_ifu_rdata),
    .io_to_ifu_rvalid(i_cache_io_to_ifu_rvalid),
    .io_to_axi_araddr(i_cache_io_to_axi_araddr),
    .io_to_axi_arvalid(i_cache_io_to_axi_arvalid),
    .io_to_axi_rready(i_cache_io_to_axi_rready),
    .io_from_axi_rdata(i_cache_io_from_axi_rdata),
    .io_from_axi_rvalid(i_cache_io_from_axi_rvalid)
  );
  D_CACHE d_cache ( // @[top.scala 23:25]
    .clock(d_cache_clock),
    .reset(d_cache_reset),
    .io_from_lsu_araddr(d_cache_io_from_lsu_araddr),
    .io_from_lsu_arvalid(d_cache_io_from_lsu_arvalid),
    .io_from_lsu_rready(d_cache_io_from_lsu_rready),
    .io_from_lsu_awaddr(d_cache_io_from_lsu_awaddr),
    .io_from_lsu_awvalid(d_cache_io_from_lsu_awvalid),
    .io_from_lsu_wdata(d_cache_io_from_lsu_wdata),
    .io_from_lsu_wstrb(d_cache_io_from_lsu_wstrb),
    .io_from_lsu_wvalid(d_cache_io_from_lsu_wvalid),
    .io_from_lsu_bready(d_cache_io_from_lsu_bready),
    .io_to_lsu_arready(d_cache_io_to_lsu_arready),
    .io_to_lsu_rdata(d_cache_io_to_lsu_rdata),
    .io_to_lsu_rvalid(d_cache_io_to_lsu_rvalid),
    .io_to_lsu_awready(d_cache_io_to_lsu_awready),
    .io_to_lsu_wready(d_cache_io_to_lsu_wready),
    .io_to_lsu_bvalid(d_cache_io_to_lsu_bvalid),
    .io_to_axi_araddr(d_cache_io_to_axi_araddr),
    .io_to_axi_arvalid(d_cache_io_to_axi_arvalid),
    .io_to_axi_rready(d_cache_io_to_axi_rready),
    .io_to_axi_awaddr(d_cache_io_to_axi_awaddr),
    .io_to_axi_awvalid(d_cache_io_to_axi_awvalid),
    .io_to_axi_wdata(d_cache_io_to_axi_wdata),
    .io_to_axi_wstrb(d_cache_io_to_axi_wstrb),
    .io_to_axi_wvalid(d_cache_io_to_axi_wvalid),
    .io_to_axi_bready(d_cache_io_to_axi_bready),
    .io_from_axi_arready(d_cache_io_from_axi_arready),
    .io_from_axi_rdata(d_cache_io_from_axi_rdata),
    .io_from_axi_rvalid(d_cache_io_from_axi_rvalid),
    .io_from_axi_awready(d_cache_io_from_axi_awready),
    .io_from_axi_wready(d_cache_io_from_axi_wready),
    .io_from_axi_bvalid(d_cache_io_from_axi_bvalid)
  );
  IDU idu_step ( // @[top.scala 46:26]
    .io_inst(idu_step_io_inst),
    .io_inst_now(idu_step_io_inst_now),
    .io_rs1(idu_step_io_rs1),
    .io_rs2(idu_step_io_rs2),
    .io_rd(idu_step_io_rd),
    .io_imm(idu_step_io_imm),
    .io_ctrl_sign_reg_write(idu_step_io_ctrl_sign_reg_write),
    .io_ctrl_sign_csr_write(idu_step_io_ctrl_sign_csr_write),
    .io_ctrl_sign_src2_is_imm(idu_step_io_ctrl_sign_src2_is_imm),
    .io_ctrl_sign_src1_is_pc(idu_step_io_ctrl_sign_src1_is_pc),
    .io_ctrl_sign_Writemem_en(idu_step_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(idu_step_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(idu_step_io_ctrl_sign_Wmask)
  );
  EXU_AXI exu_step ( // @[top.scala 51:26]
    .clock(exu_step_clock),
    .reset(exu_step_reset),
    .io_pc(exu_step_io_pc),
    .io_pc_next(exu_step_io_pc_next),
    .io_inst_now(exu_step_io_inst_now),
    .io_rs1(exu_step_io_rs1),
    .io_rs2(exu_step_io_rs2),
    .io_rd(exu_step_io_rd),
    .io_imm(exu_step_io_imm),
    .io_ctrl_sign_reg_write(exu_step_io_ctrl_sign_reg_write),
    .io_ctrl_sign_csr_write(exu_step_io_ctrl_sign_csr_write),
    .io_ctrl_sign_src2_is_imm(exu_step_io_ctrl_sign_src2_is_imm),
    .io_ctrl_sign_src1_is_pc(exu_step_io_ctrl_sign_src1_is_pc),
    .io_ctrl_sign_Writemem_en(exu_step_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(exu_step_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(exu_step_io_ctrl_sign_Wmask),
    .io_res2rd(exu_step_io_res2rd),
    .io_inst_valid(exu_step_io_inst_valid),
    .io_inst_store(exu_step_io_inst_store),
    .io_inst_load(exu_step_io_inst_load),
    .io_Mem_addr(exu_step_io_Mem_addr),
    .io_Mem_rdata(exu_step_io_Mem_rdata),
    .io_Mem_wdata(exu_step_io_Mem_wdata),
    .io_Mem_wstrb(exu_step_io_Mem_wstrb),
    .io_rdata_valid(exu_step_io_rdata_valid)
  );
  DPI dpi ( // @[top.scala 73:21]
    .flag(dpi_flag),
    .ecall_flag(dpi_ecall_flag)
  );
  assign io_inst = ifu_step_io_inst; // @[top.scala 25:13]
  assign io_pc = pc_now; // @[top.scala 16:11]
  assign io_pc_next = exu_step_io_pc_next; // @[top.scala 94:16]
  assign io_outval = exu_step_io_res2rd; // @[top.scala 69:15]
  assign io_step = diff_step; // @[top.scala 92:13]
  assign axi_clock = clock;
  assign axi_reset = reset;
  assign axi_io_axi_in_araddr = arbiter_io_axi_out_araddr; // @[top.scala 43:19]
  assign axi_io_axi_in_arvalid = arbiter_io_axi_out_arvalid; // @[top.scala 43:19]
  assign axi_io_axi_in_rready = arbiter_io_axi_out_rready; // @[top.scala 43:19]
  assign axi_io_axi_in_awaddr = arbiter_io_axi_out_awaddr; // @[top.scala 43:19]
  assign axi_io_axi_in_awvalid = arbiter_io_axi_out_awvalid; // @[top.scala 43:19]
  assign axi_io_axi_in_wdata = arbiter_io_axi_out_wdata; // @[top.scala 43:19]
  assign axi_io_axi_in_wstrb = arbiter_io_axi_out_wstrb; // @[top.scala 43:19]
  assign axi_io_axi_in_wvalid = arbiter_io_axi_out_wvalid; // @[top.scala 43:19]
  assign axi_io_axi_in_bready = arbiter_io_axi_out_bready; // @[top.scala 43:19]
  assign lsu_step_clock = clock;
  assign lsu_step_reset = reset;
  assign lsu_step_io_inst_store = exu_step_io_inst_store; // @[top.scala 61:28]
  assign lsu_step_io_inst_load = exu_step_io_inst_load; // @[top.scala 60:27]
  assign lsu_step_io_mem_addr = exu_step_io_Mem_addr; // @[top.scala 62:26]
  assign lsu_step_io_mem_wdata = exu_step_io_Mem_wdata; // @[top.scala 63:27]
  assign lsu_step_io_mem_wstrb = exu_step_io_Mem_wstrb; // @[top.scala 64:27]
  assign lsu_step_io_axi_in_arready = d_cache_io_to_lsu_arready; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_rdata = d_cache_io_to_lsu_rdata; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_rvalid = d_cache_io_to_lsu_rvalid; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_awready = d_cache_io_to_lsu_awready; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_wready = d_cache_io_to_lsu_wready; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_bvalid = d_cache_io_to_lsu_bvalid; // @[top.scala 36:24]
  assign arbiter_clock = clock;
  assign arbiter_reset = reset;
  assign arbiter_io_ifu_axi_in_araddr = i_cache_io_to_axi_araddr; // @[top.scala 26:27]
  assign arbiter_io_ifu_axi_in_arvalid = i_cache_io_to_axi_arvalid; // @[top.scala 26:27]
  assign arbiter_io_ifu_axi_in_rready = i_cache_io_to_axi_rready; // @[top.scala 26:27]
  assign arbiter_io_lsu_axi_in_araddr = d_cache_io_to_axi_araddr; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_arvalid = d_cache_io_to_axi_arvalid; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_rready = d_cache_io_to_axi_rready; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_awaddr = d_cache_io_to_axi_awaddr; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_awvalid = d_cache_io_to_axi_awvalid; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_wdata = d_cache_io_to_axi_wdata; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_wstrb = d_cache_io_to_axi_wstrb; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_wvalid = d_cache_io_to_axi_wvalid; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_bready = d_cache_io_to_axi_bready; // @[top.scala 34:27]
  assign arbiter_io_axi_in_arready = axi_io_axi_out_arready; // @[top.scala 42:23]
  assign arbiter_io_axi_in_rdata = axi_io_axi_out_rdata; // @[top.scala 42:23]
  assign arbiter_io_axi_in_rvalid = axi_io_axi_out_rvalid; // @[top.scala 42:23]
  assign arbiter_io_axi_in_awready = axi_io_axi_out_awready; // @[top.scala 42:23]
  assign arbiter_io_axi_in_wready = axi_io_axi_out_wready; // @[top.scala 42:23]
  assign arbiter_io_axi_in_bvalid = axi_io_axi_out_bvalid; // @[top.scala 42:23]
  assign ifu_step_clock = clock;
  assign ifu_step_reset = reset;
  assign ifu_step_io_pc = pc_now; // @[top.scala 24:20]
  assign ifu_step_io_pc_valid = pc_valid; // @[top.scala 89:26]
  assign ifu_step_io_axi_in_rdata = i_cache_io_to_ifu_rdata; // @[top.scala 28:24]
  assign ifu_step_io_axi_in_rvalid = i_cache_io_to_ifu_rvalid; // @[top.scala 28:24]
  assign i_cache_clock = clock;
  assign i_cache_reset = reset;
  assign i_cache_io_from_ifu_araddr = ifu_step_io_axi_out_araddr; // @[top.scala 29:25]
  assign i_cache_io_from_ifu_arvalid = ifu_step_io_axi_out_arvalid; // @[top.scala 29:25]
  assign i_cache_io_from_ifu_rready = ifu_step_io_axi_out_rready; // @[top.scala 29:25]
  assign i_cache_io_from_axi_rdata = arbiter_io_ifu_axi_out_rdata; // @[top.scala 27:25]
  assign i_cache_io_from_axi_rvalid = arbiter_io_ifu_axi_out_rvalid; // @[top.scala 27:25]
  assign d_cache_clock = clock;
  assign d_cache_reset = reset;
  assign d_cache_io_from_lsu_araddr = lsu_step_io_axi_out_araddr; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_arvalid = lsu_step_io_axi_out_arvalid; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_rready = lsu_step_io_axi_out_rready; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_awaddr = lsu_step_io_axi_out_awaddr; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_awvalid = lsu_step_io_axi_out_awvalid; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_wdata = lsu_step_io_axi_out_wdata; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_wstrb = lsu_step_io_axi_out_wstrb; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_wvalid = lsu_step_io_axi_out_wvalid; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_bready = lsu_step_io_axi_out_bready; // @[top.scala 37:25]
  assign d_cache_io_from_axi_arready = arbiter_io_lsu_axi_out_arready; // @[top.scala 35:25]
  assign d_cache_io_from_axi_rdata = arbiter_io_lsu_axi_out_rdata; // @[top.scala 35:25]
  assign d_cache_io_from_axi_rvalid = arbiter_io_lsu_axi_out_rvalid; // @[top.scala 35:25]
  assign d_cache_io_from_axi_awready = arbiter_io_lsu_axi_out_awready; // @[top.scala 35:25]
  assign d_cache_io_from_axi_wready = arbiter_io_lsu_axi_out_wready; // @[top.scala 35:25]
  assign d_cache_io_from_axi_bvalid = arbiter_io_lsu_axi_out_bvalid; // @[top.scala 35:25]
  assign idu_step_io_inst = ~ifu_step_io_inst_valid & ~pc_valid & ~execute_end ? ifu_step_io_inst_reg : ifu_step_io_inst
    ; // @[top.scala 96:28]
  assign exu_step_clock = clock;
  assign exu_step_reset = reset;
  assign exu_step_io_pc = pc_now; // @[top.scala 52:20]
  assign exu_step_io_inst_now = idu_step_io_inst_now; // @[top.scala 53:26]
  assign exu_step_io_rs1 = idu_step_io_rs1; // @[top.scala 55:21]
  assign exu_step_io_rs2 = idu_step_io_rs2; // @[top.scala 56:21]
  assign exu_step_io_rd = idu_step_io_rd; // @[top.scala 57:20]
  assign exu_step_io_imm = idu_step_io_imm; // @[top.scala 58:21]
  assign exu_step_io_ctrl_sign_reg_write = idu_step_io_ctrl_sign_reg_write; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_csr_write = idu_step_io_ctrl_sign_csr_write; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_src2_is_imm = idu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_src1_is_pc = idu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_Writemem_en = idu_step_io_ctrl_sign_Writemem_en; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_Readmem_en = idu_step_io_ctrl_sign_Readmem_en; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_Wmask = idu_step_io_ctrl_sign_Wmask; // @[top.scala 59:27]
  assign exu_step_io_inst_valid = ifu_step_io_inst_valid; // @[top.scala 68:28]
  assign exu_step_io_Mem_rdata = lsu_step_io_mem_rdata; // @[top.scala 65:27]
  assign exu_step_io_rdata_valid = lsu_step_io_axi_in_rvalid; // @[top.scala 66:29]
  assign dpi_flag = {{31'd0}, idu_step_io_inst_now == 32'h2}; // @[top.scala 74:17]
  assign dpi_ecall_flag = {{31'd0}, idu_step_io_inst_now == 32'h3d}; // @[top.scala 75:23]
  always @(posedge clock) begin
    if (reset) begin // @[top.scala 15:25]
      pc_now <= 64'h80000000; // @[top.scala 15:25]
    end else if (execute_end) begin // @[top.scala 93:18]
      pc_now <= exu_step_io_pc_next;
    end
    if (reset) begin // @[top.scala 17:30]
      execute_end <= 1'h0; // @[top.scala 17:30]
    end else if (exu_step_io_inst_store) begin // @[top.scala 85:23]
      execute_end <= lsu_step_io_axi_in_bvalid;
    end else if (exu_step_io_inst_load) begin // @[top.scala 85:76]
      execute_end <= lsu_step_io_axi_in_rvalid;
    end else begin
      execute_end <= ifu_step_io_inst_valid;
    end
    pc_valid <= reset | execute_end; // @[top.scala 87:{27,27} 88:14]
    if (reset) begin // @[top.scala 90:28]
      diff_step <= 1'h0; // @[top.scala 90:28]
    end else begin
      diff_step <= execute_end; // @[top.scala 91:15]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"pc : %x inst:%x execute_end : %d\n\n",pc_now,idu_step_io_inst,execute_end); // @[top.scala 86:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc_now = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  execute_end = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pc_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  diff_step = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
