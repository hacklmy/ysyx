module I_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_ifu_araddr,
  input         io_from_ifu_arvalid,
  input         io_from_ifu_rready,
  output [63:0] io_to_ifu_rdata,
  output        io_to_ifu_rlast,
  output        io_to_ifu_rvalid,
  output [31:0] io_to_axi_araddr,
  output [7:0]  io_to_axi_arlen,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rlast,
  input         io_from_axi_rvalid,
  output        io_cache_init,
  input         io_clear_cache
);
`ifdef RANDOMIZE_REG_INIT
  reg [511:0] _RAND_0;
  reg [511:0] _RAND_1;
  reg [511:0] _RAND_2;
  reg [511:0] _RAND_3;
  reg [511:0] _RAND_4;
  reg [511:0] _RAND_5;
  reg [511:0] _RAND_6;
  reg [511:0] _RAND_7;
  reg [511:0] _RAND_8;
  reg [511:0] _RAND_9;
  reg [511:0] _RAND_10;
  reg [511:0] _RAND_11;
  reg [511:0] _RAND_12;
  reg [511:0] _RAND_13;
  reg [511:0] _RAND_14;
  reg [511:0] _RAND_15;
  reg [511:0] _RAND_16;
  reg [511:0] _RAND_17;
  reg [511:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [511:0] _RAND_21;
  reg [511:0] _RAND_22;
  reg [511:0] _RAND_23;
  reg [511:0] _RAND_24;
  reg [511:0] _RAND_25;
  reg [511:0] _RAND_26;
  reg [511:0] _RAND_27;
  reg [511:0] _RAND_28;
  reg [511:0] _RAND_29;
  reg [511:0] _RAND_30;
  reg [511:0] _RAND_31;
  reg [511:0] _RAND_32;
  reg [511:0] _RAND_33;
  reg [511:0] _RAND_34;
  reg [511:0] _RAND_35;
  reg [511:0] _RAND_36;
  reg [511:0] _RAND_37;
  reg [511:0] _RAND_38;
  reg [511:0] _RAND_39;
  reg [511:0] _RAND_40;
  reg [511:0] _RAND_41;
  reg [511:0] _RAND_42;
  reg [511:0] _RAND_43;
  reg [511:0] _RAND_44;
  reg [511:0] _RAND_45;
  reg [511:0] _RAND_46;
  reg [511:0] _RAND_47;
  reg [511:0] _RAND_48;
  reg [511:0] _RAND_49;
  reg [511:0] _RAND_50;
  reg [511:0] _RAND_51;
  reg [511:0] _RAND_52;
  reg [511:0] _RAND_53;
  reg [511:0] _RAND_54;
  reg [511:0] _RAND_55;
  reg [511:0] _RAND_56;
  reg [511:0] _RAND_57;
  reg [511:0] _RAND_58;
  reg [511:0] _RAND_59;
  reg [511:0] _RAND_60;
  reg [511:0] _RAND_61;
  reg [511:0] _RAND_62;
  reg [511:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] ram_0_0; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_1; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_2; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_3; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_4; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_5; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_6; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_7; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_8; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_9; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_10; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_11; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_12; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_13; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_14; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_15; // @[i_cache.scala 19:24]
  reg [511:0] ram_1_0; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_1; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_2; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_3; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_4; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_5; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_6; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_7; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_8; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_9; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_10; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_11; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_12; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_13; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_14; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_15; // @[i_cache.scala 20:24]
  reg [511:0] ram_2_0; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_1; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_2; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_3; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_4; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_5; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_6; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_7; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_8; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_9; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_10; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_11; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_12; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_13; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_14; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_15; // @[i_cache.scala 21:24]
  reg [511:0] ram_3_0; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_1; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_2; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_3; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_4; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_5; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_6; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_7; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_8; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_9; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_10; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_11; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_12; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_13; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_14; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_15; // @[i_cache.scala 22:24]
  reg [31:0] tag_0_0; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_1; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_2; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_3; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_4; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_5; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_6; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_7; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_8; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_9; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_10; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_11; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_12; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_13; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_14; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_15; // @[i_cache.scala 23:24]
  reg [31:0] tag_1_0; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_1; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_2; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_3; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_4; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_5; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_6; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_7; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_8; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_9; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_10; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_11; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_12; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_13; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_14; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_15; // @[i_cache.scala 24:24]
  reg [31:0] tag_2_0; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_1; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_2; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_3; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_4; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_5; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_6; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_7; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_8; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_9; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_10; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_11; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_12; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_13; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_14; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_15; // @[i_cache.scala 25:24]
  reg [31:0] tag_3_0; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_1; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_2; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_3; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_4; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_5; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_6; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_7; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_8; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_9; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_10; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_11; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_12; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_13; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_14; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_15; // @[i_cache.scala 26:24]
  reg  valid_0_0; // @[i_cache.scala 27:26]
  reg  valid_0_1; // @[i_cache.scala 27:26]
  reg  valid_0_2; // @[i_cache.scala 27:26]
  reg  valid_0_3; // @[i_cache.scala 27:26]
  reg  valid_0_4; // @[i_cache.scala 27:26]
  reg  valid_0_5; // @[i_cache.scala 27:26]
  reg  valid_0_6; // @[i_cache.scala 27:26]
  reg  valid_0_7; // @[i_cache.scala 27:26]
  reg  valid_0_8; // @[i_cache.scala 27:26]
  reg  valid_0_9; // @[i_cache.scala 27:26]
  reg  valid_0_10; // @[i_cache.scala 27:26]
  reg  valid_0_11; // @[i_cache.scala 27:26]
  reg  valid_0_12; // @[i_cache.scala 27:26]
  reg  valid_0_13; // @[i_cache.scala 27:26]
  reg  valid_0_14; // @[i_cache.scala 27:26]
  reg  valid_0_15; // @[i_cache.scala 27:26]
  reg  valid_1_0; // @[i_cache.scala 28:26]
  reg  valid_1_1; // @[i_cache.scala 28:26]
  reg  valid_1_2; // @[i_cache.scala 28:26]
  reg  valid_1_3; // @[i_cache.scala 28:26]
  reg  valid_1_4; // @[i_cache.scala 28:26]
  reg  valid_1_5; // @[i_cache.scala 28:26]
  reg  valid_1_6; // @[i_cache.scala 28:26]
  reg  valid_1_7; // @[i_cache.scala 28:26]
  reg  valid_1_8; // @[i_cache.scala 28:26]
  reg  valid_1_9; // @[i_cache.scala 28:26]
  reg  valid_1_10; // @[i_cache.scala 28:26]
  reg  valid_1_11; // @[i_cache.scala 28:26]
  reg  valid_1_12; // @[i_cache.scala 28:26]
  reg  valid_1_13; // @[i_cache.scala 28:26]
  reg  valid_1_14; // @[i_cache.scala 28:26]
  reg  valid_1_15; // @[i_cache.scala 28:26]
  reg  valid_2_0; // @[i_cache.scala 29:26]
  reg  valid_2_1; // @[i_cache.scala 29:26]
  reg  valid_2_2; // @[i_cache.scala 29:26]
  reg  valid_2_3; // @[i_cache.scala 29:26]
  reg  valid_2_4; // @[i_cache.scala 29:26]
  reg  valid_2_5; // @[i_cache.scala 29:26]
  reg  valid_2_6; // @[i_cache.scala 29:26]
  reg  valid_2_7; // @[i_cache.scala 29:26]
  reg  valid_2_8; // @[i_cache.scala 29:26]
  reg  valid_2_9; // @[i_cache.scala 29:26]
  reg  valid_2_10; // @[i_cache.scala 29:26]
  reg  valid_2_11; // @[i_cache.scala 29:26]
  reg  valid_2_12; // @[i_cache.scala 29:26]
  reg  valid_2_13; // @[i_cache.scala 29:26]
  reg  valid_2_14; // @[i_cache.scala 29:26]
  reg  valid_2_15; // @[i_cache.scala 29:26]
  reg  valid_3_0; // @[i_cache.scala 30:26]
  reg  valid_3_1; // @[i_cache.scala 30:26]
  reg  valid_3_2; // @[i_cache.scala 30:26]
  reg  valid_3_3; // @[i_cache.scala 30:26]
  reg  valid_3_4; // @[i_cache.scala 30:26]
  reg  valid_3_5; // @[i_cache.scala 30:26]
  reg  valid_3_6; // @[i_cache.scala 30:26]
  reg  valid_3_7; // @[i_cache.scala 30:26]
  reg  valid_3_8; // @[i_cache.scala 30:26]
  reg  valid_3_9; // @[i_cache.scala 30:26]
  reg  valid_3_10; // @[i_cache.scala 30:26]
  reg  valid_3_11; // @[i_cache.scala 30:26]
  reg  valid_3_12; // @[i_cache.scala 30:26]
  reg  valid_3_13; // @[i_cache.scala 30:26]
  reg  valid_3_14; // @[i_cache.scala 30:26]
  reg  valid_3_15; // @[i_cache.scala 30:26]
  reg [63:0] receive_data_0; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_1; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_2; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_3; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_4; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_5; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_6; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_7; // @[i_cache.scala 38:31]
  reg [2:0] receive_num; // @[i_cache.scala 39:30]
  reg [7:0] quene_0; // @[i_cache.scala 40:24]
  reg [7:0] quene_1; // @[i_cache.scala 40:24]
  reg [7:0] quene_2; // @[i_cache.scala 40:24]
  reg [7:0] quene_3; // @[i_cache.scala 40:24]
  reg [7:0] quene_4; // @[i_cache.scala 40:24]
  reg [7:0] quene_5; // @[i_cache.scala 40:24]
  reg [7:0] quene_6; // @[i_cache.scala 40:24]
  reg [7:0] quene_7; // @[i_cache.scala 40:24]
  reg [7:0] quene_8; // @[i_cache.scala 40:24]
  reg [7:0] quene_9; // @[i_cache.scala 40:24]
  reg [7:0] quene_10; // @[i_cache.scala 40:24]
  reg [7:0] quene_11; // @[i_cache.scala 40:24]
  reg [7:0] quene_12; // @[i_cache.scala 40:24]
  reg [7:0] quene_13; // @[i_cache.scala 40:24]
  reg [7:0] quene_14; // @[i_cache.scala 40:24]
  reg [7:0] quene_15; // @[i_cache.scala 40:24]
  wire [5:0] offset = io_from_ifu_araddr[5:0]; // @[i_cache.scala 42:36]
  wire [3:0] index = io_from_ifu_araddr[9:6]; // @[i_cache.scala 43:35]
  wire [21:0] tag = io_from_ifu_araddr[31:10]; // @[i_cache.scala 44:33]
  wire [8:0] shift_bit = {offset, 3'h0}; // @[i_cache.scala 45:28]
  wire [31:0] _GEN_1 = 4'h1 == index ? tag_0_1 : tag_0_0; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_2 = 4'h2 == index ? tag_0_2 : _GEN_1; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_3 = 4'h3 == index ? tag_0_3 : _GEN_2; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_4 = 4'h4 == index ? tag_0_4 : _GEN_3; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_5 = 4'h5 == index ? tag_0_5 : _GEN_4; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_6 = 4'h6 == index ? tag_0_6 : _GEN_5; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_7 = 4'h7 == index ? tag_0_7 : _GEN_6; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_8 = 4'h8 == index ? tag_0_8 : _GEN_7; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_9 = 4'h9 == index ? tag_0_9 : _GEN_8; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_10 = 4'ha == index ? tag_0_10 : _GEN_9; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_11 = 4'hb == index ? tag_0_11 : _GEN_10; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_12 = 4'hc == index ? tag_0_12 : _GEN_11; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_13 = 4'hd == index ? tag_0_13 : _GEN_12; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_14 = 4'he == index ? tag_0_14 : _GEN_13; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_15 = 4'hf == index ? tag_0_15 : _GEN_14; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_2956 = {{10'd0}, tag}; // @[i_cache.scala 47:31]
  wire  _GEN_17 = 4'h1 == index ? valid_0_1 : valid_0_0; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_18 = 4'h2 == index ? valid_0_2 : _GEN_17; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_19 = 4'h3 == index ? valid_0_3 : _GEN_18; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_20 = 4'h4 == index ? valid_0_4 : _GEN_19; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_21 = 4'h5 == index ? valid_0_5 : _GEN_20; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_22 = 4'h6 == index ? valid_0_6 : _GEN_21; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_23 = 4'h7 == index ? valid_0_7 : _GEN_22; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_24 = 4'h8 == index ? valid_0_8 : _GEN_23; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_25 = 4'h9 == index ? valid_0_9 : _GEN_24; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_26 = 4'ha == index ? valid_0_10 : _GEN_25; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_27 = 4'hb == index ? valid_0_11 : _GEN_26; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_28 = 4'hc == index ? valid_0_12 : _GEN_27; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_29 = 4'hd == index ? valid_0_13 : _GEN_28; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_30 = 4'he == index ? valid_0_14 : _GEN_29; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_31 = 4'hf == index ? valid_0_15 : _GEN_30; // @[i_cache.scala 47:{57,57}]
  wire  way0_hit = _GEN_15 == _GEN_2956 & _GEN_31; // @[i_cache.scala 47:40]
  wire [31:0] _GEN_33 = 4'h1 == index ? tag_1_1 : tag_1_0; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_34 = 4'h2 == index ? tag_1_2 : _GEN_33; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_35 = 4'h3 == index ? tag_1_3 : _GEN_34; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_36 = 4'h4 == index ? tag_1_4 : _GEN_35; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_37 = 4'h5 == index ? tag_1_5 : _GEN_36; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_38 = 4'h6 == index ? tag_1_6 : _GEN_37; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_39 = 4'h7 == index ? tag_1_7 : _GEN_38; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_40 = 4'h8 == index ? tag_1_8 : _GEN_39; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_41 = 4'h9 == index ? tag_1_9 : _GEN_40; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_42 = 4'ha == index ? tag_1_10 : _GEN_41; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_43 = 4'hb == index ? tag_1_11 : _GEN_42; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_44 = 4'hc == index ? tag_1_12 : _GEN_43; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_45 = 4'hd == index ? tag_1_13 : _GEN_44; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_46 = 4'he == index ? tag_1_14 : _GEN_45; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_47 = 4'hf == index ? tag_1_15 : _GEN_46; // @[i_cache.scala 49:{31,31}]
  wire  _GEN_49 = 4'h1 == index ? valid_1_1 : valid_1_0; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_50 = 4'h2 == index ? valid_1_2 : _GEN_49; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_51 = 4'h3 == index ? valid_1_3 : _GEN_50; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_52 = 4'h4 == index ? valid_1_4 : _GEN_51; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_53 = 4'h5 == index ? valid_1_5 : _GEN_52; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_54 = 4'h6 == index ? valid_1_6 : _GEN_53; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_55 = 4'h7 == index ? valid_1_7 : _GEN_54; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_56 = 4'h8 == index ? valid_1_8 : _GEN_55; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_57 = 4'h9 == index ? valid_1_9 : _GEN_56; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_58 = 4'ha == index ? valid_1_10 : _GEN_57; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_59 = 4'hb == index ? valid_1_11 : _GEN_58; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_60 = 4'hc == index ? valid_1_12 : _GEN_59; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_61 = 4'hd == index ? valid_1_13 : _GEN_60; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_62 = 4'he == index ? valid_1_14 : _GEN_61; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_63 = 4'hf == index ? valid_1_15 : _GEN_62; // @[i_cache.scala 49:{57,57}]
  wire  way1_hit = _GEN_47 == _GEN_2956 & _GEN_63; // @[i_cache.scala 49:40]
  wire [31:0] _GEN_65 = 4'h1 == index ? tag_2_1 : tag_2_0; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_66 = 4'h2 == index ? tag_2_2 : _GEN_65; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_67 = 4'h3 == index ? tag_2_3 : _GEN_66; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_68 = 4'h4 == index ? tag_2_4 : _GEN_67; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_69 = 4'h5 == index ? tag_2_5 : _GEN_68; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_70 = 4'h6 == index ? tag_2_6 : _GEN_69; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_71 = 4'h7 == index ? tag_2_7 : _GEN_70; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_72 = 4'h8 == index ? tag_2_8 : _GEN_71; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_73 = 4'h9 == index ? tag_2_9 : _GEN_72; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_74 = 4'ha == index ? tag_2_10 : _GEN_73; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_75 = 4'hb == index ? tag_2_11 : _GEN_74; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_76 = 4'hc == index ? tag_2_12 : _GEN_75; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_77 = 4'hd == index ? tag_2_13 : _GEN_76; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_78 = 4'he == index ? tag_2_14 : _GEN_77; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_79 = 4'hf == index ? tag_2_15 : _GEN_78; // @[i_cache.scala 50:{31,31}]
  wire  _GEN_81 = 4'h1 == index ? valid_2_1 : valid_2_0; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_82 = 4'h2 == index ? valid_2_2 : _GEN_81; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_83 = 4'h3 == index ? valid_2_3 : _GEN_82; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_84 = 4'h4 == index ? valid_2_4 : _GEN_83; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_85 = 4'h5 == index ? valid_2_5 : _GEN_84; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_86 = 4'h6 == index ? valid_2_6 : _GEN_85; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_87 = 4'h7 == index ? valid_2_7 : _GEN_86; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_88 = 4'h8 == index ? valid_2_8 : _GEN_87; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_89 = 4'h9 == index ? valid_2_9 : _GEN_88; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_90 = 4'ha == index ? valid_2_10 : _GEN_89; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_91 = 4'hb == index ? valid_2_11 : _GEN_90; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_92 = 4'hc == index ? valid_2_12 : _GEN_91; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_93 = 4'hd == index ? valid_2_13 : _GEN_92; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_94 = 4'he == index ? valid_2_14 : _GEN_93; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_95 = 4'hf == index ? valid_2_15 : _GEN_94; // @[i_cache.scala 50:{57,57}]
  wire  way2_hit = _GEN_79 == _GEN_2956 & _GEN_95; // @[i_cache.scala 50:40]
  wire [31:0] _GEN_97 = 4'h1 == index ? tag_3_1 : tag_3_0; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_98 = 4'h2 == index ? tag_3_2 : _GEN_97; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_99 = 4'h3 == index ? tag_3_3 : _GEN_98; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_100 = 4'h4 == index ? tag_3_4 : _GEN_99; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_101 = 4'h5 == index ? tag_3_5 : _GEN_100; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_102 = 4'h6 == index ? tag_3_6 : _GEN_101; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_103 = 4'h7 == index ? tag_3_7 : _GEN_102; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_104 = 4'h8 == index ? tag_3_8 : _GEN_103; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_105 = 4'h9 == index ? tag_3_9 : _GEN_104; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_106 = 4'ha == index ? tag_3_10 : _GEN_105; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_107 = 4'hb == index ? tag_3_11 : _GEN_106; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_108 = 4'hc == index ? tag_3_12 : _GEN_107; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_109 = 4'hd == index ? tag_3_13 : _GEN_108; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_110 = 4'he == index ? tag_3_14 : _GEN_109; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_111 = 4'hf == index ? tag_3_15 : _GEN_110; // @[i_cache.scala 51:{31,31}]
  wire  _GEN_113 = 4'h1 == index ? valid_3_1 : valid_3_0; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_114 = 4'h2 == index ? valid_3_2 : _GEN_113; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_115 = 4'h3 == index ? valid_3_3 : _GEN_114; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_116 = 4'h4 == index ? valid_3_4 : _GEN_115; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_117 = 4'h5 == index ? valid_3_5 : _GEN_116; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_118 = 4'h6 == index ? valid_3_6 : _GEN_117; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_119 = 4'h7 == index ? valid_3_7 : _GEN_118; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_120 = 4'h8 == index ? valid_3_8 : _GEN_119; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_121 = 4'h9 == index ? valid_3_9 : _GEN_120; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_122 = 4'ha == index ? valid_3_10 : _GEN_121; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_123 = 4'hb == index ? valid_3_11 : _GEN_122; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_124 = 4'hc == index ? valid_3_12 : _GEN_123; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_125 = 4'hd == index ? valid_3_13 : _GEN_124; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_126 = 4'he == index ? valid_3_14 : _GEN_125; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_127 = 4'hf == index ? valid_3_15 : _GEN_126; // @[i_cache.scala 51:{57,57}]
  wire  way3_hit = _GEN_111 == _GEN_2956 & _GEN_127; // @[i_cache.scala 51:40]
  wire [2:0] _unuse_way_T_4 = ~_GEN_127 ? 3'h4 : 3'h0; // @[i_cache.scala 52:108]
  wire [2:0] _unuse_way_T_5 = ~_GEN_95 ? 3'h3 : _unuse_way_T_4; // @[i_cache.scala 52:79]
  wire [2:0] _unuse_way_T_6 = ~_GEN_63 ? 3'h2 : _unuse_way_T_5; // @[i_cache.scala 52:50]
  wire [2:0] unuse_way = ~_GEN_31 ? 3'h1 : _unuse_way_T_6; // @[i_cache.scala 52:21]
  reg [2:0] state; // @[i_cache.scala 54:24]
  wire  _T_4 = way0_hit | way1_hit | way2_hit | way3_hit; // @[i_cache.scala 65:46]
  wire [2:0] _GEN_130 = io_from_ifu_rready ? 3'h0 : state; // @[i_cache.scala 54:24 66:41 67:27]
  wire [63:0] _GEN_133 = 3'h0 == receive_num ? io_from_axi_rdata : receive_data_0; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_134 = 3'h1 == receive_num ? io_from_axi_rdata : receive_data_1; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_135 = 3'h2 == receive_num ? io_from_axi_rdata : receive_data_2; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_136 = 3'h3 == receive_num ? io_from_axi_rdata : receive_data_3; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_137 = 3'h4 == receive_num ? io_from_axi_rdata : receive_data_4; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_138 = 3'h5 == receive_num ? io_from_axi_rdata : receive_data_5; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_139 = 3'h6 == receive_num ? io_from_axi_rdata : receive_data_6; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_140 = 3'h7 == receive_num ? io_from_axi_rdata : receive_data_7; // @[i_cache.scala 38:31 76:{43,43}]
  wire [2:0] _receive_num_T_1 = receive_num + 3'h1; // @[i_cache.scala 77:44]
  wire [2:0] _GEN_141 = io_from_axi_rlast ? 3'h3 : state; // @[i_cache.scala 54:24 78:40 79:27]
  wire [63:0] _GEN_142 = io_from_axi_rvalid ? _GEN_133 : receive_data_0; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_143 = io_from_axi_rvalid ? _GEN_134 : receive_data_1; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_144 = io_from_axi_rvalid ? _GEN_135 : receive_data_2; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_145 = io_from_axi_rvalid ? _GEN_136 : receive_data_3; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_146 = io_from_axi_rvalid ? _GEN_137 : receive_data_4; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_147 = io_from_axi_rvalid ? _GEN_138 : receive_data_5; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_148 = io_from_axi_rvalid ? _GEN_139 : receive_data_6; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_149 = io_from_axi_rvalid ? _GEN_140 : receive_data_7; // @[i_cache.scala 38:31 75:37]
  wire [2:0] _GEN_150 = io_from_axi_rvalid ? _receive_num_T_1 : receive_num; // @[i_cache.scala 75:37 77:29 39:30]
  wire [2:0] _GEN_151 = io_from_axi_rvalid ? _GEN_141 : state; // @[i_cache.scala 54:24 75:37]
  wire [511:0] _ram_0_T = {receive_data_7,receive_data_6,receive_data_5,receive_data_4,receive_data_3,receive_data_2,
    receive_data_1,receive_data_0}; // @[Cat.scala 31:58]
  wire [511:0] _GEN_152 = 4'h0 == index ? _ram_0_T : ram_0_0; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_153 = 4'h1 == index ? _ram_0_T : ram_0_1; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_154 = 4'h2 == index ? _ram_0_T : ram_0_2; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_155 = 4'h3 == index ? _ram_0_T : ram_0_3; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_156 = 4'h4 == index ? _ram_0_T : ram_0_4; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_157 = 4'h5 == index ? _ram_0_T : ram_0_5; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_158 = 4'h6 == index ? _ram_0_T : ram_0_6; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_159 = 4'h7 == index ? _ram_0_T : ram_0_7; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_160 = 4'h8 == index ? _ram_0_T : ram_0_8; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_161 = 4'h9 == index ? _ram_0_T : ram_0_9; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_162 = 4'ha == index ? _ram_0_T : ram_0_10; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_163 = 4'hb == index ? _ram_0_T : ram_0_11; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_164 = 4'hc == index ? _ram_0_T : ram_0_12; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_165 = 4'hd == index ? _ram_0_T : ram_0_13; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_166 = 4'he == index ? _ram_0_T : ram_0_14; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_167 = 4'hf == index ? _ram_0_T : ram_0_15; // @[i_cache.scala 19:24 86:{30,30}]
  wire [31:0] _GEN_168 = 4'h0 == index ? _GEN_2956 : tag_0_0; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_169 = 4'h1 == index ? _GEN_2956 : tag_0_1; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_170 = 4'h2 == index ? _GEN_2956 : tag_0_2; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_171 = 4'h3 == index ? _GEN_2956 : tag_0_3; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_172 = 4'h4 == index ? _GEN_2956 : tag_0_4; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_173 = 4'h5 == index ? _GEN_2956 : tag_0_5; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_174 = 4'h6 == index ? _GEN_2956 : tag_0_6; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_175 = 4'h7 == index ? _GEN_2956 : tag_0_7; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_176 = 4'h8 == index ? _GEN_2956 : tag_0_8; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_177 = 4'h9 == index ? _GEN_2956 : tag_0_9; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_178 = 4'ha == index ? _GEN_2956 : tag_0_10; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_179 = 4'hb == index ? _GEN_2956 : tag_0_11; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_180 = 4'hc == index ? _GEN_2956 : tag_0_12; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_181 = 4'hd == index ? _GEN_2956 : tag_0_13; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_182 = 4'he == index ? _GEN_2956 : tag_0_14; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_183 = 4'hf == index ? _GEN_2956 : tag_0_15; // @[i_cache.scala 23:24 87:{30,30}]
  wire  _GEN_2969 = 4'h0 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_184 = 4'h0 == index | valid_0_0; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2970 = 4'h1 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_185 = 4'h1 == index | valid_0_1; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2971 = 4'h2 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_186 = 4'h2 == index | valid_0_2; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2972 = 4'h3 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_187 = 4'h3 == index | valid_0_3; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2973 = 4'h4 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_188 = 4'h4 == index | valid_0_4; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2974 = 4'h5 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_189 = 4'h5 == index | valid_0_5; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2975 = 4'h6 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_190 = 4'h6 == index | valid_0_6; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2976 = 4'h7 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_191 = 4'h7 == index | valid_0_7; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2977 = 4'h8 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_192 = 4'h8 == index | valid_0_8; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2978 = 4'h9 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_193 = 4'h9 == index | valid_0_9; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2979 = 4'ha == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_194 = 4'ha == index | valid_0_10; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2980 = 4'hb == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_195 = 4'hb == index | valid_0_11; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2981 = 4'hc == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_196 = 4'hc == index | valid_0_12; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2982 = 4'hd == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_197 = 4'hd == index | valid_0_13; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2983 = 4'he == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_198 = 4'he == index | valid_0_14; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2984 = 4'hf == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_199 = 4'hf == index | valid_0_15; // @[i_cache.scala 27:26 88:{32,32}]
  wire [7:0] _GEN_201 = 4'h1 == index ? quene_1 : quene_0; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_202 = 4'h2 == index ? quene_2 : _GEN_201; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_203 = 4'h3 == index ? quene_3 : _GEN_202; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_204 = 4'h4 == index ? quene_4 : _GEN_203; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_205 = 4'h5 == index ? quene_5 : _GEN_204; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_206 = 4'h6 == index ? quene_6 : _GEN_205; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_207 = 4'h7 == index ? quene_7 : _GEN_206; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_208 = 4'h8 == index ? quene_8 : _GEN_207; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_209 = 4'h9 == index ? quene_9 : _GEN_208; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_210 = 4'ha == index ? quene_10 : _GEN_209; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_211 = 4'hb == index ? quene_11 : _GEN_210; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_212 = 4'hc == index ? quene_12 : _GEN_211; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_213 = 4'hd == index ? quene_13 : _GEN_212; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_214 = 4'he == index ? quene_14 : _GEN_213; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_215 = 4'hf == index ? quene_15 : _GEN_214; // @[i_cache.scala 89:{46,46}]
  wire [9:0] _GEN_2985 = {_GEN_215, 2'h0}; // @[i_cache.scala 89:46]
  wire [10:0] _quene_T = {{1'd0}, _GEN_2985}; // @[i_cache.scala 89:46]
  wire [7:0] _GEN_216 = 4'h0 == index ? _quene_T[7:0] : quene_0; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_217 = 4'h1 == index ? _quene_T[7:0] : quene_1; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_218 = 4'h2 == index ? _quene_T[7:0] : quene_2; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_219 = 4'h3 == index ? _quene_T[7:0] : quene_3; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_220 = 4'h4 == index ? _quene_T[7:0] : quene_4; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_221 = 4'h5 == index ? _quene_T[7:0] : quene_5; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_222 = 4'h6 == index ? _quene_T[7:0] : quene_6; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_223 = 4'h7 == index ? _quene_T[7:0] : quene_7; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_224 = 4'h8 == index ? _quene_T[7:0] : quene_8; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_225 = 4'h9 == index ? _quene_T[7:0] : quene_9; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_226 = 4'ha == index ? _quene_T[7:0] : quene_10; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_227 = 4'hb == index ? _quene_T[7:0] : quene_11; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_228 = 4'hc == index ? _quene_T[7:0] : quene_12; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_229 = 4'hd == index ? _quene_T[7:0] : quene_13; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_230 = 4'he == index ? _quene_T[7:0] : quene_14; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_231 = 4'hf == index ? _quene_T[7:0] : quene_15; // @[i_cache.scala 40:24 89:{30,30}]
  wire [511:0] _GEN_232 = 4'h0 == index ? _ram_0_T : ram_1_0; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_233 = 4'h1 == index ? _ram_0_T : ram_1_1; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_234 = 4'h2 == index ? _ram_0_T : ram_1_2; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_235 = 4'h3 == index ? _ram_0_T : ram_1_3; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_236 = 4'h4 == index ? _ram_0_T : ram_1_4; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_237 = 4'h5 == index ? _ram_0_T : ram_1_5; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_238 = 4'h6 == index ? _ram_0_T : ram_1_6; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_239 = 4'h7 == index ? _ram_0_T : ram_1_7; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_240 = 4'h8 == index ? _ram_0_T : ram_1_8; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_241 = 4'h9 == index ? _ram_0_T : ram_1_9; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_242 = 4'ha == index ? _ram_0_T : ram_1_10; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_243 = 4'hb == index ? _ram_0_T : ram_1_11; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_244 = 4'hc == index ? _ram_0_T : ram_1_12; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_245 = 4'hd == index ? _ram_0_T : ram_1_13; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_246 = 4'he == index ? _ram_0_T : ram_1_14; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_247 = 4'hf == index ? _ram_0_T : ram_1_15; // @[i_cache.scala 20:24 91:{30,30}]
  wire [31:0] _GEN_248 = 4'h0 == index ? _GEN_2956 : tag_1_0; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_249 = 4'h1 == index ? _GEN_2956 : tag_1_1; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_250 = 4'h2 == index ? _GEN_2956 : tag_1_2; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_251 = 4'h3 == index ? _GEN_2956 : tag_1_3; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_252 = 4'h4 == index ? _GEN_2956 : tag_1_4; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_253 = 4'h5 == index ? _GEN_2956 : tag_1_5; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_254 = 4'h6 == index ? _GEN_2956 : tag_1_6; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_255 = 4'h7 == index ? _GEN_2956 : tag_1_7; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_256 = 4'h8 == index ? _GEN_2956 : tag_1_8; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_257 = 4'h9 == index ? _GEN_2956 : tag_1_9; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_258 = 4'ha == index ? _GEN_2956 : tag_1_10; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_259 = 4'hb == index ? _GEN_2956 : tag_1_11; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_260 = 4'hc == index ? _GEN_2956 : tag_1_12; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_261 = 4'hd == index ? _GEN_2956 : tag_1_13; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_262 = 4'he == index ? _GEN_2956 : tag_1_14; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_263 = 4'hf == index ? _GEN_2956 : tag_1_15; // @[i_cache.scala 24:24 92:{30,30}]
  wire  _GEN_264 = _GEN_2969 | valid_1_0; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_265 = _GEN_2970 | valid_1_1; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_266 = _GEN_2971 | valid_1_2; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_267 = _GEN_2972 | valid_1_3; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_268 = _GEN_2973 | valid_1_4; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_269 = _GEN_2974 | valid_1_5; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_270 = _GEN_2975 | valid_1_6; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_271 = _GEN_2976 | valid_1_7; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_272 = _GEN_2977 | valid_1_8; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_273 = _GEN_2978 | valid_1_9; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_274 = _GEN_2979 | valid_1_10; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_275 = _GEN_2980 | valid_1_11; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_276 = _GEN_2981 | valid_1_12; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_277 = _GEN_2982 | valid_1_13; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_278 = _GEN_2983 | valid_1_14; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_279 = _GEN_2984 | valid_1_15; // @[i_cache.scala 28:26 93:{32,32}]
  wire [10:0] _quene_T_2 = _quene_T | 11'h1; // @[i_cache.scala 94:55]
  wire [7:0] _GEN_280 = 4'h0 == index ? _quene_T_2[7:0] : quene_0; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_281 = 4'h1 == index ? _quene_T_2[7:0] : quene_1; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_282 = 4'h2 == index ? _quene_T_2[7:0] : quene_2; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_283 = 4'h3 == index ? _quene_T_2[7:0] : quene_3; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_284 = 4'h4 == index ? _quene_T_2[7:0] : quene_4; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_285 = 4'h5 == index ? _quene_T_2[7:0] : quene_5; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_286 = 4'h6 == index ? _quene_T_2[7:0] : quene_6; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_287 = 4'h7 == index ? _quene_T_2[7:0] : quene_7; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_288 = 4'h8 == index ? _quene_T_2[7:0] : quene_8; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_289 = 4'h9 == index ? _quene_T_2[7:0] : quene_9; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_290 = 4'ha == index ? _quene_T_2[7:0] : quene_10; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_291 = 4'hb == index ? _quene_T_2[7:0] : quene_11; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_292 = 4'hc == index ? _quene_T_2[7:0] : quene_12; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_293 = 4'hd == index ? _quene_T_2[7:0] : quene_13; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_294 = 4'he == index ? _quene_T_2[7:0] : quene_14; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_295 = 4'hf == index ? _quene_T_2[7:0] : quene_15; // @[i_cache.scala 40:24 94:{30,30}]
  wire [511:0] _GEN_296 = 4'h0 == index ? _ram_0_T : ram_2_0; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_297 = 4'h1 == index ? _ram_0_T : ram_2_1; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_298 = 4'h2 == index ? _ram_0_T : ram_2_2; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_299 = 4'h3 == index ? _ram_0_T : ram_2_3; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_300 = 4'h4 == index ? _ram_0_T : ram_2_4; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_301 = 4'h5 == index ? _ram_0_T : ram_2_5; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_302 = 4'h6 == index ? _ram_0_T : ram_2_6; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_303 = 4'h7 == index ? _ram_0_T : ram_2_7; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_304 = 4'h8 == index ? _ram_0_T : ram_2_8; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_305 = 4'h9 == index ? _ram_0_T : ram_2_9; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_306 = 4'ha == index ? _ram_0_T : ram_2_10; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_307 = 4'hb == index ? _ram_0_T : ram_2_11; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_308 = 4'hc == index ? _ram_0_T : ram_2_12; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_309 = 4'hd == index ? _ram_0_T : ram_2_13; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_310 = 4'he == index ? _ram_0_T : ram_2_14; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_311 = 4'hf == index ? _ram_0_T : ram_2_15; // @[i_cache.scala 21:24 96:{30,30}]
  wire [31:0] _GEN_312 = 4'h0 == index ? _GEN_2956 : tag_2_0; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_313 = 4'h1 == index ? _GEN_2956 : tag_2_1; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_314 = 4'h2 == index ? _GEN_2956 : tag_2_2; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_315 = 4'h3 == index ? _GEN_2956 : tag_2_3; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_316 = 4'h4 == index ? _GEN_2956 : tag_2_4; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_317 = 4'h5 == index ? _GEN_2956 : tag_2_5; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_318 = 4'h6 == index ? _GEN_2956 : tag_2_6; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_319 = 4'h7 == index ? _GEN_2956 : tag_2_7; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_320 = 4'h8 == index ? _GEN_2956 : tag_2_8; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_321 = 4'h9 == index ? _GEN_2956 : tag_2_9; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_322 = 4'ha == index ? _GEN_2956 : tag_2_10; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_323 = 4'hb == index ? _GEN_2956 : tag_2_11; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_324 = 4'hc == index ? _GEN_2956 : tag_2_12; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_325 = 4'hd == index ? _GEN_2956 : tag_2_13; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_326 = 4'he == index ? _GEN_2956 : tag_2_14; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_327 = 4'hf == index ? _GEN_2956 : tag_2_15; // @[i_cache.scala 25:24 97:{30,30}]
  wire  _GEN_328 = _GEN_2969 | valid_2_0; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_329 = _GEN_2970 | valid_2_1; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_330 = _GEN_2971 | valid_2_2; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_331 = _GEN_2972 | valid_2_3; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_332 = _GEN_2973 | valid_2_4; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_333 = _GEN_2974 | valid_2_5; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_334 = _GEN_2975 | valid_2_6; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_335 = _GEN_2976 | valid_2_7; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_336 = _GEN_2977 | valid_2_8; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_337 = _GEN_2978 | valid_2_9; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_338 = _GEN_2979 | valid_2_10; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_339 = _GEN_2980 | valid_2_11; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_340 = _GEN_2981 | valid_2_12; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_341 = _GEN_2982 | valid_2_13; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_342 = _GEN_2983 | valid_2_14; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_343 = _GEN_2984 | valid_2_15; // @[i_cache.scala 29:26 98:{32,32}]
  wire [10:0] _quene_T_4 = _quene_T | 11'h2; // @[i_cache.scala 99:55]
  wire [7:0] _GEN_344 = 4'h0 == index ? _quene_T_4[7:0] : quene_0; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_345 = 4'h1 == index ? _quene_T_4[7:0] : quene_1; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_346 = 4'h2 == index ? _quene_T_4[7:0] : quene_2; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_347 = 4'h3 == index ? _quene_T_4[7:0] : quene_3; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_348 = 4'h4 == index ? _quene_T_4[7:0] : quene_4; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_349 = 4'h5 == index ? _quene_T_4[7:0] : quene_5; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_350 = 4'h6 == index ? _quene_T_4[7:0] : quene_6; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_351 = 4'h7 == index ? _quene_T_4[7:0] : quene_7; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_352 = 4'h8 == index ? _quene_T_4[7:0] : quene_8; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_353 = 4'h9 == index ? _quene_T_4[7:0] : quene_9; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_354 = 4'ha == index ? _quene_T_4[7:0] : quene_10; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_355 = 4'hb == index ? _quene_T_4[7:0] : quene_11; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_356 = 4'hc == index ? _quene_T_4[7:0] : quene_12; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_357 = 4'hd == index ? _quene_T_4[7:0] : quene_13; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_358 = 4'he == index ? _quene_T_4[7:0] : quene_14; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_359 = 4'hf == index ? _quene_T_4[7:0] : quene_15; // @[i_cache.scala 40:24 99:{30,30}]
  wire [511:0] _GEN_360 = 4'h0 == index ? _ram_0_T : ram_3_0; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_361 = 4'h1 == index ? _ram_0_T : ram_3_1; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_362 = 4'h2 == index ? _ram_0_T : ram_3_2; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_363 = 4'h3 == index ? _ram_0_T : ram_3_3; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_364 = 4'h4 == index ? _ram_0_T : ram_3_4; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_365 = 4'h5 == index ? _ram_0_T : ram_3_5; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_366 = 4'h6 == index ? _ram_0_T : ram_3_6; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_367 = 4'h7 == index ? _ram_0_T : ram_3_7; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_368 = 4'h8 == index ? _ram_0_T : ram_3_8; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_369 = 4'h9 == index ? _ram_0_T : ram_3_9; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_370 = 4'ha == index ? _ram_0_T : ram_3_10; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_371 = 4'hb == index ? _ram_0_T : ram_3_11; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_372 = 4'hc == index ? _ram_0_T : ram_3_12; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_373 = 4'hd == index ? _ram_0_T : ram_3_13; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_374 = 4'he == index ? _ram_0_T : ram_3_14; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_375 = 4'hf == index ? _ram_0_T : ram_3_15; // @[i_cache.scala 101:{30,30} 22:24]
  wire [31:0] _GEN_376 = 4'h0 == index ? _GEN_2956 : tag_3_0; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_377 = 4'h1 == index ? _GEN_2956 : tag_3_1; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_378 = 4'h2 == index ? _GEN_2956 : tag_3_2; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_379 = 4'h3 == index ? _GEN_2956 : tag_3_3; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_380 = 4'h4 == index ? _GEN_2956 : tag_3_4; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_381 = 4'h5 == index ? _GEN_2956 : tag_3_5; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_382 = 4'h6 == index ? _GEN_2956 : tag_3_6; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_383 = 4'h7 == index ? _GEN_2956 : tag_3_7; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_384 = 4'h8 == index ? _GEN_2956 : tag_3_8; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_385 = 4'h9 == index ? _GEN_2956 : tag_3_9; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_386 = 4'ha == index ? _GEN_2956 : tag_3_10; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_387 = 4'hb == index ? _GEN_2956 : tag_3_11; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_388 = 4'hc == index ? _GEN_2956 : tag_3_12; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_389 = 4'hd == index ? _GEN_2956 : tag_3_13; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_390 = 4'he == index ? _GEN_2956 : tag_3_14; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_391 = 4'hf == index ? _GEN_2956 : tag_3_15; // @[i_cache.scala 102:{30,30} 26:24]
  wire  _GEN_392 = _GEN_2969 | valid_3_0; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_393 = _GEN_2970 | valid_3_1; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_394 = _GEN_2971 | valid_3_2; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_395 = _GEN_2972 | valid_3_3; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_396 = _GEN_2973 | valid_3_4; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_397 = _GEN_2974 | valid_3_5; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_398 = _GEN_2975 | valid_3_6; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_399 = _GEN_2976 | valid_3_7; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_400 = _GEN_2977 | valid_3_8; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_401 = _GEN_2978 | valid_3_9; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_402 = _GEN_2979 | valid_3_10; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_403 = _GEN_2980 | valid_3_11; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_404 = _GEN_2981 | valid_3_12; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_405 = _GEN_2982 | valid_3_13; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_406 = _GEN_2983 | valid_3_14; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_407 = _GEN_2984 | valid_3_15; // @[i_cache.scala 103:{32,32} 30:26]
  wire [10:0] _quene_T_6 = _quene_T | 11'h3; // @[i_cache.scala 104:55]
  wire [7:0] _GEN_408 = 4'h0 == index ? _quene_T_6[7:0] : quene_0; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_409 = 4'h1 == index ? _quene_T_6[7:0] : quene_1; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_410 = 4'h2 == index ? _quene_T_6[7:0] : quene_2; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_411 = 4'h3 == index ? _quene_T_6[7:0] : quene_3; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_412 = 4'h4 == index ? _quene_T_6[7:0] : quene_4; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_413 = 4'h5 == index ? _quene_T_6[7:0] : quene_5; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_414 = 4'h6 == index ? _quene_T_6[7:0] : quene_6; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_415 = 4'h7 == index ? _quene_T_6[7:0] : quene_7; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_416 = 4'h8 == index ? _quene_T_6[7:0] : quene_8; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_417 = 4'h9 == index ? _quene_T_6[7:0] : quene_9; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_418 = 4'ha == index ? _quene_T_6[7:0] : quene_10; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_419 = 4'hb == index ? _quene_T_6[7:0] : quene_11; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_420 = 4'hc == index ? _quene_T_6[7:0] : quene_12; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_421 = 4'hd == index ? _quene_T_6[7:0] : quene_13; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_422 = 4'he == index ? _quene_T_6[7:0] : quene_14; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_423 = 4'hf == index ? _quene_T_6[7:0] : quene_15; // @[i_cache.scala 104:{30,30} 40:24]
  wire [511:0] _GEN_680 = _GEN_215[7:6] == 2'h2 ? _GEN_296 : ram_2_0; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_681 = _GEN_215[7:6] == 2'h2 ? _GEN_297 : ram_2_1; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_682 = _GEN_215[7:6] == 2'h2 ? _GEN_298 : ram_2_2; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_683 = _GEN_215[7:6] == 2'h2 ? _GEN_299 : ram_2_3; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_684 = _GEN_215[7:6] == 2'h2 ? _GEN_300 : ram_2_4; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_685 = _GEN_215[7:6] == 2'h2 ? _GEN_301 : ram_2_5; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_686 = _GEN_215[7:6] == 2'h2 ? _GEN_302 : ram_2_6; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_687 = _GEN_215[7:6] == 2'h2 ? _GEN_303 : ram_2_7; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_688 = _GEN_215[7:6] == 2'h2 ? _GEN_304 : ram_2_8; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_689 = _GEN_215[7:6] == 2'h2 ? _GEN_305 : ram_2_9; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_690 = _GEN_215[7:6] == 2'h2 ? _GEN_306 : ram_2_10; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_691 = _GEN_215[7:6] == 2'h2 ? _GEN_307 : ram_2_11; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_692 = _GEN_215[7:6] == 2'h2 ? _GEN_308 : ram_2_12; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_693 = _GEN_215[7:6] == 2'h2 ? _GEN_309 : ram_2_13; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_694 = _GEN_215[7:6] == 2'h2 ? _GEN_310 : ram_2_14; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_695 = _GEN_215[7:6] == 2'h2 ? _GEN_311 : ram_2_15; // @[i_cache.scala 116:52 21:24]
  wire [31:0] _GEN_696 = _GEN_215[7:6] == 2'h2 ? _GEN_312 : tag_2_0; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_697 = _GEN_215[7:6] == 2'h2 ? _GEN_313 : tag_2_1; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_698 = _GEN_215[7:6] == 2'h2 ? _GEN_314 : tag_2_2; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_699 = _GEN_215[7:6] == 2'h2 ? _GEN_315 : tag_2_3; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_700 = _GEN_215[7:6] == 2'h2 ? _GEN_316 : tag_2_4; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_701 = _GEN_215[7:6] == 2'h2 ? _GEN_317 : tag_2_5; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_702 = _GEN_215[7:6] == 2'h2 ? _GEN_318 : tag_2_6; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_703 = _GEN_215[7:6] == 2'h2 ? _GEN_319 : tag_2_7; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_704 = _GEN_215[7:6] == 2'h2 ? _GEN_320 : tag_2_8; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_705 = _GEN_215[7:6] == 2'h2 ? _GEN_321 : tag_2_9; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_706 = _GEN_215[7:6] == 2'h2 ? _GEN_322 : tag_2_10; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_707 = _GEN_215[7:6] == 2'h2 ? _GEN_323 : tag_2_11; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_708 = _GEN_215[7:6] == 2'h2 ? _GEN_324 : tag_2_12; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_709 = _GEN_215[7:6] == 2'h2 ? _GEN_325 : tag_2_13; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_710 = _GEN_215[7:6] == 2'h2 ? _GEN_326 : tag_2_14; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_711 = _GEN_215[7:6] == 2'h2 ? _GEN_327 : tag_2_15; // @[i_cache.scala 116:52 25:24]
  wire  _GEN_712 = _GEN_215[7:6] == 2'h2 ? _GEN_328 : valid_2_0; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_713 = _GEN_215[7:6] == 2'h2 ? _GEN_329 : valid_2_1; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_714 = _GEN_215[7:6] == 2'h2 ? _GEN_330 : valid_2_2; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_715 = _GEN_215[7:6] == 2'h2 ? _GEN_331 : valid_2_3; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_716 = _GEN_215[7:6] == 2'h2 ? _GEN_332 : valid_2_4; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_717 = _GEN_215[7:6] == 2'h2 ? _GEN_333 : valid_2_5; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_718 = _GEN_215[7:6] == 2'h2 ? _GEN_334 : valid_2_6; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_719 = _GEN_215[7:6] == 2'h2 ? _GEN_335 : valid_2_7; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_720 = _GEN_215[7:6] == 2'h2 ? _GEN_336 : valid_2_8; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_721 = _GEN_215[7:6] == 2'h2 ? _GEN_337 : valid_2_9; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_722 = _GEN_215[7:6] == 2'h2 ? _GEN_338 : valid_2_10; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_723 = _GEN_215[7:6] == 2'h2 ? _GEN_339 : valid_2_11; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_724 = _GEN_215[7:6] == 2'h2 ? _GEN_340 : valid_2_12; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_725 = _GEN_215[7:6] == 2'h2 ? _GEN_341 : valid_2_13; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_726 = _GEN_215[7:6] == 2'h2 ? _GEN_342 : valid_2_14; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_727 = _GEN_215[7:6] == 2'h2 ? _GEN_343 : valid_2_15; // @[i_cache.scala 116:52 29:26]
  wire [7:0] _GEN_728 = _GEN_215[7:6] == 2'h2 ? _GEN_344 : _GEN_408; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_729 = _GEN_215[7:6] == 2'h2 ? _GEN_345 : _GEN_409; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_730 = _GEN_215[7:6] == 2'h2 ? _GEN_346 : _GEN_410; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_731 = _GEN_215[7:6] == 2'h2 ? _GEN_347 : _GEN_411; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_732 = _GEN_215[7:6] == 2'h2 ? _GEN_348 : _GEN_412; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_733 = _GEN_215[7:6] == 2'h2 ? _GEN_349 : _GEN_413; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_734 = _GEN_215[7:6] == 2'h2 ? _GEN_350 : _GEN_414; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_735 = _GEN_215[7:6] == 2'h2 ? _GEN_351 : _GEN_415; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_736 = _GEN_215[7:6] == 2'h2 ? _GEN_352 : _GEN_416; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_737 = _GEN_215[7:6] == 2'h2 ? _GEN_353 : _GEN_417; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_738 = _GEN_215[7:6] == 2'h2 ? _GEN_354 : _GEN_418; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_739 = _GEN_215[7:6] == 2'h2 ? _GEN_355 : _GEN_419; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_740 = _GEN_215[7:6] == 2'h2 ? _GEN_356 : _GEN_420; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_741 = _GEN_215[7:6] == 2'h2 ? _GEN_357 : _GEN_421; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_742 = _GEN_215[7:6] == 2'h2 ? _GEN_358 : _GEN_422; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_743 = _GEN_215[7:6] == 2'h2 ? _GEN_359 : _GEN_423; // @[i_cache.scala 116:52]
  wire [511:0] _GEN_744 = _GEN_215[7:6] == 2'h2 ? ram_3_0 : _GEN_360; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_745 = _GEN_215[7:6] == 2'h2 ? ram_3_1 : _GEN_361; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_746 = _GEN_215[7:6] == 2'h2 ? ram_3_2 : _GEN_362; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_747 = _GEN_215[7:6] == 2'h2 ? ram_3_3 : _GEN_363; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_748 = _GEN_215[7:6] == 2'h2 ? ram_3_4 : _GEN_364; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_749 = _GEN_215[7:6] == 2'h2 ? ram_3_5 : _GEN_365; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_750 = _GEN_215[7:6] == 2'h2 ? ram_3_6 : _GEN_366; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_751 = _GEN_215[7:6] == 2'h2 ? ram_3_7 : _GEN_367; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_752 = _GEN_215[7:6] == 2'h2 ? ram_3_8 : _GEN_368; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_753 = _GEN_215[7:6] == 2'h2 ? ram_3_9 : _GEN_369; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_754 = _GEN_215[7:6] == 2'h2 ? ram_3_10 : _GEN_370; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_755 = _GEN_215[7:6] == 2'h2 ? ram_3_11 : _GEN_371; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_756 = _GEN_215[7:6] == 2'h2 ? ram_3_12 : _GEN_372; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_757 = _GEN_215[7:6] == 2'h2 ? ram_3_13 : _GEN_373; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_758 = _GEN_215[7:6] == 2'h2 ? ram_3_14 : _GEN_374; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_759 = _GEN_215[7:6] == 2'h2 ? ram_3_15 : _GEN_375; // @[i_cache.scala 116:52 22:24]
  wire [31:0] _GEN_760 = _GEN_215[7:6] == 2'h2 ? tag_3_0 : _GEN_376; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_761 = _GEN_215[7:6] == 2'h2 ? tag_3_1 : _GEN_377; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_762 = _GEN_215[7:6] == 2'h2 ? tag_3_2 : _GEN_378; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_763 = _GEN_215[7:6] == 2'h2 ? tag_3_3 : _GEN_379; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_764 = _GEN_215[7:6] == 2'h2 ? tag_3_4 : _GEN_380; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_765 = _GEN_215[7:6] == 2'h2 ? tag_3_5 : _GEN_381; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_766 = _GEN_215[7:6] == 2'h2 ? tag_3_6 : _GEN_382; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_767 = _GEN_215[7:6] == 2'h2 ? tag_3_7 : _GEN_383; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_768 = _GEN_215[7:6] == 2'h2 ? tag_3_8 : _GEN_384; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_769 = _GEN_215[7:6] == 2'h2 ? tag_3_9 : _GEN_385; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_770 = _GEN_215[7:6] == 2'h2 ? tag_3_10 : _GEN_386; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_771 = _GEN_215[7:6] == 2'h2 ? tag_3_11 : _GEN_387; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_772 = _GEN_215[7:6] == 2'h2 ? tag_3_12 : _GEN_388; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_773 = _GEN_215[7:6] == 2'h2 ? tag_3_13 : _GEN_389; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_774 = _GEN_215[7:6] == 2'h2 ? tag_3_14 : _GEN_390; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_775 = _GEN_215[7:6] == 2'h2 ? tag_3_15 : _GEN_391; // @[i_cache.scala 116:52 26:24]
  wire  _GEN_776 = _GEN_215[7:6] == 2'h2 ? valid_3_0 : _GEN_392; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_777 = _GEN_215[7:6] == 2'h2 ? valid_3_1 : _GEN_393; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_778 = _GEN_215[7:6] == 2'h2 ? valid_3_2 : _GEN_394; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_779 = _GEN_215[7:6] == 2'h2 ? valid_3_3 : _GEN_395; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_780 = _GEN_215[7:6] == 2'h2 ? valid_3_4 : _GEN_396; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_781 = _GEN_215[7:6] == 2'h2 ? valid_3_5 : _GEN_397; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_782 = _GEN_215[7:6] == 2'h2 ? valid_3_6 : _GEN_398; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_783 = _GEN_215[7:6] == 2'h2 ? valid_3_7 : _GEN_399; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_784 = _GEN_215[7:6] == 2'h2 ? valid_3_8 : _GEN_400; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_785 = _GEN_215[7:6] == 2'h2 ? valid_3_9 : _GEN_401; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_786 = _GEN_215[7:6] == 2'h2 ? valid_3_10 : _GEN_402; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_787 = _GEN_215[7:6] == 2'h2 ? valid_3_11 : _GEN_403; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_788 = _GEN_215[7:6] == 2'h2 ? valid_3_12 : _GEN_404; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_789 = _GEN_215[7:6] == 2'h2 ? valid_3_13 : _GEN_405; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_790 = _GEN_215[7:6] == 2'h2 ? valid_3_14 : _GEN_406; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_791 = _GEN_215[7:6] == 2'h2 ? valid_3_15 : _GEN_407; // @[i_cache.scala 116:52 30:26]
  wire [511:0] _GEN_792 = _GEN_215[7:6] == 2'h1 ? _GEN_232 : ram_1_0; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_793 = _GEN_215[7:6] == 2'h1 ? _GEN_233 : ram_1_1; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_794 = _GEN_215[7:6] == 2'h1 ? _GEN_234 : ram_1_2; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_795 = _GEN_215[7:6] == 2'h1 ? _GEN_235 : ram_1_3; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_796 = _GEN_215[7:6] == 2'h1 ? _GEN_236 : ram_1_4; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_797 = _GEN_215[7:6] == 2'h1 ? _GEN_237 : ram_1_5; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_798 = _GEN_215[7:6] == 2'h1 ? _GEN_238 : ram_1_6; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_799 = _GEN_215[7:6] == 2'h1 ? _GEN_239 : ram_1_7; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_800 = _GEN_215[7:6] == 2'h1 ? _GEN_240 : ram_1_8; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_801 = _GEN_215[7:6] == 2'h1 ? _GEN_241 : ram_1_9; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_802 = _GEN_215[7:6] == 2'h1 ? _GEN_242 : ram_1_10; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_803 = _GEN_215[7:6] == 2'h1 ? _GEN_243 : ram_1_11; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_804 = _GEN_215[7:6] == 2'h1 ? _GEN_244 : ram_1_12; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_805 = _GEN_215[7:6] == 2'h1 ? _GEN_245 : ram_1_13; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_806 = _GEN_215[7:6] == 2'h1 ? _GEN_246 : ram_1_14; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_807 = _GEN_215[7:6] == 2'h1 ? _GEN_247 : ram_1_15; // @[i_cache.scala 111:52 20:24]
  wire [31:0] _GEN_808 = _GEN_215[7:6] == 2'h1 ? _GEN_248 : tag_1_0; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_809 = _GEN_215[7:6] == 2'h1 ? _GEN_249 : tag_1_1; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_810 = _GEN_215[7:6] == 2'h1 ? _GEN_250 : tag_1_2; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_811 = _GEN_215[7:6] == 2'h1 ? _GEN_251 : tag_1_3; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_812 = _GEN_215[7:6] == 2'h1 ? _GEN_252 : tag_1_4; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_813 = _GEN_215[7:6] == 2'h1 ? _GEN_253 : tag_1_5; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_814 = _GEN_215[7:6] == 2'h1 ? _GEN_254 : tag_1_6; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_815 = _GEN_215[7:6] == 2'h1 ? _GEN_255 : tag_1_7; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_816 = _GEN_215[7:6] == 2'h1 ? _GEN_256 : tag_1_8; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_817 = _GEN_215[7:6] == 2'h1 ? _GEN_257 : tag_1_9; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_818 = _GEN_215[7:6] == 2'h1 ? _GEN_258 : tag_1_10; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_819 = _GEN_215[7:6] == 2'h1 ? _GEN_259 : tag_1_11; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_820 = _GEN_215[7:6] == 2'h1 ? _GEN_260 : tag_1_12; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_821 = _GEN_215[7:6] == 2'h1 ? _GEN_261 : tag_1_13; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_822 = _GEN_215[7:6] == 2'h1 ? _GEN_262 : tag_1_14; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_823 = _GEN_215[7:6] == 2'h1 ? _GEN_263 : tag_1_15; // @[i_cache.scala 111:52 24:24]
  wire  _GEN_824 = _GEN_215[7:6] == 2'h1 ? _GEN_264 : valid_1_0; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_825 = _GEN_215[7:6] == 2'h1 ? _GEN_265 : valid_1_1; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_826 = _GEN_215[7:6] == 2'h1 ? _GEN_266 : valid_1_2; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_827 = _GEN_215[7:6] == 2'h1 ? _GEN_267 : valid_1_3; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_828 = _GEN_215[7:6] == 2'h1 ? _GEN_268 : valid_1_4; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_829 = _GEN_215[7:6] == 2'h1 ? _GEN_269 : valid_1_5; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_830 = _GEN_215[7:6] == 2'h1 ? _GEN_270 : valid_1_6; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_831 = _GEN_215[7:6] == 2'h1 ? _GEN_271 : valid_1_7; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_832 = _GEN_215[7:6] == 2'h1 ? _GEN_272 : valid_1_8; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_833 = _GEN_215[7:6] == 2'h1 ? _GEN_273 : valid_1_9; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_834 = _GEN_215[7:6] == 2'h1 ? _GEN_274 : valid_1_10; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_835 = _GEN_215[7:6] == 2'h1 ? _GEN_275 : valid_1_11; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_836 = _GEN_215[7:6] == 2'h1 ? _GEN_276 : valid_1_12; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_837 = _GEN_215[7:6] == 2'h1 ? _GEN_277 : valid_1_13; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_838 = _GEN_215[7:6] == 2'h1 ? _GEN_278 : valid_1_14; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_839 = _GEN_215[7:6] == 2'h1 ? _GEN_279 : valid_1_15; // @[i_cache.scala 111:52 28:26]
  wire [7:0] _GEN_840 = _GEN_215[7:6] == 2'h1 ? _GEN_280 : _GEN_728; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_841 = _GEN_215[7:6] == 2'h1 ? _GEN_281 : _GEN_729; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_842 = _GEN_215[7:6] == 2'h1 ? _GEN_282 : _GEN_730; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_843 = _GEN_215[7:6] == 2'h1 ? _GEN_283 : _GEN_731; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_844 = _GEN_215[7:6] == 2'h1 ? _GEN_284 : _GEN_732; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_845 = _GEN_215[7:6] == 2'h1 ? _GEN_285 : _GEN_733; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_846 = _GEN_215[7:6] == 2'h1 ? _GEN_286 : _GEN_734; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_847 = _GEN_215[7:6] == 2'h1 ? _GEN_287 : _GEN_735; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_848 = _GEN_215[7:6] == 2'h1 ? _GEN_288 : _GEN_736; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_849 = _GEN_215[7:6] == 2'h1 ? _GEN_289 : _GEN_737; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_850 = _GEN_215[7:6] == 2'h1 ? _GEN_290 : _GEN_738; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_851 = _GEN_215[7:6] == 2'h1 ? _GEN_291 : _GEN_739; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_852 = _GEN_215[7:6] == 2'h1 ? _GEN_292 : _GEN_740; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_853 = _GEN_215[7:6] == 2'h1 ? _GEN_293 : _GEN_741; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_854 = _GEN_215[7:6] == 2'h1 ? _GEN_294 : _GEN_742; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_855 = _GEN_215[7:6] == 2'h1 ? _GEN_295 : _GEN_743; // @[i_cache.scala 111:52]
  wire [511:0] _GEN_856 = _GEN_215[7:6] == 2'h1 ? ram_2_0 : _GEN_680; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_857 = _GEN_215[7:6] == 2'h1 ? ram_2_1 : _GEN_681; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_858 = _GEN_215[7:6] == 2'h1 ? ram_2_2 : _GEN_682; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_859 = _GEN_215[7:6] == 2'h1 ? ram_2_3 : _GEN_683; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_860 = _GEN_215[7:6] == 2'h1 ? ram_2_4 : _GEN_684; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_861 = _GEN_215[7:6] == 2'h1 ? ram_2_5 : _GEN_685; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_862 = _GEN_215[7:6] == 2'h1 ? ram_2_6 : _GEN_686; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_863 = _GEN_215[7:6] == 2'h1 ? ram_2_7 : _GEN_687; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_864 = _GEN_215[7:6] == 2'h1 ? ram_2_8 : _GEN_688; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_865 = _GEN_215[7:6] == 2'h1 ? ram_2_9 : _GEN_689; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_866 = _GEN_215[7:6] == 2'h1 ? ram_2_10 : _GEN_690; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_867 = _GEN_215[7:6] == 2'h1 ? ram_2_11 : _GEN_691; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_868 = _GEN_215[7:6] == 2'h1 ? ram_2_12 : _GEN_692; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_869 = _GEN_215[7:6] == 2'h1 ? ram_2_13 : _GEN_693; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_870 = _GEN_215[7:6] == 2'h1 ? ram_2_14 : _GEN_694; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_871 = _GEN_215[7:6] == 2'h1 ? ram_2_15 : _GEN_695; // @[i_cache.scala 111:52 21:24]
  wire [31:0] _GEN_872 = _GEN_215[7:6] == 2'h1 ? tag_2_0 : _GEN_696; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_873 = _GEN_215[7:6] == 2'h1 ? tag_2_1 : _GEN_697; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_874 = _GEN_215[7:6] == 2'h1 ? tag_2_2 : _GEN_698; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_875 = _GEN_215[7:6] == 2'h1 ? tag_2_3 : _GEN_699; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_876 = _GEN_215[7:6] == 2'h1 ? tag_2_4 : _GEN_700; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_877 = _GEN_215[7:6] == 2'h1 ? tag_2_5 : _GEN_701; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_878 = _GEN_215[7:6] == 2'h1 ? tag_2_6 : _GEN_702; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_879 = _GEN_215[7:6] == 2'h1 ? tag_2_7 : _GEN_703; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_880 = _GEN_215[7:6] == 2'h1 ? tag_2_8 : _GEN_704; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_881 = _GEN_215[7:6] == 2'h1 ? tag_2_9 : _GEN_705; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_882 = _GEN_215[7:6] == 2'h1 ? tag_2_10 : _GEN_706; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_883 = _GEN_215[7:6] == 2'h1 ? tag_2_11 : _GEN_707; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_884 = _GEN_215[7:6] == 2'h1 ? tag_2_12 : _GEN_708; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_885 = _GEN_215[7:6] == 2'h1 ? tag_2_13 : _GEN_709; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_886 = _GEN_215[7:6] == 2'h1 ? tag_2_14 : _GEN_710; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_887 = _GEN_215[7:6] == 2'h1 ? tag_2_15 : _GEN_711; // @[i_cache.scala 111:52 25:24]
  wire  _GEN_888 = _GEN_215[7:6] == 2'h1 ? valid_2_0 : _GEN_712; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_889 = _GEN_215[7:6] == 2'h1 ? valid_2_1 : _GEN_713; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_890 = _GEN_215[7:6] == 2'h1 ? valid_2_2 : _GEN_714; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_891 = _GEN_215[7:6] == 2'h1 ? valid_2_3 : _GEN_715; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_892 = _GEN_215[7:6] == 2'h1 ? valid_2_4 : _GEN_716; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_893 = _GEN_215[7:6] == 2'h1 ? valid_2_5 : _GEN_717; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_894 = _GEN_215[7:6] == 2'h1 ? valid_2_6 : _GEN_718; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_895 = _GEN_215[7:6] == 2'h1 ? valid_2_7 : _GEN_719; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_896 = _GEN_215[7:6] == 2'h1 ? valid_2_8 : _GEN_720; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_897 = _GEN_215[7:6] == 2'h1 ? valid_2_9 : _GEN_721; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_898 = _GEN_215[7:6] == 2'h1 ? valid_2_10 : _GEN_722; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_899 = _GEN_215[7:6] == 2'h1 ? valid_2_11 : _GEN_723; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_900 = _GEN_215[7:6] == 2'h1 ? valid_2_12 : _GEN_724; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_901 = _GEN_215[7:6] == 2'h1 ? valid_2_13 : _GEN_725; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_902 = _GEN_215[7:6] == 2'h1 ? valid_2_14 : _GEN_726; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_903 = _GEN_215[7:6] == 2'h1 ? valid_2_15 : _GEN_727; // @[i_cache.scala 111:52 29:26]
  wire [511:0] _GEN_904 = _GEN_215[7:6] == 2'h1 ? ram_3_0 : _GEN_744; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_905 = _GEN_215[7:6] == 2'h1 ? ram_3_1 : _GEN_745; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_906 = _GEN_215[7:6] == 2'h1 ? ram_3_2 : _GEN_746; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_907 = _GEN_215[7:6] == 2'h1 ? ram_3_3 : _GEN_747; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_908 = _GEN_215[7:6] == 2'h1 ? ram_3_4 : _GEN_748; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_909 = _GEN_215[7:6] == 2'h1 ? ram_3_5 : _GEN_749; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_910 = _GEN_215[7:6] == 2'h1 ? ram_3_6 : _GEN_750; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_911 = _GEN_215[7:6] == 2'h1 ? ram_3_7 : _GEN_751; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_912 = _GEN_215[7:6] == 2'h1 ? ram_3_8 : _GEN_752; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_913 = _GEN_215[7:6] == 2'h1 ? ram_3_9 : _GEN_753; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_914 = _GEN_215[7:6] == 2'h1 ? ram_3_10 : _GEN_754; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_915 = _GEN_215[7:6] == 2'h1 ? ram_3_11 : _GEN_755; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_916 = _GEN_215[7:6] == 2'h1 ? ram_3_12 : _GEN_756; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_917 = _GEN_215[7:6] == 2'h1 ? ram_3_13 : _GEN_757; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_918 = _GEN_215[7:6] == 2'h1 ? ram_3_14 : _GEN_758; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_919 = _GEN_215[7:6] == 2'h1 ? ram_3_15 : _GEN_759; // @[i_cache.scala 111:52 22:24]
  wire [31:0] _GEN_920 = _GEN_215[7:6] == 2'h1 ? tag_3_0 : _GEN_760; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_921 = _GEN_215[7:6] == 2'h1 ? tag_3_1 : _GEN_761; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_922 = _GEN_215[7:6] == 2'h1 ? tag_3_2 : _GEN_762; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_923 = _GEN_215[7:6] == 2'h1 ? tag_3_3 : _GEN_763; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_924 = _GEN_215[7:6] == 2'h1 ? tag_3_4 : _GEN_764; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_925 = _GEN_215[7:6] == 2'h1 ? tag_3_5 : _GEN_765; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_926 = _GEN_215[7:6] == 2'h1 ? tag_3_6 : _GEN_766; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_927 = _GEN_215[7:6] == 2'h1 ? tag_3_7 : _GEN_767; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_928 = _GEN_215[7:6] == 2'h1 ? tag_3_8 : _GEN_768; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_929 = _GEN_215[7:6] == 2'h1 ? tag_3_9 : _GEN_769; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_930 = _GEN_215[7:6] == 2'h1 ? tag_3_10 : _GEN_770; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_931 = _GEN_215[7:6] == 2'h1 ? tag_3_11 : _GEN_771; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_932 = _GEN_215[7:6] == 2'h1 ? tag_3_12 : _GEN_772; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_933 = _GEN_215[7:6] == 2'h1 ? tag_3_13 : _GEN_773; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_934 = _GEN_215[7:6] == 2'h1 ? tag_3_14 : _GEN_774; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_935 = _GEN_215[7:6] == 2'h1 ? tag_3_15 : _GEN_775; // @[i_cache.scala 111:52 26:24]
  wire  _GEN_936 = _GEN_215[7:6] == 2'h1 ? valid_3_0 : _GEN_776; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_937 = _GEN_215[7:6] == 2'h1 ? valid_3_1 : _GEN_777; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_938 = _GEN_215[7:6] == 2'h1 ? valid_3_2 : _GEN_778; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_939 = _GEN_215[7:6] == 2'h1 ? valid_3_3 : _GEN_779; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_940 = _GEN_215[7:6] == 2'h1 ? valid_3_4 : _GEN_780; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_941 = _GEN_215[7:6] == 2'h1 ? valid_3_5 : _GEN_781; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_942 = _GEN_215[7:6] == 2'h1 ? valid_3_6 : _GEN_782; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_943 = _GEN_215[7:6] == 2'h1 ? valid_3_7 : _GEN_783; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_944 = _GEN_215[7:6] == 2'h1 ? valid_3_8 : _GEN_784; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_945 = _GEN_215[7:6] == 2'h1 ? valid_3_9 : _GEN_785; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_946 = _GEN_215[7:6] == 2'h1 ? valid_3_10 : _GEN_786; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_947 = _GEN_215[7:6] == 2'h1 ? valid_3_11 : _GEN_787; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_948 = _GEN_215[7:6] == 2'h1 ? valid_3_12 : _GEN_788; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_949 = _GEN_215[7:6] == 2'h1 ? valid_3_13 : _GEN_789; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_950 = _GEN_215[7:6] == 2'h1 ? valid_3_14 : _GEN_790; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_951 = _GEN_215[7:6] == 2'h1 ? valid_3_15 : _GEN_791; // @[i_cache.scala 111:52 30:26]
  wire [511:0] _GEN_952 = _GEN_215[7:6] == 2'h0 ? _GEN_152 : ram_0_0; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_953 = _GEN_215[7:6] == 2'h0 ? _GEN_153 : ram_0_1; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_954 = _GEN_215[7:6] == 2'h0 ? _GEN_154 : ram_0_2; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_955 = _GEN_215[7:6] == 2'h0 ? _GEN_155 : ram_0_3; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_956 = _GEN_215[7:6] == 2'h0 ? _GEN_156 : ram_0_4; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_957 = _GEN_215[7:6] == 2'h0 ? _GEN_157 : ram_0_5; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_958 = _GEN_215[7:6] == 2'h0 ? _GEN_158 : ram_0_6; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_959 = _GEN_215[7:6] == 2'h0 ? _GEN_159 : ram_0_7; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_960 = _GEN_215[7:6] == 2'h0 ? _GEN_160 : ram_0_8; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_961 = _GEN_215[7:6] == 2'h0 ? _GEN_161 : ram_0_9; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_962 = _GEN_215[7:6] == 2'h0 ? _GEN_162 : ram_0_10; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_963 = _GEN_215[7:6] == 2'h0 ? _GEN_163 : ram_0_11; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_964 = _GEN_215[7:6] == 2'h0 ? _GEN_164 : ram_0_12; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_965 = _GEN_215[7:6] == 2'h0 ? _GEN_165 : ram_0_13; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_966 = _GEN_215[7:6] == 2'h0 ? _GEN_166 : ram_0_14; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_967 = _GEN_215[7:6] == 2'h0 ? _GEN_167 : ram_0_15; // @[i_cache.scala 106:46 19:24]
  wire [31:0] _GEN_968 = _GEN_215[7:6] == 2'h0 ? _GEN_168 : tag_0_0; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_969 = _GEN_215[7:6] == 2'h0 ? _GEN_169 : tag_0_1; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_970 = _GEN_215[7:6] == 2'h0 ? _GEN_170 : tag_0_2; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_971 = _GEN_215[7:6] == 2'h0 ? _GEN_171 : tag_0_3; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_972 = _GEN_215[7:6] == 2'h0 ? _GEN_172 : tag_0_4; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_973 = _GEN_215[7:6] == 2'h0 ? _GEN_173 : tag_0_5; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_974 = _GEN_215[7:6] == 2'h0 ? _GEN_174 : tag_0_6; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_975 = _GEN_215[7:6] == 2'h0 ? _GEN_175 : tag_0_7; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_976 = _GEN_215[7:6] == 2'h0 ? _GEN_176 : tag_0_8; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_977 = _GEN_215[7:6] == 2'h0 ? _GEN_177 : tag_0_9; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_978 = _GEN_215[7:6] == 2'h0 ? _GEN_178 : tag_0_10; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_979 = _GEN_215[7:6] == 2'h0 ? _GEN_179 : tag_0_11; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_980 = _GEN_215[7:6] == 2'h0 ? _GEN_180 : tag_0_12; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_981 = _GEN_215[7:6] == 2'h0 ? _GEN_181 : tag_0_13; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_982 = _GEN_215[7:6] == 2'h0 ? _GEN_182 : tag_0_14; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_983 = _GEN_215[7:6] == 2'h0 ? _GEN_183 : tag_0_15; // @[i_cache.scala 106:46 23:24]
  wire  _GEN_984 = _GEN_215[7:6] == 2'h0 ? _GEN_184 : valid_0_0; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_985 = _GEN_215[7:6] == 2'h0 ? _GEN_185 : valid_0_1; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_986 = _GEN_215[7:6] == 2'h0 ? _GEN_186 : valid_0_2; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_987 = _GEN_215[7:6] == 2'h0 ? _GEN_187 : valid_0_3; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_988 = _GEN_215[7:6] == 2'h0 ? _GEN_188 : valid_0_4; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_989 = _GEN_215[7:6] == 2'h0 ? _GEN_189 : valid_0_5; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_990 = _GEN_215[7:6] == 2'h0 ? _GEN_190 : valid_0_6; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_991 = _GEN_215[7:6] == 2'h0 ? _GEN_191 : valid_0_7; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_992 = _GEN_215[7:6] == 2'h0 ? _GEN_192 : valid_0_8; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_993 = _GEN_215[7:6] == 2'h0 ? _GEN_193 : valid_0_9; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_994 = _GEN_215[7:6] == 2'h0 ? _GEN_194 : valid_0_10; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_995 = _GEN_215[7:6] == 2'h0 ? _GEN_195 : valid_0_11; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_996 = _GEN_215[7:6] == 2'h0 ? _GEN_196 : valid_0_12; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_997 = _GEN_215[7:6] == 2'h0 ? _GEN_197 : valid_0_13; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_998 = _GEN_215[7:6] == 2'h0 ? _GEN_198 : valid_0_14; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_999 = _GEN_215[7:6] == 2'h0 ? _GEN_199 : valid_0_15; // @[i_cache.scala 106:46 27:26]
  wire [7:0] _GEN_1000 = _GEN_215[7:6] == 2'h0 ? _GEN_216 : _GEN_840; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1001 = _GEN_215[7:6] == 2'h0 ? _GEN_217 : _GEN_841; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1002 = _GEN_215[7:6] == 2'h0 ? _GEN_218 : _GEN_842; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1003 = _GEN_215[7:6] == 2'h0 ? _GEN_219 : _GEN_843; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1004 = _GEN_215[7:6] == 2'h0 ? _GEN_220 : _GEN_844; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1005 = _GEN_215[7:6] == 2'h0 ? _GEN_221 : _GEN_845; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1006 = _GEN_215[7:6] == 2'h0 ? _GEN_222 : _GEN_846; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1007 = _GEN_215[7:6] == 2'h0 ? _GEN_223 : _GEN_847; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1008 = _GEN_215[7:6] == 2'h0 ? _GEN_224 : _GEN_848; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1009 = _GEN_215[7:6] == 2'h0 ? _GEN_225 : _GEN_849; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1010 = _GEN_215[7:6] == 2'h0 ? _GEN_226 : _GEN_850; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1011 = _GEN_215[7:6] == 2'h0 ? _GEN_227 : _GEN_851; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1012 = _GEN_215[7:6] == 2'h0 ? _GEN_228 : _GEN_852; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1013 = _GEN_215[7:6] == 2'h0 ? _GEN_229 : _GEN_853; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1014 = _GEN_215[7:6] == 2'h0 ? _GEN_230 : _GEN_854; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1015 = _GEN_215[7:6] == 2'h0 ? _GEN_231 : _GEN_855; // @[i_cache.scala 106:46]
  wire [511:0] _GEN_1016 = _GEN_215[7:6] == 2'h0 ? ram_1_0 : _GEN_792; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1017 = _GEN_215[7:6] == 2'h0 ? ram_1_1 : _GEN_793; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1018 = _GEN_215[7:6] == 2'h0 ? ram_1_2 : _GEN_794; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1019 = _GEN_215[7:6] == 2'h0 ? ram_1_3 : _GEN_795; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1020 = _GEN_215[7:6] == 2'h0 ? ram_1_4 : _GEN_796; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1021 = _GEN_215[7:6] == 2'h0 ? ram_1_5 : _GEN_797; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1022 = _GEN_215[7:6] == 2'h0 ? ram_1_6 : _GEN_798; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1023 = _GEN_215[7:6] == 2'h0 ? ram_1_7 : _GEN_799; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1024 = _GEN_215[7:6] == 2'h0 ? ram_1_8 : _GEN_800; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1025 = _GEN_215[7:6] == 2'h0 ? ram_1_9 : _GEN_801; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1026 = _GEN_215[7:6] == 2'h0 ? ram_1_10 : _GEN_802; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1027 = _GEN_215[7:6] == 2'h0 ? ram_1_11 : _GEN_803; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1028 = _GEN_215[7:6] == 2'h0 ? ram_1_12 : _GEN_804; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1029 = _GEN_215[7:6] == 2'h0 ? ram_1_13 : _GEN_805; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1030 = _GEN_215[7:6] == 2'h0 ? ram_1_14 : _GEN_806; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1031 = _GEN_215[7:6] == 2'h0 ? ram_1_15 : _GEN_807; // @[i_cache.scala 106:46 20:24]
  wire [31:0] _GEN_1032 = _GEN_215[7:6] == 2'h0 ? tag_1_0 : _GEN_808; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1033 = _GEN_215[7:6] == 2'h0 ? tag_1_1 : _GEN_809; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1034 = _GEN_215[7:6] == 2'h0 ? tag_1_2 : _GEN_810; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1035 = _GEN_215[7:6] == 2'h0 ? tag_1_3 : _GEN_811; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1036 = _GEN_215[7:6] == 2'h0 ? tag_1_4 : _GEN_812; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1037 = _GEN_215[7:6] == 2'h0 ? tag_1_5 : _GEN_813; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1038 = _GEN_215[7:6] == 2'h0 ? tag_1_6 : _GEN_814; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1039 = _GEN_215[7:6] == 2'h0 ? tag_1_7 : _GEN_815; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1040 = _GEN_215[7:6] == 2'h0 ? tag_1_8 : _GEN_816; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1041 = _GEN_215[7:6] == 2'h0 ? tag_1_9 : _GEN_817; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1042 = _GEN_215[7:6] == 2'h0 ? tag_1_10 : _GEN_818; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1043 = _GEN_215[7:6] == 2'h0 ? tag_1_11 : _GEN_819; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1044 = _GEN_215[7:6] == 2'h0 ? tag_1_12 : _GEN_820; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1045 = _GEN_215[7:6] == 2'h0 ? tag_1_13 : _GEN_821; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1046 = _GEN_215[7:6] == 2'h0 ? tag_1_14 : _GEN_822; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1047 = _GEN_215[7:6] == 2'h0 ? tag_1_15 : _GEN_823; // @[i_cache.scala 106:46 24:24]
  wire  _GEN_1048 = _GEN_215[7:6] == 2'h0 ? valid_1_0 : _GEN_824; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1049 = _GEN_215[7:6] == 2'h0 ? valid_1_1 : _GEN_825; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1050 = _GEN_215[7:6] == 2'h0 ? valid_1_2 : _GEN_826; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1051 = _GEN_215[7:6] == 2'h0 ? valid_1_3 : _GEN_827; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1052 = _GEN_215[7:6] == 2'h0 ? valid_1_4 : _GEN_828; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1053 = _GEN_215[7:6] == 2'h0 ? valid_1_5 : _GEN_829; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1054 = _GEN_215[7:6] == 2'h0 ? valid_1_6 : _GEN_830; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1055 = _GEN_215[7:6] == 2'h0 ? valid_1_7 : _GEN_831; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1056 = _GEN_215[7:6] == 2'h0 ? valid_1_8 : _GEN_832; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1057 = _GEN_215[7:6] == 2'h0 ? valid_1_9 : _GEN_833; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1058 = _GEN_215[7:6] == 2'h0 ? valid_1_10 : _GEN_834; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1059 = _GEN_215[7:6] == 2'h0 ? valid_1_11 : _GEN_835; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1060 = _GEN_215[7:6] == 2'h0 ? valid_1_12 : _GEN_836; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1061 = _GEN_215[7:6] == 2'h0 ? valid_1_13 : _GEN_837; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1062 = _GEN_215[7:6] == 2'h0 ? valid_1_14 : _GEN_838; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1063 = _GEN_215[7:6] == 2'h0 ? valid_1_15 : _GEN_839; // @[i_cache.scala 106:46 28:26]
  wire [511:0] _GEN_1064 = _GEN_215[7:6] == 2'h0 ? ram_2_0 : _GEN_856; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1065 = _GEN_215[7:6] == 2'h0 ? ram_2_1 : _GEN_857; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1066 = _GEN_215[7:6] == 2'h0 ? ram_2_2 : _GEN_858; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1067 = _GEN_215[7:6] == 2'h0 ? ram_2_3 : _GEN_859; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1068 = _GEN_215[7:6] == 2'h0 ? ram_2_4 : _GEN_860; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1069 = _GEN_215[7:6] == 2'h0 ? ram_2_5 : _GEN_861; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1070 = _GEN_215[7:6] == 2'h0 ? ram_2_6 : _GEN_862; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1071 = _GEN_215[7:6] == 2'h0 ? ram_2_7 : _GEN_863; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1072 = _GEN_215[7:6] == 2'h0 ? ram_2_8 : _GEN_864; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1073 = _GEN_215[7:6] == 2'h0 ? ram_2_9 : _GEN_865; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1074 = _GEN_215[7:6] == 2'h0 ? ram_2_10 : _GEN_866; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1075 = _GEN_215[7:6] == 2'h0 ? ram_2_11 : _GEN_867; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1076 = _GEN_215[7:6] == 2'h0 ? ram_2_12 : _GEN_868; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1077 = _GEN_215[7:6] == 2'h0 ? ram_2_13 : _GEN_869; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1078 = _GEN_215[7:6] == 2'h0 ? ram_2_14 : _GEN_870; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1079 = _GEN_215[7:6] == 2'h0 ? ram_2_15 : _GEN_871; // @[i_cache.scala 106:46 21:24]
  wire [31:0] _GEN_1080 = _GEN_215[7:6] == 2'h0 ? tag_2_0 : _GEN_872; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1081 = _GEN_215[7:6] == 2'h0 ? tag_2_1 : _GEN_873; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1082 = _GEN_215[7:6] == 2'h0 ? tag_2_2 : _GEN_874; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1083 = _GEN_215[7:6] == 2'h0 ? tag_2_3 : _GEN_875; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1084 = _GEN_215[7:6] == 2'h0 ? tag_2_4 : _GEN_876; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1085 = _GEN_215[7:6] == 2'h0 ? tag_2_5 : _GEN_877; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1086 = _GEN_215[7:6] == 2'h0 ? tag_2_6 : _GEN_878; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1087 = _GEN_215[7:6] == 2'h0 ? tag_2_7 : _GEN_879; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1088 = _GEN_215[7:6] == 2'h0 ? tag_2_8 : _GEN_880; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1089 = _GEN_215[7:6] == 2'h0 ? tag_2_9 : _GEN_881; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1090 = _GEN_215[7:6] == 2'h0 ? tag_2_10 : _GEN_882; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1091 = _GEN_215[7:6] == 2'h0 ? tag_2_11 : _GEN_883; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1092 = _GEN_215[7:6] == 2'h0 ? tag_2_12 : _GEN_884; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1093 = _GEN_215[7:6] == 2'h0 ? tag_2_13 : _GEN_885; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1094 = _GEN_215[7:6] == 2'h0 ? tag_2_14 : _GEN_886; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1095 = _GEN_215[7:6] == 2'h0 ? tag_2_15 : _GEN_887; // @[i_cache.scala 106:46 25:24]
  wire  _GEN_1096 = _GEN_215[7:6] == 2'h0 ? valid_2_0 : _GEN_888; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1097 = _GEN_215[7:6] == 2'h0 ? valid_2_1 : _GEN_889; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1098 = _GEN_215[7:6] == 2'h0 ? valid_2_2 : _GEN_890; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1099 = _GEN_215[7:6] == 2'h0 ? valid_2_3 : _GEN_891; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1100 = _GEN_215[7:6] == 2'h0 ? valid_2_4 : _GEN_892; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1101 = _GEN_215[7:6] == 2'h0 ? valid_2_5 : _GEN_893; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1102 = _GEN_215[7:6] == 2'h0 ? valid_2_6 : _GEN_894; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1103 = _GEN_215[7:6] == 2'h0 ? valid_2_7 : _GEN_895; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1104 = _GEN_215[7:6] == 2'h0 ? valid_2_8 : _GEN_896; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1105 = _GEN_215[7:6] == 2'h0 ? valid_2_9 : _GEN_897; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1106 = _GEN_215[7:6] == 2'h0 ? valid_2_10 : _GEN_898; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1107 = _GEN_215[7:6] == 2'h0 ? valid_2_11 : _GEN_899; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1108 = _GEN_215[7:6] == 2'h0 ? valid_2_12 : _GEN_900; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1109 = _GEN_215[7:6] == 2'h0 ? valid_2_13 : _GEN_901; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1110 = _GEN_215[7:6] == 2'h0 ? valid_2_14 : _GEN_902; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1111 = _GEN_215[7:6] == 2'h0 ? valid_2_15 : _GEN_903; // @[i_cache.scala 106:46 29:26]
  wire [511:0] _GEN_1112 = _GEN_215[7:6] == 2'h0 ? ram_3_0 : _GEN_904; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1113 = _GEN_215[7:6] == 2'h0 ? ram_3_1 : _GEN_905; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1114 = _GEN_215[7:6] == 2'h0 ? ram_3_2 : _GEN_906; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1115 = _GEN_215[7:6] == 2'h0 ? ram_3_3 : _GEN_907; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1116 = _GEN_215[7:6] == 2'h0 ? ram_3_4 : _GEN_908; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1117 = _GEN_215[7:6] == 2'h0 ? ram_3_5 : _GEN_909; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1118 = _GEN_215[7:6] == 2'h0 ? ram_3_6 : _GEN_910; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1119 = _GEN_215[7:6] == 2'h0 ? ram_3_7 : _GEN_911; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1120 = _GEN_215[7:6] == 2'h0 ? ram_3_8 : _GEN_912; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1121 = _GEN_215[7:6] == 2'h0 ? ram_3_9 : _GEN_913; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1122 = _GEN_215[7:6] == 2'h0 ? ram_3_10 : _GEN_914; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1123 = _GEN_215[7:6] == 2'h0 ? ram_3_11 : _GEN_915; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1124 = _GEN_215[7:6] == 2'h0 ? ram_3_12 : _GEN_916; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1125 = _GEN_215[7:6] == 2'h0 ? ram_3_13 : _GEN_917; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1126 = _GEN_215[7:6] == 2'h0 ? ram_3_14 : _GEN_918; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1127 = _GEN_215[7:6] == 2'h0 ? ram_3_15 : _GEN_919; // @[i_cache.scala 106:46 22:24]
  wire [31:0] _GEN_1128 = _GEN_215[7:6] == 2'h0 ? tag_3_0 : _GEN_920; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1129 = _GEN_215[7:6] == 2'h0 ? tag_3_1 : _GEN_921; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1130 = _GEN_215[7:6] == 2'h0 ? tag_3_2 : _GEN_922; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1131 = _GEN_215[7:6] == 2'h0 ? tag_3_3 : _GEN_923; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1132 = _GEN_215[7:6] == 2'h0 ? tag_3_4 : _GEN_924; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1133 = _GEN_215[7:6] == 2'h0 ? tag_3_5 : _GEN_925; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1134 = _GEN_215[7:6] == 2'h0 ? tag_3_6 : _GEN_926; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1135 = _GEN_215[7:6] == 2'h0 ? tag_3_7 : _GEN_927; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1136 = _GEN_215[7:6] == 2'h0 ? tag_3_8 : _GEN_928; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1137 = _GEN_215[7:6] == 2'h0 ? tag_3_9 : _GEN_929; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1138 = _GEN_215[7:6] == 2'h0 ? tag_3_10 : _GEN_930; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1139 = _GEN_215[7:6] == 2'h0 ? tag_3_11 : _GEN_931; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1140 = _GEN_215[7:6] == 2'h0 ? tag_3_12 : _GEN_932; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1141 = _GEN_215[7:6] == 2'h0 ? tag_3_13 : _GEN_933; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1142 = _GEN_215[7:6] == 2'h0 ? tag_3_14 : _GEN_934; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1143 = _GEN_215[7:6] == 2'h0 ? tag_3_15 : _GEN_935; // @[i_cache.scala 106:46 26:24]
  wire  _GEN_1144 = _GEN_215[7:6] == 2'h0 ? valid_3_0 : _GEN_936; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1145 = _GEN_215[7:6] == 2'h0 ? valid_3_1 : _GEN_937; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1146 = _GEN_215[7:6] == 2'h0 ? valid_3_2 : _GEN_938; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1147 = _GEN_215[7:6] == 2'h0 ? valid_3_3 : _GEN_939; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1148 = _GEN_215[7:6] == 2'h0 ? valid_3_4 : _GEN_940; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1149 = _GEN_215[7:6] == 2'h0 ? valid_3_5 : _GEN_941; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1150 = _GEN_215[7:6] == 2'h0 ? valid_3_6 : _GEN_942; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1151 = _GEN_215[7:6] == 2'h0 ? valid_3_7 : _GEN_943; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1152 = _GEN_215[7:6] == 2'h0 ? valid_3_8 : _GEN_944; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1153 = _GEN_215[7:6] == 2'h0 ? valid_3_9 : _GEN_945; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1154 = _GEN_215[7:6] == 2'h0 ? valid_3_10 : _GEN_946; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1155 = _GEN_215[7:6] == 2'h0 ? valid_3_11 : _GEN_947; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1156 = _GEN_215[7:6] == 2'h0 ? valid_3_12 : _GEN_948; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1157 = _GEN_215[7:6] == 2'h0 ? valid_3_13 : _GEN_949; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1158 = _GEN_215[7:6] == 2'h0 ? valid_3_14 : _GEN_950; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1159 = _GEN_215[7:6] == 2'h0 ? valid_3_15 : _GEN_951; // @[i_cache.scala 106:46 30:26]
  wire [511:0] _GEN_1160 = unuse_way == 3'h4 ? _GEN_360 : _GEN_1112; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1161 = unuse_way == 3'h4 ? _GEN_361 : _GEN_1113; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1162 = unuse_way == 3'h4 ? _GEN_362 : _GEN_1114; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1163 = unuse_way == 3'h4 ? _GEN_363 : _GEN_1115; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1164 = unuse_way == 3'h4 ? _GEN_364 : _GEN_1116; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1165 = unuse_way == 3'h4 ? _GEN_365 : _GEN_1117; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1166 = unuse_way == 3'h4 ? _GEN_366 : _GEN_1118; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1167 = unuse_way == 3'h4 ? _GEN_367 : _GEN_1119; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1168 = unuse_way == 3'h4 ? _GEN_368 : _GEN_1120; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1169 = unuse_way == 3'h4 ? _GEN_369 : _GEN_1121; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1170 = unuse_way == 3'h4 ? _GEN_370 : _GEN_1122; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1171 = unuse_way == 3'h4 ? _GEN_371 : _GEN_1123; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1172 = unuse_way == 3'h4 ? _GEN_372 : _GEN_1124; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1173 = unuse_way == 3'h4 ? _GEN_373 : _GEN_1125; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1174 = unuse_way == 3'h4 ? _GEN_374 : _GEN_1126; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1175 = unuse_way == 3'h4 ? _GEN_375 : _GEN_1127; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1176 = unuse_way == 3'h4 ? _GEN_376 : _GEN_1128; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1177 = unuse_way == 3'h4 ? _GEN_377 : _GEN_1129; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1178 = unuse_way == 3'h4 ? _GEN_378 : _GEN_1130; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1179 = unuse_way == 3'h4 ? _GEN_379 : _GEN_1131; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1180 = unuse_way == 3'h4 ? _GEN_380 : _GEN_1132; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1181 = unuse_way == 3'h4 ? _GEN_381 : _GEN_1133; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1182 = unuse_way == 3'h4 ? _GEN_382 : _GEN_1134; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1183 = unuse_way == 3'h4 ? _GEN_383 : _GEN_1135; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1184 = unuse_way == 3'h4 ? _GEN_384 : _GEN_1136; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1185 = unuse_way == 3'h4 ? _GEN_385 : _GEN_1137; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1186 = unuse_way == 3'h4 ? _GEN_386 : _GEN_1138; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1187 = unuse_way == 3'h4 ? _GEN_387 : _GEN_1139; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1188 = unuse_way == 3'h4 ? _GEN_388 : _GEN_1140; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1189 = unuse_way == 3'h4 ? _GEN_389 : _GEN_1141; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1190 = unuse_way == 3'h4 ? _GEN_390 : _GEN_1142; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1191 = unuse_way == 3'h4 ? _GEN_391 : _GEN_1143; // @[i_cache.scala 100:40]
  wire  _GEN_1192 = unuse_way == 3'h4 ? _GEN_392 : _GEN_1144; // @[i_cache.scala 100:40]
  wire  _GEN_1193 = unuse_way == 3'h4 ? _GEN_393 : _GEN_1145; // @[i_cache.scala 100:40]
  wire  _GEN_1194 = unuse_way == 3'h4 ? _GEN_394 : _GEN_1146; // @[i_cache.scala 100:40]
  wire  _GEN_1195 = unuse_way == 3'h4 ? _GEN_395 : _GEN_1147; // @[i_cache.scala 100:40]
  wire  _GEN_1196 = unuse_way == 3'h4 ? _GEN_396 : _GEN_1148; // @[i_cache.scala 100:40]
  wire  _GEN_1197 = unuse_way == 3'h4 ? _GEN_397 : _GEN_1149; // @[i_cache.scala 100:40]
  wire  _GEN_1198 = unuse_way == 3'h4 ? _GEN_398 : _GEN_1150; // @[i_cache.scala 100:40]
  wire  _GEN_1199 = unuse_way == 3'h4 ? _GEN_399 : _GEN_1151; // @[i_cache.scala 100:40]
  wire  _GEN_1200 = unuse_way == 3'h4 ? _GEN_400 : _GEN_1152; // @[i_cache.scala 100:40]
  wire  _GEN_1201 = unuse_way == 3'h4 ? _GEN_401 : _GEN_1153; // @[i_cache.scala 100:40]
  wire  _GEN_1202 = unuse_way == 3'h4 ? _GEN_402 : _GEN_1154; // @[i_cache.scala 100:40]
  wire  _GEN_1203 = unuse_way == 3'h4 ? _GEN_403 : _GEN_1155; // @[i_cache.scala 100:40]
  wire  _GEN_1204 = unuse_way == 3'h4 ? _GEN_404 : _GEN_1156; // @[i_cache.scala 100:40]
  wire  _GEN_1205 = unuse_way == 3'h4 ? _GEN_405 : _GEN_1157; // @[i_cache.scala 100:40]
  wire  _GEN_1206 = unuse_way == 3'h4 ? _GEN_406 : _GEN_1158; // @[i_cache.scala 100:40]
  wire  _GEN_1207 = unuse_way == 3'h4 ? _GEN_407 : _GEN_1159; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1208 = unuse_way == 3'h4 ? _GEN_408 : _GEN_1000; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1209 = unuse_way == 3'h4 ? _GEN_409 : _GEN_1001; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1210 = unuse_way == 3'h4 ? _GEN_410 : _GEN_1002; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1211 = unuse_way == 3'h4 ? _GEN_411 : _GEN_1003; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1212 = unuse_way == 3'h4 ? _GEN_412 : _GEN_1004; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1213 = unuse_way == 3'h4 ? _GEN_413 : _GEN_1005; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1214 = unuse_way == 3'h4 ? _GEN_414 : _GEN_1006; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1215 = unuse_way == 3'h4 ? _GEN_415 : _GEN_1007; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1216 = unuse_way == 3'h4 ? _GEN_416 : _GEN_1008; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1217 = unuse_way == 3'h4 ? _GEN_417 : _GEN_1009; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1218 = unuse_way == 3'h4 ? _GEN_418 : _GEN_1010; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1219 = unuse_way == 3'h4 ? _GEN_419 : _GEN_1011; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1220 = unuse_way == 3'h4 ? _GEN_420 : _GEN_1012; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1221 = unuse_way == 3'h4 ? _GEN_421 : _GEN_1013; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1222 = unuse_way == 3'h4 ? _GEN_422 : _GEN_1014; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1223 = unuse_way == 3'h4 ? _GEN_423 : _GEN_1015; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1224 = unuse_way == 3'h4 ? ram_0_0 : _GEN_952; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1225 = unuse_way == 3'h4 ? ram_0_1 : _GEN_953; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1226 = unuse_way == 3'h4 ? ram_0_2 : _GEN_954; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1227 = unuse_way == 3'h4 ? ram_0_3 : _GEN_955; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1228 = unuse_way == 3'h4 ? ram_0_4 : _GEN_956; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1229 = unuse_way == 3'h4 ? ram_0_5 : _GEN_957; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1230 = unuse_way == 3'h4 ? ram_0_6 : _GEN_958; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1231 = unuse_way == 3'h4 ? ram_0_7 : _GEN_959; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1232 = unuse_way == 3'h4 ? ram_0_8 : _GEN_960; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1233 = unuse_way == 3'h4 ? ram_0_9 : _GEN_961; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1234 = unuse_way == 3'h4 ? ram_0_10 : _GEN_962; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1235 = unuse_way == 3'h4 ? ram_0_11 : _GEN_963; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1236 = unuse_way == 3'h4 ? ram_0_12 : _GEN_964; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1237 = unuse_way == 3'h4 ? ram_0_13 : _GEN_965; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1238 = unuse_way == 3'h4 ? ram_0_14 : _GEN_966; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1239 = unuse_way == 3'h4 ? ram_0_15 : _GEN_967; // @[i_cache.scala 100:40 19:24]
  wire [31:0] _GEN_1240 = unuse_way == 3'h4 ? tag_0_0 : _GEN_968; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1241 = unuse_way == 3'h4 ? tag_0_1 : _GEN_969; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1242 = unuse_way == 3'h4 ? tag_0_2 : _GEN_970; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1243 = unuse_way == 3'h4 ? tag_0_3 : _GEN_971; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1244 = unuse_way == 3'h4 ? tag_0_4 : _GEN_972; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1245 = unuse_way == 3'h4 ? tag_0_5 : _GEN_973; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1246 = unuse_way == 3'h4 ? tag_0_6 : _GEN_974; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1247 = unuse_way == 3'h4 ? tag_0_7 : _GEN_975; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1248 = unuse_way == 3'h4 ? tag_0_8 : _GEN_976; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1249 = unuse_way == 3'h4 ? tag_0_9 : _GEN_977; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1250 = unuse_way == 3'h4 ? tag_0_10 : _GEN_978; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1251 = unuse_way == 3'h4 ? tag_0_11 : _GEN_979; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1252 = unuse_way == 3'h4 ? tag_0_12 : _GEN_980; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1253 = unuse_way == 3'h4 ? tag_0_13 : _GEN_981; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1254 = unuse_way == 3'h4 ? tag_0_14 : _GEN_982; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1255 = unuse_way == 3'h4 ? tag_0_15 : _GEN_983; // @[i_cache.scala 100:40 23:24]
  wire  _GEN_1256 = unuse_way == 3'h4 ? valid_0_0 : _GEN_984; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1257 = unuse_way == 3'h4 ? valid_0_1 : _GEN_985; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1258 = unuse_way == 3'h4 ? valid_0_2 : _GEN_986; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1259 = unuse_way == 3'h4 ? valid_0_3 : _GEN_987; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1260 = unuse_way == 3'h4 ? valid_0_4 : _GEN_988; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1261 = unuse_way == 3'h4 ? valid_0_5 : _GEN_989; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1262 = unuse_way == 3'h4 ? valid_0_6 : _GEN_990; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1263 = unuse_way == 3'h4 ? valid_0_7 : _GEN_991; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1264 = unuse_way == 3'h4 ? valid_0_8 : _GEN_992; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1265 = unuse_way == 3'h4 ? valid_0_9 : _GEN_993; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1266 = unuse_way == 3'h4 ? valid_0_10 : _GEN_994; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1267 = unuse_way == 3'h4 ? valid_0_11 : _GEN_995; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1268 = unuse_way == 3'h4 ? valid_0_12 : _GEN_996; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1269 = unuse_way == 3'h4 ? valid_0_13 : _GEN_997; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1270 = unuse_way == 3'h4 ? valid_0_14 : _GEN_998; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1271 = unuse_way == 3'h4 ? valid_0_15 : _GEN_999; // @[i_cache.scala 100:40 27:26]
  wire [511:0] _GEN_1272 = unuse_way == 3'h4 ? ram_1_0 : _GEN_1016; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1273 = unuse_way == 3'h4 ? ram_1_1 : _GEN_1017; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1274 = unuse_way == 3'h4 ? ram_1_2 : _GEN_1018; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1275 = unuse_way == 3'h4 ? ram_1_3 : _GEN_1019; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1276 = unuse_way == 3'h4 ? ram_1_4 : _GEN_1020; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1277 = unuse_way == 3'h4 ? ram_1_5 : _GEN_1021; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1278 = unuse_way == 3'h4 ? ram_1_6 : _GEN_1022; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1279 = unuse_way == 3'h4 ? ram_1_7 : _GEN_1023; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1280 = unuse_way == 3'h4 ? ram_1_8 : _GEN_1024; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1281 = unuse_way == 3'h4 ? ram_1_9 : _GEN_1025; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1282 = unuse_way == 3'h4 ? ram_1_10 : _GEN_1026; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1283 = unuse_way == 3'h4 ? ram_1_11 : _GEN_1027; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1284 = unuse_way == 3'h4 ? ram_1_12 : _GEN_1028; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1285 = unuse_way == 3'h4 ? ram_1_13 : _GEN_1029; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1286 = unuse_way == 3'h4 ? ram_1_14 : _GEN_1030; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1287 = unuse_way == 3'h4 ? ram_1_15 : _GEN_1031; // @[i_cache.scala 100:40 20:24]
  wire [31:0] _GEN_1288 = unuse_way == 3'h4 ? tag_1_0 : _GEN_1032; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1289 = unuse_way == 3'h4 ? tag_1_1 : _GEN_1033; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1290 = unuse_way == 3'h4 ? tag_1_2 : _GEN_1034; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1291 = unuse_way == 3'h4 ? tag_1_3 : _GEN_1035; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1292 = unuse_way == 3'h4 ? tag_1_4 : _GEN_1036; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1293 = unuse_way == 3'h4 ? tag_1_5 : _GEN_1037; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1294 = unuse_way == 3'h4 ? tag_1_6 : _GEN_1038; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1295 = unuse_way == 3'h4 ? tag_1_7 : _GEN_1039; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1296 = unuse_way == 3'h4 ? tag_1_8 : _GEN_1040; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1297 = unuse_way == 3'h4 ? tag_1_9 : _GEN_1041; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1298 = unuse_way == 3'h4 ? tag_1_10 : _GEN_1042; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1299 = unuse_way == 3'h4 ? tag_1_11 : _GEN_1043; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1300 = unuse_way == 3'h4 ? tag_1_12 : _GEN_1044; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1301 = unuse_way == 3'h4 ? tag_1_13 : _GEN_1045; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1302 = unuse_way == 3'h4 ? tag_1_14 : _GEN_1046; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1303 = unuse_way == 3'h4 ? tag_1_15 : _GEN_1047; // @[i_cache.scala 100:40 24:24]
  wire  _GEN_1304 = unuse_way == 3'h4 ? valid_1_0 : _GEN_1048; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1305 = unuse_way == 3'h4 ? valid_1_1 : _GEN_1049; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1306 = unuse_way == 3'h4 ? valid_1_2 : _GEN_1050; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1307 = unuse_way == 3'h4 ? valid_1_3 : _GEN_1051; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1308 = unuse_way == 3'h4 ? valid_1_4 : _GEN_1052; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1309 = unuse_way == 3'h4 ? valid_1_5 : _GEN_1053; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1310 = unuse_way == 3'h4 ? valid_1_6 : _GEN_1054; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1311 = unuse_way == 3'h4 ? valid_1_7 : _GEN_1055; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1312 = unuse_way == 3'h4 ? valid_1_8 : _GEN_1056; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1313 = unuse_way == 3'h4 ? valid_1_9 : _GEN_1057; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1314 = unuse_way == 3'h4 ? valid_1_10 : _GEN_1058; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1315 = unuse_way == 3'h4 ? valid_1_11 : _GEN_1059; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1316 = unuse_way == 3'h4 ? valid_1_12 : _GEN_1060; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1317 = unuse_way == 3'h4 ? valid_1_13 : _GEN_1061; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1318 = unuse_way == 3'h4 ? valid_1_14 : _GEN_1062; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1319 = unuse_way == 3'h4 ? valid_1_15 : _GEN_1063; // @[i_cache.scala 100:40 28:26]
  wire [511:0] _GEN_1320 = unuse_way == 3'h4 ? ram_2_0 : _GEN_1064; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1321 = unuse_way == 3'h4 ? ram_2_1 : _GEN_1065; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1322 = unuse_way == 3'h4 ? ram_2_2 : _GEN_1066; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1323 = unuse_way == 3'h4 ? ram_2_3 : _GEN_1067; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1324 = unuse_way == 3'h4 ? ram_2_4 : _GEN_1068; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1325 = unuse_way == 3'h4 ? ram_2_5 : _GEN_1069; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1326 = unuse_way == 3'h4 ? ram_2_6 : _GEN_1070; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1327 = unuse_way == 3'h4 ? ram_2_7 : _GEN_1071; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1328 = unuse_way == 3'h4 ? ram_2_8 : _GEN_1072; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1329 = unuse_way == 3'h4 ? ram_2_9 : _GEN_1073; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1330 = unuse_way == 3'h4 ? ram_2_10 : _GEN_1074; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1331 = unuse_way == 3'h4 ? ram_2_11 : _GEN_1075; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1332 = unuse_way == 3'h4 ? ram_2_12 : _GEN_1076; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1333 = unuse_way == 3'h4 ? ram_2_13 : _GEN_1077; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1334 = unuse_way == 3'h4 ? ram_2_14 : _GEN_1078; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1335 = unuse_way == 3'h4 ? ram_2_15 : _GEN_1079; // @[i_cache.scala 100:40 21:24]
  wire [31:0] _GEN_1336 = unuse_way == 3'h4 ? tag_2_0 : _GEN_1080; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1337 = unuse_way == 3'h4 ? tag_2_1 : _GEN_1081; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1338 = unuse_way == 3'h4 ? tag_2_2 : _GEN_1082; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1339 = unuse_way == 3'h4 ? tag_2_3 : _GEN_1083; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1340 = unuse_way == 3'h4 ? tag_2_4 : _GEN_1084; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1341 = unuse_way == 3'h4 ? tag_2_5 : _GEN_1085; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1342 = unuse_way == 3'h4 ? tag_2_6 : _GEN_1086; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1343 = unuse_way == 3'h4 ? tag_2_7 : _GEN_1087; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1344 = unuse_way == 3'h4 ? tag_2_8 : _GEN_1088; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1345 = unuse_way == 3'h4 ? tag_2_9 : _GEN_1089; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1346 = unuse_way == 3'h4 ? tag_2_10 : _GEN_1090; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1347 = unuse_way == 3'h4 ? tag_2_11 : _GEN_1091; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1348 = unuse_way == 3'h4 ? tag_2_12 : _GEN_1092; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1349 = unuse_way == 3'h4 ? tag_2_13 : _GEN_1093; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1350 = unuse_way == 3'h4 ? tag_2_14 : _GEN_1094; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1351 = unuse_way == 3'h4 ? tag_2_15 : _GEN_1095; // @[i_cache.scala 100:40 25:24]
  wire  _GEN_1352 = unuse_way == 3'h4 ? valid_2_0 : _GEN_1096; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1353 = unuse_way == 3'h4 ? valid_2_1 : _GEN_1097; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1354 = unuse_way == 3'h4 ? valid_2_2 : _GEN_1098; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1355 = unuse_way == 3'h4 ? valid_2_3 : _GEN_1099; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1356 = unuse_way == 3'h4 ? valid_2_4 : _GEN_1100; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1357 = unuse_way == 3'h4 ? valid_2_5 : _GEN_1101; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1358 = unuse_way == 3'h4 ? valid_2_6 : _GEN_1102; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1359 = unuse_way == 3'h4 ? valid_2_7 : _GEN_1103; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1360 = unuse_way == 3'h4 ? valid_2_8 : _GEN_1104; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1361 = unuse_way == 3'h4 ? valid_2_9 : _GEN_1105; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1362 = unuse_way == 3'h4 ? valid_2_10 : _GEN_1106; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1363 = unuse_way == 3'h4 ? valid_2_11 : _GEN_1107; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1364 = unuse_way == 3'h4 ? valid_2_12 : _GEN_1108; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1365 = unuse_way == 3'h4 ? valid_2_13 : _GEN_1109; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1366 = unuse_way == 3'h4 ? valid_2_14 : _GEN_1110; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1367 = unuse_way == 3'h4 ? valid_2_15 : _GEN_1111; // @[i_cache.scala 100:40 29:26]
  wire [511:0] _GEN_1368 = unuse_way == 3'h3 ? _GEN_296 : _GEN_1320; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1369 = unuse_way == 3'h3 ? _GEN_297 : _GEN_1321; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1370 = unuse_way == 3'h3 ? _GEN_298 : _GEN_1322; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1371 = unuse_way == 3'h3 ? _GEN_299 : _GEN_1323; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1372 = unuse_way == 3'h3 ? _GEN_300 : _GEN_1324; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1373 = unuse_way == 3'h3 ? _GEN_301 : _GEN_1325; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1374 = unuse_way == 3'h3 ? _GEN_302 : _GEN_1326; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1375 = unuse_way == 3'h3 ? _GEN_303 : _GEN_1327; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1376 = unuse_way == 3'h3 ? _GEN_304 : _GEN_1328; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1377 = unuse_way == 3'h3 ? _GEN_305 : _GEN_1329; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1378 = unuse_way == 3'h3 ? _GEN_306 : _GEN_1330; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1379 = unuse_way == 3'h3 ? _GEN_307 : _GEN_1331; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1380 = unuse_way == 3'h3 ? _GEN_308 : _GEN_1332; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1381 = unuse_way == 3'h3 ? _GEN_309 : _GEN_1333; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1382 = unuse_way == 3'h3 ? _GEN_310 : _GEN_1334; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1383 = unuse_way == 3'h3 ? _GEN_311 : _GEN_1335; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1384 = unuse_way == 3'h3 ? _GEN_312 : _GEN_1336; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1385 = unuse_way == 3'h3 ? _GEN_313 : _GEN_1337; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1386 = unuse_way == 3'h3 ? _GEN_314 : _GEN_1338; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1387 = unuse_way == 3'h3 ? _GEN_315 : _GEN_1339; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1388 = unuse_way == 3'h3 ? _GEN_316 : _GEN_1340; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1389 = unuse_way == 3'h3 ? _GEN_317 : _GEN_1341; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1390 = unuse_way == 3'h3 ? _GEN_318 : _GEN_1342; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1391 = unuse_way == 3'h3 ? _GEN_319 : _GEN_1343; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1392 = unuse_way == 3'h3 ? _GEN_320 : _GEN_1344; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1393 = unuse_way == 3'h3 ? _GEN_321 : _GEN_1345; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1394 = unuse_way == 3'h3 ? _GEN_322 : _GEN_1346; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1395 = unuse_way == 3'h3 ? _GEN_323 : _GEN_1347; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1396 = unuse_way == 3'h3 ? _GEN_324 : _GEN_1348; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1397 = unuse_way == 3'h3 ? _GEN_325 : _GEN_1349; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1398 = unuse_way == 3'h3 ? _GEN_326 : _GEN_1350; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1399 = unuse_way == 3'h3 ? _GEN_327 : _GEN_1351; // @[i_cache.scala 95:40]
  wire  _GEN_1400 = unuse_way == 3'h3 ? _GEN_328 : _GEN_1352; // @[i_cache.scala 95:40]
  wire  _GEN_1401 = unuse_way == 3'h3 ? _GEN_329 : _GEN_1353; // @[i_cache.scala 95:40]
  wire  _GEN_1402 = unuse_way == 3'h3 ? _GEN_330 : _GEN_1354; // @[i_cache.scala 95:40]
  wire  _GEN_1403 = unuse_way == 3'h3 ? _GEN_331 : _GEN_1355; // @[i_cache.scala 95:40]
  wire  _GEN_1404 = unuse_way == 3'h3 ? _GEN_332 : _GEN_1356; // @[i_cache.scala 95:40]
  wire  _GEN_1405 = unuse_way == 3'h3 ? _GEN_333 : _GEN_1357; // @[i_cache.scala 95:40]
  wire  _GEN_1406 = unuse_way == 3'h3 ? _GEN_334 : _GEN_1358; // @[i_cache.scala 95:40]
  wire  _GEN_1407 = unuse_way == 3'h3 ? _GEN_335 : _GEN_1359; // @[i_cache.scala 95:40]
  wire  _GEN_1408 = unuse_way == 3'h3 ? _GEN_336 : _GEN_1360; // @[i_cache.scala 95:40]
  wire  _GEN_1409 = unuse_way == 3'h3 ? _GEN_337 : _GEN_1361; // @[i_cache.scala 95:40]
  wire  _GEN_1410 = unuse_way == 3'h3 ? _GEN_338 : _GEN_1362; // @[i_cache.scala 95:40]
  wire  _GEN_1411 = unuse_way == 3'h3 ? _GEN_339 : _GEN_1363; // @[i_cache.scala 95:40]
  wire  _GEN_1412 = unuse_way == 3'h3 ? _GEN_340 : _GEN_1364; // @[i_cache.scala 95:40]
  wire  _GEN_1413 = unuse_way == 3'h3 ? _GEN_341 : _GEN_1365; // @[i_cache.scala 95:40]
  wire  _GEN_1414 = unuse_way == 3'h3 ? _GEN_342 : _GEN_1366; // @[i_cache.scala 95:40]
  wire  _GEN_1415 = unuse_way == 3'h3 ? _GEN_343 : _GEN_1367; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1416 = unuse_way == 3'h3 ? _GEN_344 : _GEN_1208; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1417 = unuse_way == 3'h3 ? _GEN_345 : _GEN_1209; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1418 = unuse_way == 3'h3 ? _GEN_346 : _GEN_1210; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1419 = unuse_way == 3'h3 ? _GEN_347 : _GEN_1211; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1420 = unuse_way == 3'h3 ? _GEN_348 : _GEN_1212; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1421 = unuse_way == 3'h3 ? _GEN_349 : _GEN_1213; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1422 = unuse_way == 3'h3 ? _GEN_350 : _GEN_1214; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1423 = unuse_way == 3'h3 ? _GEN_351 : _GEN_1215; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1424 = unuse_way == 3'h3 ? _GEN_352 : _GEN_1216; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1425 = unuse_way == 3'h3 ? _GEN_353 : _GEN_1217; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1426 = unuse_way == 3'h3 ? _GEN_354 : _GEN_1218; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1427 = unuse_way == 3'h3 ? _GEN_355 : _GEN_1219; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1428 = unuse_way == 3'h3 ? _GEN_356 : _GEN_1220; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1429 = unuse_way == 3'h3 ? _GEN_357 : _GEN_1221; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1430 = unuse_way == 3'h3 ? _GEN_358 : _GEN_1222; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1431 = unuse_way == 3'h3 ? _GEN_359 : _GEN_1223; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1432 = unuse_way == 3'h3 ? ram_3_0 : _GEN_1160; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1433 = unuse_way == 3'h3 ? ram_3_1 : _GEN_1161; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1434 = unuse_way == 3'h3 ? ram_3_2 : _GEN_1162; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1435 = unuse_way == 3'h3 ? ram_3_3 : _GEN_1163; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1436 = unuse_way == 3'h3 ? ram_3_4 : _GEN_1164; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1437 = unuse_way == 3'h3 ? ram_3_5 : _GEN_1165; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1438 = unuse_way == 3'h3 ? ram_3_6 : _GEN_1166; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1439 = unuse_way == 3'h3 ? ram_3_7 : _GEN_1167; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1440 = unuse_way == 3'h3 ? ram_3_8 : _GEN_1168; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1441 = unuse_way == 3'h3 ? ram_3_9 : _GEN_1169; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1442 = unuse_way == 3'h3 ? ram_3_10 : _GEN_1170; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1443 = unuse_way == 3'h3 ? ram_3_11 : _GEN_1171; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1444 = unuse_way == 3'h3 ? ram_3_12 : _GEN_1172; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1445 = unuse_way == 3'h3 ? ram_3_13 : _GEN_1173; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1446 = unuse_way == 3'h3 ? ram_3_14 : _GEN_1174; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1447 = unuse_way == 3'h3 ? ram_3_15 : _GEN_1175; // @[i_cache.scala 22:24 95:40]
  wire [31:0] _GEN_1448 = unuse_way == 3'h3 ? tag_3_0 : _GEN_1176; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1449 = unuse_way == 3'h3 ? tag_3_1 : _GEN_1177; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1450 = unuse_way == 3'h3 ? tag_3_2 : _GEN_1178; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1451 = unuse_way == 3'h3 ? tag_3_3 : _GEN_1179; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1452 = unuse_way == 3'h3 ? tag_3_4 : _GEN_1180; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1453 = unuse_way == 3'h3 ? tag_3_5 : _GEN_1181; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1454 = unuse_way == 3'h3 ? tag_3_6 : _GEN_1182; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1455 = unuse_way == 3'h3 ? tag_3_7 : _GEN_1183; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1456 = unuse_way == 3'h3 ? tag_3_8 : _GEN_1184; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1457 = unuse_way == 3'h3 ? tag_3_9 : _GEN_1185; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1458 = unuse_way == 3'h3 ? tag_3_10 : _GEN_1186; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1459 = unuse_way == 3'h3 ? tag_3_11 : _GEN_1187; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1460 = unuse_way == 3'h3 ? tag_3_12 : _GEN_1188; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1461 = unuse_way == 3'h3 ? tag_3_13 : _GEN_1189; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1462 = unuse_way == 3'h3 ? tag_3_14 : _GEN_1190; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1463 = unuse_way == 3'h3 ? tag_3_15 : _GEN_1191; // @[i_cache.scala 26:24 95:40]
  wire  _GEN_1464 = unuse_way == 3'h3 ? valid_3_0 : _GEN_1192; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1465 = unuse_way == 3'h3 ? valid_3_1 : _GEN_1193; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1466 = unuse_way == 3'h3 ? valid_3_2 : _GEN_1194; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1467 = unuse_way == 3'h3 ? valid_3_3 : _GEN_1195; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1468 = unuse_way == 3'h3 ? valid_3_4 : _GEN_1196; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1469 = unuse_way == 3'h3 ? valid_3_5 : _GEN_1197; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1470 = unuse_way == 3'h3 ? valid_3_6 : _GEN_1198; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1471 = unuse_way == 3'h3 ? valid_3_7 : _GEN_1199; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1472 = unuse_way == 3'h3 ? valid_3_8 : _GEN_1200; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1473 = unuse_way == 3'h3 ? valid_3_9 : _GEN_1201; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1474 = unuse_way == 3'h3 ? valid_3_10 : _GEN_1202; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1475 = unuse_way == 3'h3 ? valid_3_11 : _GEN_1203; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1476 = unuse_way == 3'h3 ? valid_3_12 : _GEN_1204; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1477 = unuse_way == 3'h3 ? valid_3_13 : _GEN_1205; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1478 = unuse_way == 3'h3 ? valid_3_14 : _GEN_1206; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1479 = unuse_way == 3'h3 ? valid_3_15 : _GEN_1207; // @[i_cache.scala 30:26 95:40]
  wire [511:0] _GEN_1480 = unuse_way == 3'h3 ? ram_0_0 : _GEN_1224; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1481 = unuse_way == 3'h3 ? ram_0_1 : _GEN_1225; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1482 = unuse_way == 3'h3 ? ram_0_2 : _GEN_1226; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1483 = unuse_way == 3'h3 ? ram_0_3 : _GEN_1227; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1484 = unuse_way == 3'h3 ? ram_0_4 : _GEN_1228; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1485 = unuse_way == 3'h3 ? ram_0_5 : _GEN_1229; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1486 = unuse_way == 3'h3 ? ram_0_6 : _GEN_1230; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1487 = unuse_way == 3'h3 ? ram_0_7 : _GEN_1231; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1488 = unuse_way == 3'h3 ? ram_0_8 : _GEN_1232; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1489 = unuse_way == 3'h3 ? ram_0_9 : _GEN_1233; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1490 = unuse_way == 3'h3 ? ram_0_10 : _GEN_1234; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1491 = unuse_way == 3'h3 ? ram_0_11 : _GEN_1235; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1492 = unuse_way == 3'h3 ? ram_0_12 : _GEN_1236; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1493 = unuse_way == 3'h3 ? ram_0_13 : _GEN_1237; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1494 = unuse_way == 3'h3 ? ram_0_14 : _GEN_1238; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1495 = unuse_way == 3'h3 ? ram_0_15 : _GEN_1239; // @[i_cache.scala 19:24 95:40]
  wire [31:0] _GEN_1496 = unuse_way == 3'h3 ? tag_0_0 : _GEN_1240; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1497 = unuse_way == 3'h3 ? tag_0_1 : _GEN_1241; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1498 = unuse_way == 3'h3 ? tag_0_2 : _GEN_1242; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1499 = unuse_way == 3'h3 ? tag_0_3 : _GEN_1243; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1500 = unuse_way == 3'h3 ? tag_0_4 : _GEN_1244; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1501 = unuse_way == 3'h3 ? tag_0_5 : _GEN_1245; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1502 = unuse_way == 3'h3 ? tag_0_6 : _GEN_1246; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1503 = unuse_way == 3'h3 ? tag_0_7 : _GEN_1247; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1504 = unuse_way == 3'h3 ? tag_0_8 : _GEN_1248; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1505 = unuse_way == 3'h3 ? tag_0_9 : _GEN_1249; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1506 = unuse_way == 3'h3 ? tag_0_10 : _GEN_1250; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1507 = unuse_way == 3'h3 ? tag_0_11 : _GEN_1251; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1508 = unuse_way == 3'h3 ? tag_0_12 : _GEN_1252; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1509 = unuse_way == 3'h3 ? tag_0_13 : _GEN_1253; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1510 = unuse_way == 3'h3 ? tag_0_14 : _GEN_1254; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1511 = unuse_way == 3'h3 ? tag_0_15 : _GEN_1255; // @[i_cache.scala 23:24 95:40]
  wire  _GEN_1512 = unuse_way == 3'h3 ? valid_0_0 : _GEN_1256; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1513 = unuse_way == 3'h3 ? valid_0_1 : _GEN_1257; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1514 = unuse_way == 3'h3 ? valid_0_2 : _GEN_1258; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1515 = unuse_way == 3'h3 ? valid_0_3 : _GEN_1259; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1516 = unuse_way == 3'h3 ? valid_0_4 : _GEN_1260; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1517 = unuse_way == 3'h3 ? valid_0_5 : _GEN_1261; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1518 = unuse_way == 3'h3 ? valid_0_6 : _GEN_1262; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1519 = unuse_way == 3'h3 ? valid_0_7 : _GEN_1263; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1520 = unuse_way == 3'h3 ? valid_0_8 : _GEN_1264; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1521 = unuse_way == 3'h3 ? valid_0_9 : _GEN_1265; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1522 = unuse_way == 3'h3 ? valid_0_10 : _GEN_1266; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1523 = unuse_way == 3'h3 ? valid_0_11 : _GEN_1267; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1524 = unuse_way == 3'h3 ? valid_0_12 : _GEN_1268; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1525 = unuse_way == 3'h3 ? valid_0_13 : _GEN_1269; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1526 = unuse_way == 3'h3 ? valid_0_14 : _GEN_1270; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1527 = unuse_way == 3'h3 ? valid_0_15 : _GEN_1271; // @[i_cache.scala 27:26 95:40]
  wire [511:0] _GEN_1528 = unuse_way == 3'h3 ? ram_1_0 : _GEN_1272; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1529 = unuse_way == 3'h3 ? ram_1_1 : _GEN_1273; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1530 = unuse_way == 3'h3 ? ram_1_2 : _GEN_1274; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1531 = unuse_way == 3'h3 ? ram_1_3 : _GEN_1275; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1532 = unuse_way == 3'h3 ? ram_1_4 : _GEN_1276; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1533 = unuse_way == 3'h3 ? ram_1_5 : _GEN_1277; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1534 = unuse_way == 3'h3 ? ram_1_6 : _GEN_1278; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1535 = unuse_way == 3'h3 ? ram_1_7 : _GEN_1279; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1536 = unuse_way == 3'h3 ? ram_1_8 : _GEN_1280; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1537 = unuse_way == 3'h3 ? ram_1_9 : _GEN_1281; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1538 = unuse_way == 3'h3 ? ram_1_10 : _GEN_1282; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1539 = unuse_way == 3'h3 ? ram_1_11 : _GEN_1283; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1540 = unuse_way == 3'h3 ? ram_1_12 : _GEN_1284; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1541 = unuse_way == 3'h3 ? ram_1_13 : _GEN_1285; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1542 = unuse_way == 3'h3 ? ram_1_14 : _GEN_1286; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1543 = unuse_way == 3'h3 ? ram_1_15 : _GEN_1287; // @[i_cache.scala 20:24 95:40]
  wire [31:0] _GEN_1544 = unuse_way == 3'h3 ? tag_1_0 : _GEN_1288; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1545 = unuse_way == 3'h3 ? tag_1_1 : _GEN_1289; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1546 = unuse_way == 3'h3 ? tag_1_2 : _GEN_1290; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1547 = unuse_way == 3'h3 ? tag_1_3 : _GEN_1291; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1548 = unuse_way == 3'h3 ? tag_1_4 : _GEN_1292; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1549 = unuse_way == 3'h3 ? tag_1_5 : _GEN_1293; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1550 = unuse_way == 3'h3 ? tag_1_6 : _GEN_1294; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1551 = unuse_way == 3'h3 ? tag_1_7 : _GEN_1295; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1552 = unuse_way == 3'h3 ? tag_1_8 : _GEN_1296; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1553 = unuse_way == 3'h3 ? tag_1_9 : _GEN_1297; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1554 = unuse_way == 3'h3 ? tag_1_10 : _GEN_1298; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1555 = unuse_way == 3'h3 ? tag_1_11 : _GEN_1299; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1556 = unuse_way == 3'h3 ? tag_1_12 : _GEN_1300; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1557 = unuse_way == 3'h3 ? tag_1_13 : _GEN_1301; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1558 = unuse_way == 3'h3 ? tag_1_14 : _GEN_1302; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1559 = unuse_way == 3'h3 ? tag_1_15 : _GEN_1303; // @[i_cache.scala 24:24 95:40]
  wire  _GEN_1560 = unuse_way == 3'h3 ? valid_1_0 : _GEN_1304; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1561 = unuse_way == 3'h3 ? valid_1_1 : _GEN_1305; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1562 = unuse_way == 3'h3 ? valid_1_2 : _GEN_1306; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1563 = unuse_way == 3'h3 ? valid_1_3 : _GEN_1307; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1564 = unuse_way == 3'h3 ? valid_1_4 : _GEN_1308; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1565 = unuse_way == 3'h3 ? valid_1_5 : _GEN_1309; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1566 = unuse_way == 3'h3 ? valid_1_6 : _GEN_1310; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1567 = unuse_way == 3'h3 ? valid_1_7 : _GEN_1311; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1568 = unuse_way == 3'h3 ? valid_1_8 : _GEN_1312; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1569 = unuse_way == 3'h3 ? valid_1_9 : _GEN_1313; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1570 = unuse_way == 3'h3 ? valid_1_10 : _GEN_1314; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1571 = unuse_way == 3'h3 ? valid_1_11 : _GEN_1315; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1572 = unuse_way == 3'h3 ? valid_1_12 : _GEN_1316; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1573 = unuse_way == 3'h3 ? valid_1_13 : _GEN_1317; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1574 = unuse_way == 3'h3 ? valid_1_14 : _GEN_1318; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1575 = unuse_way == 3'h3 ? valid_1_15 : _GEN_1319; // @[i_cache.scala 28:26 95:40]
  wire [511:0] _GEN_1576 = unuse_way == 3'h2 ? _GEN_232 : _GEN_1528; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1577 = unuse_way == 3'h2 ? _GEN_233 : _GEN_1529; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1578 = unuse_way == 3'h2 ? _GEN_234 : _GEN_1530; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1579 = unuse_way == 3'h2 ? _GEN_235 : _GEN_1531; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1580 = unuse_way == 3'h2 ? _GEN_236 : _GEN_1532; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1581 = unuse_way == 3'h2 ? _GEN_237 : _GEN_1533; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1582 = unuse_way == 3'h2 ? _GEN_238 : _GEN_1534; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1583 = unuse_way == 3'h2 ? _GEN_239 : _GEN_1535; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1584 = unuse_way == 3'h2 ? _GEN_240 : _GEN_1536; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1585 = unuse_way == 3'h2 ? _GEN_241 : _GEN_1537; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1586 = unuse_way == 3'h2 ? _GEN_242 : _GEN_1538; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1587 = unuse_way == 3'h2 ? _GEN_243 : _GEN_1539; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1588 = unuse_way == 3'h2 ? _GEN_244 : _GEN_1540; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1589 = unuse_way == 3'h2 ? _GEN_245 : _GEN_1541; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1590 = unuse_way == 3'h2 ? _GEN_246 : _GEN_1542; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1591 = unuse_way == 3'h2 ? _GEN_247 : _GEN_1543; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1592 = unuse_way == 3'h2 ? _GEN_248 : _GEN_1544; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1593 = unuse_way == 3'h2 ? _GEN_249 : _GEN_1545; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1594 = unuse_way == 3'h2 ? _GEN_250 : _GEN_1546; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1595 = unuse_way == 3'h2 ? _GEN_251 : _GEN_1547; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1596 = unuse_way == 3'h2 ? _GEN_252 : _GEN_1548; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1597 = unuse_way == 3'h2 ? _GEN_253 : _GEN_1549; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1598 = unuse_way == 3'h2 ? _GEN_254 : _GEN_1550; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1599 = unuse_way == 3'h2 ? _GEN_255 : _GEN_1551; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1600 = unuse_way == 3'h2 ? _GEN_256 : _GEN_1552; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1601 = unuse_way == 3'h2 ? _GEN_257 : _GEN_1553; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1602 = unuse_way == 3'h2 ? _GEN_258 : _GEN_1554; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1603 = unuse_way == 3'h2 ? _GEN_259 : _GEN_1555; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1604 = unuse_way == 3'h2 ? _GEN_260 : _GEN_1556; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1605 = unuse_way == 3'h2 ? _GEN_261 : _GEN_1557; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1606 = unuse_way == 3'h2 ? _GEN_262 : _GEN_1558; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1607 = unuse_way == 3'h2 ? _GEN_263 : _GEN_1559; // @[i_cache.scala 90:40]
  wire  _GEN_1608 = unuse_way == 3'h2 ? _GEN_264 : _GEN_1560; // @[i_cache.scala 90:40]
  wire  _GEN_1609 = unuse_way == 3'h2 ? _GEN_265 : _GEN_1561; // @[i_cache.scala 90:40]
  wire  _GEN_1610 = unuse_way == 3'h2 ? _GEN_266 : _GEN_1562; // @[i_cache.scala 90:40]
  wire  _GEN_1611 = unuse_way == 3'h2 ? _GEN_267 : _GEN_1563; // @[i_cache.scala 90:40]
  wire  _GEN_1612 = unuse_way == 3'h2 ? _GEN_268 : _GEN_1564; // @[i_cache.scala 90:40]
  wire  _GEN_1613 = unuse_way == 3'h2 ? _GEN_269 : _GEN_1565; // @[i_cache.scala 90:40]
  wire  _GEN_1614 = unuse_way == 3'h2 ? _GEN_270 : _GEN_1566; // @[i_cache.scala 90:40]
  wire  _GEN_1615 = unuse_way == 3'h2 ? _GEN_271 : _GEN_1567; // @[i_cache.scala 90:40]
  wire  _GEN_1616 = unuse_way == 3'h2 ? _GEN_272 : _GEN_1568; // @[i_cache.scala 90:40]
  wire  _GEN_1617 = unuse_way == 3'h2 ? _GEN_273 : _GEN_1569; // @[i_cache.scala 90:40]
  wire  _GEN_1618 = unuse_way == 3'h2 ? _GEN_274 : _GEN_1570; // @[i_cache.scala 90:40]
  wire  _GEN_1619 = unuse_way == 3'h2 ? _GEN_275 : _GEN_1571; // @[i_cache.scala 90:40]
  wire  _GEN_1620 = unuse_way == 3'h2 ? _GEN_276 : _GEN_1572; // @[i_cache.scala 90:40]
  wire  _GEN_1621 = unuse_way == 3'h2 ? _GEN_277 : _GEN_1573; // @[i_cache.scala 90:40]
  wire  _GEN_1622 = unuse_way == 3'h2 ? _GEN_278 : _GEN_1574; // @[i_cache.scala 90:40]
  wire  _GEN_1623 = unuse_way == 3'h2 ? _GEN_279 : _GEN_1575; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1624 = unuse_way == 3'h2 ? _GEN_280 : _GEN_1416; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1625 = unuse_way == 3'h2 ? _GEN_281 : _GEN_1417; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1626 = unuse_way == 3'h2 ? _GEN_282 : _GEN_1418; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1627 = unuse_way == 3'h2 ? _GEN_283 : _GEN_1419; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1628 = unuse_way == 3'h2 ? _GEN_284 : _GEN_1420; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1629 = unuse_way == 3'h2 ? _GEN_285 : _GEN_1421; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1630 = unuse_way == 3'h2 ? _GEN_286 : _GEN_1422; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1631 = unuse_way == 3'h2 ? _GEN_287 : _GEN_1423; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1632 = unuse_way == 3'h2 ? _GEN_288 : _GEN_1424; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1633 = unuse_way == 3'h2 ? _GEN_289 : _GEN_1425; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1634 = unuse_way == 3'h2 ? _GEN_290 : _GEN_1426; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1635 = unuse_way == 3'h2 ? _GEN_291 : _GEN_1427; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1636 = unuse_way == 3'h2 ? _GEN_292 : _GEN_1428; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1637 = unuse_way == 3'h2 ? _GEN_293 : _GEN_1429; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1638 = unuse_way == 3'h2 ? _GEN_294 : _GEN_1430; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1639 = unuse_way == 3'h2 ? _GEN_295 : _GEN_1431; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1640 = unuse_way == 3'h2 ? ram_2_0 : _GEN_1368; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1641 = unuse_way == 3'h2 ? ram_2_1 : _GEN_1369; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1642 = unuse_way == 3'h2 ? ram_2_2 : _GEN_1370; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1643 = unuse_way == 3'h2 ? ram_2_3 : _GEN_1371; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1644 = unuse_way == 3'h2 ? ram_2_4 : _GEN_1372; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1645 = unuse_way == 3'h2 ? ram_2_5 : _GEN_1373; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1646 = unuse_way == 3'h2 ? ram_2_6 : _GEN_1374; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1647 = unuse_way == 3'h2 ? ram_2_7 : _GEN_1375; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1648 = unuse_way == 3'h2 ? ram_2_8 : _GEN_1376; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1649 = unuse_way == 3'h2 ? ram_2_9 : _GEN_1377; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1650 = unuse_way == 3'h2 ? ram_2_10 : _GEN_1378; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1651 = unuse_way == 3'h2 ? ram_2_11 : _GEN_1379; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1652 = unuse_way == 3'h2 ? ram_2_12 : _GEN_1380; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1653 = unuse_way == 3'h2 ? ram_2_13 : _GEN_1381; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1654 = unuse_way == 3'h2 ? ram_2_14 : _GEN_1382; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1655 = unuse_way == 3'h2 ? ram_2_15 : _GEN_1383; // @[i_cache.scala 21:24 90:40]
  wire [31:0] _GEN_1656 = unuse_way == 3'h2 ? tag_2_0 : _GEN_1384; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1657 = unuse_way == 3'h2 ? tag_2_1 : _GEN_1385; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1658 = unuse_way == 3'h2 ? tag_2_2 : _GEN_1386; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1659 = unuse_way == 3'h2 ? tag_2_3 : _GEN_1387; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1660 = unuse_way == 3'h2 ? tag_2_4 : _GEN_1388; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1661 = unuse_way == 3'h2 ? tag_2_5 : _GEN_1389; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1662 = unuse_way == 3'h2 ? tag_2_6 : _GEN_1390; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1663 = unuse_way == 3'h2 ? tag_2_7 : _GEN_1391; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1664 = unuse_way == 3'h2 ? tag_2_8 : _GEN_1392; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1665 = unuse_way == 3'h2 ? tag_2_9 : _GEN_1393; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1666 = unuse_way == 3'h2 ? tag_2_10 : _GEN_1394; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1667 = unuse_way == 3'h2 ? tag_2_11 : _GEN_1395; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1668 = unuse_way == 3'h2 ? tag_2_12 : _GEN_1396; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1669 = unuse_way == 3'h2 ? tag_2_13 : _GEN_1397; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1670 = unuse_way == 3'h2 ? tag_2_14 : _GEN_1398; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1671 = unuse_way == 3'h2 ? tag_2_15 : _GEN_1399; // @[i_cache.scala 25:24 90:40]
  wire  _GEN_1672 = unuse_way == 3'h2 ? valid_2_0 : _GEN_1400; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1673 = unuse_way == 3'h2 ? valid_2_1 : _GEN_1401; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1674 = unuse_way == 3'h2 ? valid_2_2 : _GEN_1402; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1675 = unuse_way == 3'h2 ? valid_2_3 : _GEN_1403; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1676 = unuse_way == 3'h2 ? valid_2_4 : _GEN_1404; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1677 = unuse_way == 3'h2 ? valid_2_5 : _GEN_1405; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1678 = unuse_way == 3'h2 ? valid_2_6 : _GEN_1406; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1679 = unuse_way == 3'h2 ? valid_2_7 : _GEN_1407; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1680 = unuse_way == 3'h2 ? valid_2_8 : _GEN_1408; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1681 = unuse_way == 3'h2 ? valid_2_9 : _GEN_1409; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1682 = unuse_way == 3'h2 ? valid_2_10 : _GEN_1410; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1683 = unuse_way == 3'h2 ? valid_2_11 : _GEN_1411; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1684 = unuse_way == 3'h2 ? valid_2_12 : _GEN_1412; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1685 = unuse_way == 3'h2 ? valid_2_13 : _GEN_1413; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1686 = unuse_way == 3'h2 ? valid_2_14 : _GEN_1414; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1687 = unuse_way == 3'h2 ? valid_2_15 : _GEN_1415; // @[i_cache.scala 29:26 90:40]
  wire [511:0] _GEN_1688 = unuse_way == 3'h2 ? ram_3_0 : _GEN_1432; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1689 = unuse_way == 3'h2 ? ram_3_1 : _GEN_1433; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1690 = unuse_way == 3'h2 ? ram_3_2 : _GEN_1434; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1691 = unuse_way == 3'h2 ? ram_3_3 : _GEN_1435; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1692 = unuse_way == 3'h2 ? ram_3_4 : _GEN_1436; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1693 = unuse_way == 3'h2 ? ram_3_5 : _GEN_1437; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1694 = unuse_way == 3'h2 ? ram_3_6 : _GEN_1438; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1695 = unuse_way == 3'h2 ? ram_3_7 : _GEN_1439; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1696 = unuse_way == 3'h2 ? ram_3_8 : _GEN_1440; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1697 = unuse_way == 3'h2 ? ram_3_9 : _GEN_1441; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1698 = unuse_way == 3'h2 ? ram_3_10 : _GEN_1442; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1699 = unuse_way == 3'h2 ? ram_3_11 : _GEN_1443; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1700 = unuse_way == 3'h2 ? ram_3_12 : _GEN_1444; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1701 = unuse_way == 3'h2 ? ram_3_13 : _GEN_1445; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1702 = unuse_way == 3'h2 ? ram_3_14 : _GEN_1446; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1703 = unuse_way == 3'h2 ? ram_3_15 : _GEN_1447; // @[i_cache.scala 22:24 90:40]
  wire [31:0] _GEN_1704 = unuse_way == 3'h2 ? tag_3_0 : _GEN_1448; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1705 = unuse_way == 3'h2 ? tag_3_1 : _GEN_1449; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1706 = unuse_way == 3'h2 ? tag_3_2 : _GEN_1450; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1707 = unuse_way == 3'h2 ? tag_3_3 : _GEN_1451; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1708 = unuse_way == 3'h2 ? tag_3_4 : _GEN_1452; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1709 = unuse_way == 3'h2 ? tag_3_5 : _GEN_1453; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1710 = unuse_way == 3'h2 ? tag_3_6 : _GEN_1454; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1711 = unuse_way == 3'h2 ? tag_3_7 : _GEN_1455; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1712 = unuse_way == 3'h2 ? tag_3_8 : _GEN_1456; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1713 = unuse_way == 3'h2 ? tag_3_9 : _GEN_1457; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1714 = unuse_way == 3'h2 ? tag_3_10 : _GEN_1458; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1715 = unuse_way == 3'h2 ? tag_3_11 : _GEN_1459; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1716 = unuse_way == 3'h2 ? tag_3_12 : _GEN_1460; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1717 = unuse_way == 3'h2 ? tag_3_13 : _GEN_1461; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1718 = unuse_way == 3'h2 ? tag_3_14 : _GEN_1462; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1719 = unuse_way == 3'h2 ? tag_3_15 : _GEN_1463; // @[i_cache.scala 26:24 90:40]
  wire  _GEN_1720 = unuse_way == 3'h2 ? valid_3_0 : _GEN_1464; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1721 = unuse_way == 3'h2 ? valid_3_1 : _GEN_1465; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1722 = unuse_way == 3'h2 ? valid_3_2 : _GEN_1466; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1723 = unuse_way == 3'h2 ? valid_3_3 : _GEN_1467; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1724 = unuse_way == 3'h2 ? valid_3_4 : _GEN_1468; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1725 = unuse_way == 3'h2 ? valid_3_5 : _GEN_1469; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1726 = unuse_way == 3'h2 ? valid_3_6 : _GEN_1470; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1727 = unuse_way == 3'h2 ? valid_3_7 : _GEN_1471; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1728 = unuse_way == 3'h2 ? valid_3_8 : _GEN_1472; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1729 = unuse_way == 3'h2 ? valid_3_9 : _GEN_1473; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1730 = unuse_way == 3'h2 ? valid_3_10 : _GEN_1474; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1731 = unuse_way == 3'h2 ? valid_3_11 : _GEN_1475; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1732 = unuse_way == 3'h2 ? valid_3_12 : _GEN_1476; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1733 = unuse_way == 3'h2 ? valid_3_13 : _GEN_1477; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1734 = unuse_way == 3'h2 ? valid_3_14 : _GEN_1478; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1735 = unuse_way == 3'h2 ? valid_3_15 : _GEN_1479; // @[i_cache.scala 30:26 90:40]
  wire [511:0] _GEN_1736 = unuse_way == 3'h2 ? ram_0_0 : _GEN_1480; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1737 = unuse_way == 3'h2 ? ram_0_1 : _GEN_1481; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1738 = unuse_way == 3'h2 ? ram_0_2 : _GEN_1482; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1739 = unuse_way == 3'h2 ? ram_0_3 : _GEN_1483; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1740 = unuse_way == 3'h2 ? ram_0_4 : _GEN_1484; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1741 = unuse_way == 3'h2 ? ram_0_5 : _GEN_1485; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1742 = unuse_way == 3'h2 ? ram_0_6 : _GEN_1486; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1743 = unuse_way == 3'h2 ? ram_0_7 : _GEN_1487; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1744 = unuse_way == 3'h2 ? ram_0_8 : _GEN_1488; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1745 = unuse_way == 3'h2 ? ram_0_9 : _GEN_1489; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1746 = unuse_way == 3'h2 ? ram_0_10 : _GEN_1490; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1747 = unuse_way == 3'h2 ? ram_0_11 : _GEN_1491; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1748 = unuse_way == 3'h2 ? ram_0_12 : _GEN_1492; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1749 = unuse_way == 3'h2 ? ram_0_13 : _GEN_1493; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1750 = unuse_way == 3'h2 ? ram_0_14 : _GEN_1494; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1751 = unuse_way == 3'h2 ? ram_0_15 : _GEN_1495; // @[i_cache.scala 19:24 90:40]
  wire [31:0] _GEN_1752 = unuse_way == 3'h2 ? tag_0_0 : _GEN_1496; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1753 = unuse_way == 3'h2 ? tag_0_1 : _GEN_1497; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1754 = unuse_way == 3'h2 ? tag_0_2 : _GEN_1498; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1755 = unuse_way == 3'h2 ? tag_0_3 : _GEN_1499; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1756 = unuse_way == 3'h2 ? tag_0_4 : _GEN_1500; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1757 = unuse_way == 3'h2 ? tag_0_5 : _GEN_1501; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1758 = unuse_way == 3'h2 ? tag_0_6 : _GEN_1502; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1759 = unuse_way == 3'h2 ? tag_0_7 : _GEN_1503; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1760 = unuse_way == 3'h2 ? tag_0_8 : _GEN_1504; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1761 = unuse_way == 3'h2 ? tag_0_9 : _GEN_1505; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1762 = unuse_way == 3'h2 ? tag_0_10 : _GEN_1506; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1763 = unuse_way == 3'h2 ? tag_0_11 : _GEN_1507; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1764 = unuse_way == 3'h2 ? tag_0_12 : _GEN_1508; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1765 = unuse_way == 3'h2 ? tag_0_13 : _GEN_1509; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1766 = unuse_way == 3'h2 ? tag_0_14 : _GEN_1510; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1767 = unuse_way == 3'h2 ? tag_0_15 : _GEN_1511; // @[i_cache.scala 23:24 90:40]
  wire  _GEN_1768 = unuse_way == 3'h2 ? valid_0_0 : _GEN_1512; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1769 = unuse_way == 3'h2 ? valid_0_1 : _GEN_1513; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1770 = unuse_way == 3'h2 ? valid_0_2 : _GEN_1514; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1771 = unuse_way == 3'h2 ? valid_0_3 : _GEN_1515; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1772 = unuse_way == 3'h2 ? valid_0_4 : _GEN_1516; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1773 = unuse_way == 3'h2 ? valid_0_5 : _GEN_1517; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1774 = unuse_way == 3'h2 ? valid_0_6 : _GEN_1518; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1775 = unuse_way == 3'h2 ? valid_0_7 : _GEN_1519; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1776 = unuse_way == 3'h2 ? valid_0_8 : _GEN_1520; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1777 = unuse_way == 3'h2 ? valid_0_9 : _GEN_1521; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1778 = unuse_way == 3'h2 ? valid_0_10 : _GEN_1522; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1779 = unuse_way == 3'h2 ? valid_0_11 : _GEN_1523; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1780 = unuse_way == 3'h2 ? valid_0_12 : _GEN_1524; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1781 = unuse_way == 3'h2 ? valid_0_13 : _GEN_1525; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1782 = unuse_way == 3'h2 ? valid_0_14 : _GEN_1526; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1783 = unuse_way == 3'h2 ? valid_0_15 : _GEN_1527; // @[i_cache.scala 27:26 90:40]
  wire [511:0] _GEN_1784 = unuse_way == 3'h1 ? _GEN_152 : _GEN_1736; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1785 = unuse_way == 3'h1 ? _GEN_153 : _GEN_1737; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1786 = unuse_way == 3'h1 ? _GEN_154 : _GEN_1738; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1787 = unuse_way == 3'h1 ? _GEN_155 : _GEN_1739; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1788 = unuse_way == 3'h1 ? _GEN_156 : _GEN_1740; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1789 = unuse_way == 3'h1 ? _GEN_157 : _GEN_1741; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1790 = unuse_way == 3'h1 ? _GEN_158 : _GEN_1742; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1791 = unuse_way == 3'h1 ? _GEN_159 : _GEN_1743; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1792 = unuse_way == 3'h1 ? _GEN_160 : _GEN_1744; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1793 = unuse_way == 3'h1 ? _GEN_161 : _GEN_1745; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1794 = unuse_way == 3'h1 ? _GEN_162 : _GEN_1746; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1795 = unuse_way == 3'h1 ? _GEN_163 : _GEN_1747; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1796 = unuse_way == 3'h1 ? _GEN_164 : _GEN_1748; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1797 = unuse_way == 3'h1 ? _GEN_165 : _GEN_1749; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1798 = unuse_way == 3'h1 ? _GEN_166 : _GEN_1750; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1799 = unuse_way == 3'h1 ? _GEN_167 : _GEN_1751; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1800 = unuse_way == 3'h1 ? _GEN_168 : _GEN_1752; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1801 = unuse_way == 3'h1 ? _GEN_169 : _GEN_1753; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1802 = unuse_way == 3'h1 ? _GEN_170 : _GEN_1754; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1803 = unuse_way == 3'h1 ? _GEN_171 : _GEN_1755; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1804 = unuse_way == 3'h1 ? _GEN_172 : _GEN_1756; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1805 = unuse_way == 3'h1 ? _GEN_173 : _GEN_1757; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1806 = unuse_way == 3'h1 ? _GEN_174 : _GEN_1758; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1807 = unuse_way == 3'h1 ? _GEN_175 : _GEN_1759; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1808 = unuse_way == 3'h1 ? _GEN_176 : _GEN_1760; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1809 = unuse_way == 3'h1 ? _GEN_177 : _GEN_1761; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1810 = unuse_way == 3'h1 ? _GEN_178 : _GEN_1762; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1811 = unuse_way == 3'h1 ? _GEN_179 : _GEN_1763; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1812 = unuse_way == 3'h1 ? _GEN_180 : _GEN_1764; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1813 = unuse_way == 3'h1 ? _GEN_181 : _GEN_1765; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1814 = unuse_way == 3'h1 ? _GEN_182 : _GEN_1766; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1815 = unuse_way == 3'h1 ? _GEN_183 : _GEN_1767; // @[i_cache.scala 85:34]
  wire  _GEN_1816 = unuse_way == 3'h1 ? _GEN_184 : _GEN_1768; // @[i_cache.scala 85:34]
  wire  _GEN_1817 = unuse_way == 3'h1 ? _GEN_185 : _GEN_1769; // @[i_cache.scala 85:34]
  wire  _GEN_1818 = unuse_way == 3'h1 ? _GEN_186 : _GEN_1770; // @[i_cache.scala 85:34]
  wire  _GEN_1819 = unuse_way == 3'h1 ? _GEN_187 : _GEN_1771; // @[i_cache.scala 85:34]
  wire  _GEN_1820 = unuse_way == 3'h1 ? _GEN_188 : _GEN_1772; // @[i_cache.scala 85:34]
  wire  _GEN_1821 = unuse_way == 3'h1 ? _GEN_189 : _GEN_1773; // @[i_cache.scala 85:34]
  wire  _GEN_1822 = unuse_way == 3'h1 ? _GEN_190 : _GEN_1774; // @[i_cache.scala 85:34]
  wire  _GEN_1823 = unuse_way == 3'h1 ? _GEN_191 : _GEN_1775; // @[i_cache.scala 85:34]
  wire  _GEN_1824 = unuse_way == 3'h1 ? _GEN_192 : _GEN_1776; // @[i_cache.scala 85:34]
  wire  _GEN_1825 = unuse_way == 3'h1 ? _GEN_193 : _GEN_1777; // @[i_cache.scala 85:34]
  wire  _GEN_1826 = unuse_way == 3'h1 ? _GEN_194 : _GEN_1778; // @[i_cache.scala 85:34]
  wire  _GEN_1827 = unuse_way == 3'h1 ? _GEN_195 : _GEN_1779; // @[i_cache.scala 85:34]
  wire  _GEN_1828 = unuse_way == 3'h1 ? _GEN_196 : _GEN_1780; // @[i_cache.scala 85:34]
  wire  _GEN_1829 = unuse_way == 3'h1 ? _GEN_197 : _GEN_1781; // @[i_cache.scala 85:34]
  wire  _GEN_1830 = unuse_way == 3'h1 ? _GEN_198 : _GEN_1782; // @[i_cache.scala 85:34]
  wire  _GEN_1831 = unuse_way == 3'h1 ? _GEN_199 : _GEN_1783; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1832 = unuse_way == 3'h1 ? _GEN_216 : _GEN_1624; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1833 = unuse_way == 3'h1 ? _GEN_217 : _GEN_1625; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1834 = unuse_way == 3'h1 ? _GEN_218 : _GEN_1626; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1835 = unuse_way == 3'h1 ? _GEN_219 : _GEN_1627; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1836 = unuse_way == 3'h1 ? _GEN_220 : _GEN_1628; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1837 = unuse_way == 3'h1 ? _GEN_221 : _GEN_1629; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1838 = unuse_way == 3'h1 ? _GEN_222 : _GEN_1630; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1839 = unuse_way == 3'h1 ? _GEN_223 : _GEN_1631; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1840 = unuse_way == 3'h1 ? _GEN_224 : _GEN_1632; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1841 = unuse_way == 3'h1 ? _GEN_225 : _GEN_1633; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1842 = unuse_way == 3'h1 ? _GEN_226 : _GEN_1634; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1843 = unuse_way == 3'h1 ? _GEN_227 : _GEN_1635; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1844 = unuse_way == 3'h1 ? _GEN_228 : _GEN_1636; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1845 = unuse_way == 3'h1 ? _GEN_229 : _GEN_1637; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1846 = unuse_way == 3'h1 ? _GEN_230 : _GEN_1638; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1847 = unuse_way == 3'h1 ? _GEN_231 : _GEN_1639; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1848 = unuse_way == 3'h1 ? ram_1_0 : _GEN_1576; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1849 = unuse_way == 3'h1 ? ram_1_1 : _GEN_1577; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1850 = unuse_way == 3'h1 ? ram_1_2 : _GEN_1578; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1851 = unuse_way == 3'h1 ? ram_1_3 : _GEN_1579; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1852 = unuse_way == 3'h1 ? ram_1_4 : _GEN_1580; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1853 = unuse_way == 3'h1 ? ram_1_5 : _GEN_1581; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1854 = unuse_way == 3'h1 ? ram_1_6 : _GEN_1582; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1855 = unuse_way == 3'h1 ? ram_1_7 : _GEN_1583; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1856 = unuse_way == 3'h1 ? ram_1_8 : _GEN_1584; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1857 = unuse_way == 3'h1 ? ram_1_9 : _GEN_1585; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1858 = unuse_way == 3'h1 ? ram_1_10 : _GEN_1586; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1859 = unuse_way == 3'h1 ? ram_1_11 : _GEN_1587; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1860 = unuse_way == 3'h1 ? ram_1_12 : _GEN_1588; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1861 = unuse_way == 3'h1 ? ram_1_13 : _GEN_1589; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1862 = unuse_way == 3'h1 ? ram_1_14 : _GEN_1590; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1863 = unuse_way == 3'h1 ? ram_1_15 : _GEN_1591; // @[i_cache.scala 20:24 85:34]
  wire [31:0] _GEN_1864 = unuse_way == 3'h1 ? tag_1_0 : _GEN_1592; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1865 = unuse_way == 3'h1 ? tag_1_1 : _GEN_1593; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1866 = unuse_way == 3'h1 ? tag_1_2 : _GEN_1594; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1867 = unuse_way == 3'h1 ? tag_1_3 : _GEN_1595; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1868 = unuse_way == 3'h1 ? tag_1_4 : _GEN_1596; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1869 = unuse_way == 3'h1 ? tag_1_5 : _GEN_1597; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1870 = unuse_way == 3'h1 ? tag_1_6 : _GEN_1598; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1871 = unuse_way == 3'h1 ? tag_1_7 : _GEN_1599; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1872 = unuse_way == 3'h1 ? tag_1_8 : _GEN_1600; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1873 = unuse_way == 3'h1 ? tag_1_9 : _GEN_1601; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1874 = unuse_way == 3'h1 ? tag_1_10 : _GEN_1602; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1875 = unuse_way == 3'h1 ? tag_1_11 : _GEN_1603; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1876 = unuse_way == 3'h1 ? tag_1_12 : _GEN_1604; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1877 = unuse_way == 3'h1 ? tag_1_13 : _GEN_1605; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1878 = unuse_way == 3'h1 ? tag_1_14 : _GEN_1606; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1879 = unuse_way == 3'h1 ? tag_1_15 : _GEN_1607; // @[i_cache.scala 24:24 85:34]
  wire  _GEN_1880 = unuse_way == 3'h1 ? valid_1_0 : _GEN_1608; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1881 = unuse_way == 3'h1 ? valid_1_1 : _GEN_1609; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1882 = unuse_way == 3'h1 ? valid_1_2 : _GEN_1610; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1883 = unuse_way == 3'h1 ? valid_1_3 : _GEN_1611; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1884 = unuse_way == 3'h1 ? valid_1_4 : _GEN_1612; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1885 = unuse_way == 3'h1 ? valid_1_5 : _GEN_1613; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1886 = unuse_way == 3'h1 ? valid_1_6 : _GEN_1614; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1887 = unuse_way == 3'h1 ? valid_1_7 : _GEN_1615; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1888 = unuse_way == 3'h1 ? valid_1_8 : _GEN_1616; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1889 = unuse_way == 3'h1 ? valid_1_9 : _GEN_1617; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1890 = unuse_way == 3'h1 ? valid_1_10 : _GEN_1618; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1891 = unuse_way == 3'h1 ? valid_1_11 : _GEN_1619; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1892 = unuse_way == 3'h1 ? valid_1_12 : _GEN_1620; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1893 = unuse_way == 3'h1 ? valid_1_13 : _GEN_1621; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1894 = unuse_way == 3'h1 ? valid_1_14 : _GEN_1622; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1895 = unuse_way == 3'h1 ? valid_1_15 : _GEN_1623; // @[i_cache.scala 28:26 85:34]
  wire [511:0] _GEN_1896 = unuse_way == 3'h1 ? ram_2_0 : _GEN_1640; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1897 = unuse_way == 3'h1 ? ram_2_1 : _GEN_1641; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1898 = unuse_way == 3'h1 ? ram_2_2 : _GEN_1642; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1899 = unuse_way == 3'h1 ? ram_2_3 : _GEN_1643; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1900 = unuse_way == 3'h1 ? ram_2_4 : _GEN_1644; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1901 = unuse_way == 3'h1 ? ram_2_5 : _GEN_1645; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1902 = unuse_way == 3'h1 ? ram_2_6 : _GEN_1646; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1903 = unuse_way == 3'h1 ? ram_2_7 : _GEN_1647; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1904 = unuse_way == 3'h1 ? ram_2_8 : _GEN_1648; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1905 = unuse_way == 3'h1 ? ram_2_9 : _GEN_1649; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1906 = unuse_way == 3'h1 ? ram_2_10 : _GEN_1650; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1907 = unuse_way == 3'h1 ? ram_2_11 : _GEN_1651; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1908 = unuse_way == 3'h1 ? ram_2_12 : _GEN_1652; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1909 = unuse_way == 3'h1 ? ram_2_13 : _GEN_1653; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1910 = unuse_way == 3'h1 ? ram_2_14 : _GEN_1654; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1911 = unuse_way == 3'h1 ? ram_2_15 : _GEN_1655; // @[i_cache.scala 21:24 85:34]
  wire [31:0] _GEN_1912 = unuse_way == 3'h1 ? tag_2_0 : _GEN_1656; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1913 = unuse_way == 3'h1 ? tag_2_1 : _GEN_1657; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1914 = unuse_way == 3'h1 ? tag_2_2 : _GEN_1658; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1915 = unuse_way == 3'h1 ? tag_2_3 : _GEN_1659; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1916 = unuse_way == 3'h1 ? tag_2_4 : _GEN_1660; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1917 = unuse_way == 3'h1 ? tag_2_5 : _GEN_1661; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1918 = unuse_way == 3'h1 ? tag_2_6 : _GEN_1662; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1919 = unuse_way == 3'h1 ? tag_2_7 : _GEN_1663; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1920 = unuse_way == 3'h1 ? tag_2_8 : _GEN_1664; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1921 = unuse_way == 3'h1 ? tag_2_9 : _GEN_1665; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1922 = unuse_way == 3'h1 ? tag_2_10 : _GEN_1666; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1923 = unuse_way == 3'h1 ? tag_2_11 : _GEN_1667; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1924 = unuse_way == 3'h1 ? tag_2_12 : _GEN_1668; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1925 = unuse_way == 3'h1 ? tag_2_13 : _GEN_1669; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1926 = unuse_way == 3'h1 ? tag_2_14 : _GEN_1670; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1927 = unuse_way == 3'h1 ? tag_2_15 : _GEN_1671; // @[i_cache.scala 25:24 85:34]
  wire  _GEN_1928 = unuse_way == 3'h1 ? valid_2_0 : _GEN_1672; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1929 = unuse_way == 3'h1 ? valid_2_1 : _GEN_1673; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1930 = unuse_way == 3'h1 ? valid_2_2 : _GEN_1674; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1931 = unuse_way == 3'h1 ? valid_2_3 : _GEN_1675; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1932 = unuse_way == 3'h1 ? valid_2_4 : _GEN_1676; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1933 = unuse_way == 3'h1 ? valid_2_5 : _GEN_1677; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1934 = unuse_way == 3'h1 ? valid_2_6 : _GEN_1678; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1935 = unuse_way == 3'h1 ? valid_2_7 : _GEN_1679; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1936 = unuse_way == 3'h1 ? valid_2_8 : _GEN_1680; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1937 = unuse_way == 3'h1 ? valid_2_9 : _GEN_1681; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1938 = unuse_way == 3'h1 ? valid_2_10 : _GEN_1682; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1939 = unuse_way == 3'h1 ? valid_2_11 : _GEN_1683; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1940 = unuse_way == 3'h1 ? valid_2_12 : _GEN_1684; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1941 = unuse_way == 3'h1 ? valid_2_13 : _GEN_1685; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1942 = unuse_way == 3'h1 ? valid_2_14 : _GEN_1686; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1943 = unuse_way == 3'h1 ? valid_2_15 : _GEN_1687; // @[i_cache.scala 29:26 85:34]
  wire [511:0] _GEN_1944 = unuse_way == 3'h1 ? ram_3_0 : _GEN_1688; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1945 = unuse_way == 3'h1 ? ram_3_1 : _GEN_1689; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1946 = unuse_way == 3'h1 ? ram_3_2 : _GEN_1690; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1947 = unuse_way == 3'h1 ? ram_3_3 : _GEN_1691; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1948 = unuse_way == 3'h1 ? ram_3_4 : _GEN_1692; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1949 = unuse_way == 3'h1 ? ram_3_5 : _GEN_1693; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1950 = unuse_way == 3'h1 ? ram_3_6 : _GEN_1694; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1951 = unuse_way == 3'h1 ? ram_3_7 : _GEN_1695; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1952 = unuse_way == 3'h1 ? ram_3_8 : _GEN_1696; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1953 = unuse_way == 3'h1 ? ram_3_9 : _GEN_1697; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1954 = unuse_way == 3'h1 ? ram_3_10 : _GEN_1698; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1955 = unuse_way == 3'h1 ? ram_3_11 : _GEN_1699; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1956 = unuse_way == 3'h1 ? ram_3_12 : _GEN_1700; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1957 = unuse_way == 3'h1 ? ram_3_13 : _GEN_1701; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1958 = unuse_way == 3'h1 ? ram_3_14 : _GEN_1702; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1959 = unuse_way == 3'h1 ? ram_3_15 : _GEN_1703; // @[i_cache.scala 22:24 85:34]
  wire [31:0] _GEN_1960 = unuse_way == 3'h1 ? tag_3_0 : _GEN_1704; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1961 = unuse_way == 3'h1 ? tag_3_1 : _GEN_1705; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1962 = unuse_way == 3'h1 ? tag_3_2 : _GEN_1706; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1963 = unuse_way == 3'h1 ? tag_3_3 : _GEN_1707; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1964 = unuse_way == 3'h1 ? tag_3_4 : _GEN_1708; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1965 = unuse_way == 3'h1 ? tag_3_5 : _GEN_1709; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1966 = unuse_way == 3'h1 ? tag_3_6 : _GEN_1710; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1967 = unuse_way == 3'h1 ? tag_3_7 : _GEN_1711; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1968 = unuse_way == 3'h1 ? tag_3_8 : _GEN_1712; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1969 = unuse_way == 3'h1 ? tag_3_9 : _GEN_1713; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1970 = unuse_way == 3'h1 ? tag_3_10 : _GEN_1714; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1971 = unuse_way == 3'h1 ? tag_3_11 : _GEN_1715; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1972 = unuse_way == 3'h1 ? tag_3_12 : _GEN_1716; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1973 = unuse_way == 3'h1 ? tag_3_13 : _GEN_1717; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1974 = unuse_way == 3'h1 ? tag_3_14 : _GEN_1718; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1975 = unuse_way == 3'h1 ? tag_3_15 : _GEN_1719; // @[i_cache.scala 26:24 85:34]
  wire  _GEN_1976 = unuse_way == 3'h1 ? valid_3_0 : _GEN_1720; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1977 = unuse_way == 3'h1 ? valid_3_1 : _GEN_1721; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1978 = unuse_way == 3'h1 ? valid_3_2 : _GEN_1722; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1979 = unuse_way == 3'h1 ? valid_3_3 : _GEN_1723; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1980 = unuse_way == 3'h1 ? valid_3_4 : _GEN_1724; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1981 = unuse_way == 3'h1 ? valid_3_5 : _GEN_1725; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1982 = unuse_way == 3'h1 ? valid_3_6 : _GEN_1726; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1983 = unuse_way == 3'h1 ? valid_3_7 : _GEN_1727; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1984 = unuse_way == 3'h1 ? valid_3_8 : _GEN_1728; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1985 = unuse_way == 3'h1 ? valid_3_9 : _GEN_1729; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1986 = unuse_way == 3'h1 ? valid_3_10 : _GEN_1730; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1987 = unuse_way == 3'h1 ? valid_3_11 : _GEN_1731; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1988 = unuse_way == 3'h1 ? valid_3_12 : _GEN_1732; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1989 = unuse_way == 3'h1 ? valid_3_13 : _GEN_1733; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1990 = unuse_way == 3'h1 ? valid_3_14 : _GEN_1734; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1991 = unuse_way == 3'h1 ? valid_3_15 : _GEN_1735; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1992 = 3'h4 == state ? 1'h0 : valid_0_0; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1993 = 3'h4 == state ? 1'h0 : valid_0_1; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1994 = 3'h4 == state ? 1'h0 : valid_0_2; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1995 = 3'h4 == state ? 1'h0 : valid_0_3; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1996 = 3'h4 == state ? 1'h0 : valid_0_4; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1997 = 3'h4 == state ? 1'h0 : valid_0_5; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1998 = 3'h4 == state ? 1'h0 : valid_0_6; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1999 = 3'h4 == state ? 1'h0 : valid_0_7; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2000 = 3'h4 == state ? 1'h0 : valid_0_8; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2001 = 3'h4 == state ? 1'h0 : valid_0_9; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2002 = 3'h4 == state ? 1'h0 : valid_0_10; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2003 = 3'h4 == state ? 1'h0 : valid_0_11; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2004 = 3'h4 == state ? 1'h0 : valid_0_12; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2005 = 3'h4 == state ? 1'h0 : valid_0_13; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2006 = 3'h4 == state ? 1'h0 : valid_0_14; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2007 = 3'h4 == state ? 1'h0 : valid_0_15; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2008 = 3'h4 == state ? 1'h0 : valid_1_0; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2009 = 3'h4 == state ? 1'h0 : valid_1_1; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2010 = 3'h4 == state ? 1'h0 : valid_1_2; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2011 = 3'h4 == state ? 1'h0 : valid_1_3; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2012 = 3'h4 == state ? 1'h0 : valid_1_4; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2013 = 3'h4 == state ? 1'h0 : valid_1_5; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2014 = 3'h4 == state ? 1'h0 : valid_1_6; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2015 = 3'h4 == state ? 1'h0 : valid_1_7; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2016 = 3'h4 == state ? 1'h0 : valid_1_8; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2017 = 3'h4 == state ? 1'h0 : valid_1_9; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2018 = 3'h4 == state ? 1'h0 : valid_1_10; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2019 = 3'h4 == state ? 1'h0 : valid_1_11; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2020 = 3'h4 == state ? 1'h0 : valid_1_12; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2021 = 3'h4 == state ? 1'h0 : valid_1_13; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2022 = 3'h4 == state ? 1'h0 : valid_1_14; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2023 = 3'h4 == state ? 1'h0 : valid_1_15; // @[i_cache.scala 56:18 131:49 28:26]
  wire [2:0] _GEN_2024 = 3'h4 == state ? 3'h0 : state; // @[i_cache.scala 132:18 56:18 54:24]
  wire [2:0] _GEN_2025 = 3'h3 == state ? 3'h1 : _GEN_2024; // @[i_cache.scala 56:18 84:19]
  wire [511:0] _GEN_2026 = 3'h3 == state ? _GEN_1784 : ram_0_0; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2027 = 3'h3 == state ? _GEN_1785 : ram_0_1; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2028 = 3'h3 == state ? _GEN_1786 : ram_0_2; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2029 = 3'h3 == state ? _GEN_1787 : ram_0_3; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2030 = 3'h3 == state ? _GEN_1788 : ram_0_4; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2031 = 3'h3 == state ? _GEN_1789 : ram_0_5; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2032 = 3'h3 == state ? _GEN_1790 : ram_0_6; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2033 = 3'h3 == state ? _GEN_1791 : ram_0_7; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2034 = 3'h3 == state ? _GEN_1792 : ram_0_8; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2035 = 3'h3 == state ? _GEN_1793 : ram_0_9; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2036 = 3'h3 == state ? _GEN_1794 : ram_0_10; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2037 = 3'h3 == state ? _GEN_1795 : ram_0_11; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2038 = 3'h3 == state ? _GEN_1796 : ram_0_12; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2039 = 3'h3 == state ? _GEN_1797 : ram_0_13; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2040 = 3'h3 == state ? _GEN_1798 : ram_0_14; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2041 = 3'h3 == state ? _GEN_1799 : ram_0_15; // @[i_cache.scala 56:18 19:24]
  wire [31:0] _GEN_2042 = 3'h3 == state ? _GEN_1800 : tag_0_0; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2043 = 3'h3 == state ? _GEN_1801 : tag_0_1; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2044 = 3'h3 == state ? _GEN_1802 : tag_0_2; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2045 = 3'h3 == state ? _GEN_1803 : tag_0_3; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2046 = 3'h3 == state ? _GEN_1804 : tag_0_4; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2047 = 3'h3 == state ? _GEN_1805 : tag_0_5; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2048 = 3'h3 == state ? _GEN_1806 : tag_0_6; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2049 = 3'h3 == state ? _GEN_1807 : tag_0_7; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2050 = 3'h3 == state ? _GEN_1808 : tag_0_8; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2051 = 3'h3 == state ? _GEN_1809 : tag_0_9; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2052 = 3'h3 == state ? _GEN_1810 : tag_0_10; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2053 = 3'h3 == state ? _GEN_1811 : tag_0_11; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2054 = 3'h3 == state ? _GEN_1812 : tag_0_12; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2055 = 3'h3 == state ? _GEN_1813 : tag_0_13; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2056 = 3'h3 == state ? _GEN_1814 : tag_0_14; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2057 = 3'h3 == state ? _GEN_1815 : tag_0_15; // @[i_cache.scala 56:18 23:24]
  wire  _GEN_2058 = 3'h3 == state ? _GEN_1816 : _GEN_1992; // @[i_cache.scala 56:18]
  wire  _GEN_2059 = 3'h3 == state ? _GEN_1817 : _GEN_1993; // @[i_cache.scala 56:18]
  wire  _GEN_2060 = 3'h3 == state ? _GEN_1818 : _GEN_1994; // @[i_cache.scala 56:18]
  wire  _GEN_2061 = 3'h3 == state ? _GEN_1819 : _GEN_1995; // @[i_cache.scala 56:18]
  wire  _GEN_2062 = 3'h3 == state ? _GEN_1820 : _GEN_1996; // @[i_cache.scala 56:18]
  wire  _GEN_2063 = 3'h3 == state ? _GEN_1821 : _GEN_1997; // @[i_cache.scala 56:18]
  wire  _GEN_2064 = 3'h3 == state ? _GEN_1822 : _GEN_1998; // @[i_cache.scala 56:18]
  wire  _GEN_2065 = 3'h3 == state ? _GEN_1823 : _GEN_1999; // @[i_cache.scala 56:18]
  wire  _GEN_2066 = 3'h3 == state ? _GEN_1824 : _GEN_2000; // @[i_cache.scala 56:18]
  wire  _GEN_2067 = 3'h3 == state ? _GEN_1825 : _GEN_2001; // @[i_cache.scala 56:18]
  wire  _GEN_2068 = 3'h3 == state ? _GEN_1826 : _GEN_2002; // @[i_cache.scala 56:18]
  wire  _GEN_2069 = 3'h3 == state ? _GEN_1827 : _GEN_2003; // @[i_cache.scala 56:18]
  wire  _GEN_2070 = 3'h3 == state ? _GEN_1828 : _GEN_2004; // @[i_cache.scala 56:18]
  wire  _GEN_2071 = 3'h3 == state ? _GEN_1829 : _GEN_2005; // @[i_cache.scala 56:18]
  wire  _GEN_2072 = 3'h3 == state ? _GEN_1830 : _GEN_2006; // @[i_cache.scala 56:18]
  wire  _GEN_2073 = 3'h3 == state ? _GEN_1831 : _GEN_2007; // @[i_cache.scala 56:18]
  wire [7:0] _GEN_2074 = 3'h3 == state ? _GEN_1832 : quene_0; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2075 = 3'h3 == state ? _GEN_1833 : quene_1; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2076 = 3'h3 == state ? _GEN_1834 : quene_2; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2077 = 3'h3 == state ? _GEN_1835 : quene_3; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2078 = 3'h3 == state ? _GEN_1836 : quene_4; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2079 = 3'h3 == state ? _GEN_1837 : quene_5; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2080 = 3'h3 == state ? _GEN_1838 : quene_6; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2081 = 3'h3 == state ? _GEN_1839 : quene_7; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2082 = 3'h3 == state ? _GEN_1840 : quene_8; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2083 = 3'h3 == state ? _GEN_1841 : quene_9; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2084 = 3'h3 == state ? _GEN_1842 : quene_10; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2085 = 3'h3 == state ? _GEN_1843 : quene_11; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2086 = 3'h3 == state ? _GEN_1844 : quene_12; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2087 = 3'h3 == state ? _GEN_1845 : quene_13; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2088 = 3'h3 == state ? _GEN_1846 : quene_14; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2089 = 3'h3 == state ? _GEN_1847 : quene_15; // @[i_cache.scala 56:18 40:24]
  wire [511:0] _GEN_2090 = 3'h3 == state ? _GEN_1848 : ram_1_0; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2091 = 3'h3 == state ? _GEN_1849 : ram_1_1; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2092 = 3'h3 == state ? _GEN_1850 : ram_1_2; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2093 = 3'h3 == state ? _GEN_1851 : ram_1_3; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2094 = 3'h3 == state ? _GEN_1852 : ram_1_4; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2095 = 3'h3 == state ? _GEN_1853 : ram_1_5; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2096 = 3'h3 == state ? _GEN_1854 : ram_1_6; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2097 = 3'h3 == state ? _GEN_1855 : ram_1_7; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2098 = 3'h3 == state ? _GEN_1856 : ram_1_8; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2099 = 3'h3 == state ? _GEN_1857 : ram_1_9; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2100 = 3'h3 == state ? _GEN_1858 : ram_1_10; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2101 = 3'h3 == state ? _GEN_1859 : ram_1_11; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2102 = 3'h3 == state ? _GEN_1860 : ram_1_12; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2103 = 3'h3 == state ? _GEN_1861 : ram_1_13; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2104 = 3'h3 == state ? _GEN_1862 : ram_1_14; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2105 = 3'h3 == state ? _GEN_1863 : ram_1_15; // @[i_cache.scala 56:18 20:24]
  wire [31:0] _GEN_2106 = 3'h3 == state ? _GEN_1864 : tag_1_0; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2107 = 3'h3 == state ? _GEN_1865 : tag_1_1; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2108 = 3'h3 == state ? _GEN_1866 : tag_1_2; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2109 = 3'h3 == state ? _GEN_1867 : tag_1_3; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2110 = 3'h3 == state ? _GEN_1868 : tag_1_4; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2111 = 3'h3 == state ? _GEN_1869 : tag_1_5; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2112 = 3'h3 == state ? _GEN_1870 : tag_1_6; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2113 = 3'h3 == state ? _GEN_1871 : tag_1_7; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2114 = 3'h3 == state ? _GEN_1872 : tag_1_8; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2115 = 3'h3 == state ? _GEN_1873 : tag_1_9; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2116 = 3'h3 == state ? _GEN_1874 : tag_1_10; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2117 = 3'h3 == state ? _GEN_1875 : tag_1_11; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2118 = 3'h3 == state ? _GEN_1876 : tag_1_12; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2119 = 3'h3 == state ? _GEN_1877 : tag_1_13; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2120 = 3'h3 == state ? _GEN_1878 : tag_1_14; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2121 = 3'h3 == state ? _GEN_1879 : tag_1_15; // @[i_cache.scala 56:18 24:24]
  wire  _GEN_2122 = 3'h3 == state ? _GEN_1880 : _GEN_2008; // @[i_cache.scala 56:18]
  wire  _GEN_2123 = 3'h3 == state ? _GEN_1881 : _GEN_2009; // @[i_cache.scala 56:18]
  wire  _GEN_2124 = 3'h3 == state ? _GEN_1882 : _GEN_2010; // @[i_cache.scala 56:18]
  wire  _GEN_2125 = 3'h3 == state ? _GEN_1883 : _GEN_2011; // @[i_cache.scala 56:18]
  wire  _GEN_2126 = 3'h3 == state ? _GEN_1884 : _GEN_2012; // @[i_cache.scala 56:18]
  wire  _GEN_2127 = 3'h3 == state ? _GEN_1885 : _GEN_2013; // @[i_cache.scala 56:18]
  wire  _GEN_2128 = 3'h3 == state ? _GEN_1886 : _GEN_2014; // @[i_cache.scala 56:18]
  wire  _GEN_2129 = 3'h3 == state ? _GEN_1887 : _GEN_2015; // @[i_cache.scala 56:18]
  wire  _GEN_2130 = 3'h3 == state ? _GEN_1888 : _GEN_2016; // @[i_cache.scala 56:18]
  wire  _GEN_2131 = 3'h3 == state ? _GEN_1889 : _GEN_2017; // @[i_cache.scala 56:18]
  wire  _GEN_2132 = 3'h3 == state ? _GEN_1890 : _GEN_2018; // @[i_cache.scala 56:18]
  wire  _GEN_2133 = 3'h3 == state ? _GEN_1891 : _GEN_2019; // @[i_cache.scala 56:18]
  wire  _GEN_2134 = 3'h3 == state ? _GEN_1892 : _GEN_2020; // @[i_cache.scala 56:18]
  wire  _GEN_2135 = 3'h3 == state ? _GEN_1893 : _GEN_2021; // @[i_cache.scala 56:18]
  wire  _GEN_2136 = 3'h3 == state ? _GEN_1894 : _GEN_2022; // @[i_cache.scala 56:18]
  wire  _GEN_2137 = 3'h3 == state ? _GEN_1895 : _GEN_2023; // @[i_cache.scala 56:18]
  wire [511:0] _GEN_2138 = 3'h3 == state ? _GEN_1896 : ram_2_0; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2139 = 3'h3 == state ? _GEN_1897 : ram_2_1; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2140 = 3'h3 == state ? _GEN_1898 : ram_2_2; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2141 = 3'h3 == state ? _GEN_1899 : ram_2_3; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2142 = 3'h3 == state ? _GEN_1900 : ram_2_4; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2143 = 3'h3 == state ? _GEN_1901 : ram_2_5; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2144 = 3'h3 == state ? _GEN_1902 : ram_2_6; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2145 = 3'h3 == state ? _GEN_1903 : ram_2_7; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2146 = 3'h3 == state ? _GEN_1904 : ram_2_8; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2147 = 3'h3 == state ? _GEN_1905 : ram_2_9; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2148 = 3'h3 == state ? _GEN_1906 : ram_2_10; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2149 = 3'h3 == state ? _GEN_1907 : ram_2_11; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2150 = 3'h3 == state ? _GEN_1908 : ram_2_12; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2151 = 3'h3 == state ? _GEN_1909 : ram_2_13; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2152 = 3'h3 == state ? _GEN_1910 : ram_2_14; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2153 = 3'h3 == state ? _GEN_1911 : ram_2_15; // @[i_cache.scala 56:18 21:24]
  wire [31:0] _GEN_2154 = 3'h3 == state ? _GEN_1912 : tag_2_0; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2155 = 3'h3 == state ? _GEN_1913 : tag_2_1; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2156 = 3'h3 == state ? _GEN_1914 : tag_2_2; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2157 = 3'h3 == state ? _GEN_1915 : tag_2_3; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2158 = 3'h3 == state ? _GEN_1916 : tag_2_4; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2159 = 3'h3 == state ? _GEN_1917 : tag_2_5; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2160 = 3'h3 == state ? _GEN_1918 : tag_2_6; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2161 = 3'h3 == state ? _GEN_1919 : tag_2_7; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2162 = 3'h3 == state ? _GEN_1920 : tag_2_8; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2163 = 3'h3 == state ? _GEN_1921 : tag_2_9; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2164 = 3'h3 == state ? _GEN_1922 : tag_2_10; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2165 = 3'h3 == state ? _GEN_1923 : tag_2_11; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2166 = 3'h3 == state ? _GEN_1924 : tag_2_12; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2167 = 3'h3 == state ? _GEN_1925 : tag_2_13; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2168 = 3'h3 == state ? _GEN_1926 : tag_2_14; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2169 = 3'h3 == state ? _GEN_1927 : tag_2_15; // @[i_cache.scala 56:18 25:24]
  wire  _GEN_2170 = 3'h3 == state ? _GEN_1928 : valid_2_0; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2171 = 3'h3 == state ? _GEN_1929 : valid_2_1; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2172 = 3'h3 == state ? _GEN_1930 : valid_2_2; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2173 = 3'h3 == state ? _GEN_1931 : valid_2_3; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2174 = 3'h3 == state ? _GEN_1932 : valid_2_4; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2175 = 3'h3 == state ? _GEN_1933 : valid_2_5; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2176 = 3'h3 == state ? _GEN_1934 : valid_2_6; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2177 = 3'h3 == state ? _GEN_1935 : valid_2_7; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2178 = 3'h3 == state ? _GEN_1936 : valid_2_8; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2179 = 3'h3 == state ? _GEN_1937 : valid_2_9; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2180 = 3'h3 == state ? _GEN_1938 : valid_2_10; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2181 = 3'h3 == state ? _GEN_1939 : valid_2_11; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2182 = 3'h3 == state ? _GEN_1940 : valid_2_12; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2183 = 3'h3 == state ? _GEN_1941 : valid_2_13; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2184 = 3'h3 == state ? _GEN_1942 : valid_2_14; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2185 = 3'h3 == state ? _GEN_1943 : valid_2_15; // @[i_cache.scala 56:18 29:26]
  wire [511:0] _GEN_2186 = 3'h3 == state ? _GEN_1944 : ram_3_0; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2187 = 3'h3 == state ? _GEN_1945 : ram_3_1; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2188 = 3'h3 == state ? _GEN_1946 : ram_3_2; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2189 = 3'h3 == state ? _GEN_1947 : ram_3_3; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2190 = 3'h3 == state ? _GEN_1948 : ram_3_4; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2191 = 3'h3 == state ? _GEN_1949 : ram_3_5; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2192 = 3'h3 == state ? _GEN_1950 : ram_3_6; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2193 = 3'h3 == state ? _GEN_1951 : ram_3_7; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2194 = 3'h3 == state ? _GEN_1952 : ram_3_8; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2195 = 3'h3 == state ? _GEN_1953 : ram_3_9; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2196 = 3'h3 == state ? _GEN_1954 : ram_3_10; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2197 = 3'h3 == state ? _GEN_1955 : ram_3_11; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2198 = 3'h3 == state ? _GEN_1956 : ram_3_12; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2199 = 3'h3 == state ? _GEN_1957 : ram_3_13; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2200 = 3'h3 == state ? _GEN_1958 : ram_3_14; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2201 = 3'h3 == state ? _GEN_1959 : ram_3_15; // @[i_cache.scala 56:18 22:24]
  wire [31:0] _GEN_2202 = 3'h3 == state ? _GEN_1960 : tag_3_0; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2203 = 3'h3 == state ? _GEN_1961 : tag_3_1; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2204 = 3'h3 == state ? _GEN_1962 : tag_3_2; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2205 = 3'h3 == state ? _GEN_1963 : tag_3_3; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2206 = 3'h3 == state ? _GEN_1964 : tag_3_4; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2207 = 3'h3 == state ? _GEN_1965 : tag_3_5; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2208 = 3'h3 == state ? _GEN_1966 : tag_3_6; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2209 = 3'h3 == state ? _GEN_1967 : tag_3_7; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2210 = 3'h3 == state ? _GEN_1968 : tag_3_8; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2211 = 3'h3 == state ? _GEN_1969 : tag_3_9; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2212 = 3'h3 == state ? _GEN_1970 : tag_3_10; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2213 = 3'h3 == state ? _GEN_1971 : tag_3_11; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2214 = 3'h3 == state ? _GEN_1972 : tag_3_12; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2215 = 3'h3 == state ? _GEN_1973 : tag_3_13; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2216 = 3'h3 == state ? _GEN_1974 : tag_3_14; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2217 = 3'h3 == state ? _GEN_1975 : tag_3_15; // @[i_cache.scala 56:18 26:24]
  wire  _GEN_2218 = 3'h3 == state ? _GEN_1976 : valid_3_0; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2219 = 3'h3 == state ? _GEN_1977 : valid_3_1; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2220 = 3'h3 == state ? _GEN_1978 : valid_3_2; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2221 = 3'h3 == state ? _GEN_1979 : valid_3_3; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2222 = 3'h3 == state ? _GEN_1980 : valid_3_4; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2223 = 3'h3 == state ? _GEN_1981 : valid_3_5; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2224 = 3'h3 == state ? _GEN_1982 : valid_3_6; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2225 = 3'h3 == state ? _GEN_1983 : valid_3_7; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2226 = 3'h3 == state ? _GEN_1984 : valid_3_8; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2227 = 3'h3 == state ? _GEN_1985 : valid_3_9; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2228 = 3'h3 == state ? _GEN_1986 : valid_3_10; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2229 = 3'h3 == state ? _GEN_1987 : valid_3_11; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2230 = 3'h3 == state ? _GEN_1988 : valid_3_12; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2231 = 3'h3 == state ? _GEN_1989 : valid_3_13; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2232 = 3'h3 == state ? _GEN_1990 : valid_3_14; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2233 = 3'h3 == state ? _GEN_1991 : valid_3_15; // @[i_cache.scala 56:18 30:26]
  wire [511:0] _GEN_2889 = 4'h1 == index ? ram_0_1 : ram_0_0; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2890 = 4'h2 == index ? ram_0_2 : _GEN_2889; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2891 = 4'h3 == index ? ram_0_3 : _GEN_2890; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2892 = 4'h4 == index ? ram_0_4 : _GEN_2891; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2893 = 4'h5 == index ? ram_0_5 : _GEN_2892; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2894 = 4'h6 == index ? ram_0_6 : _GEN_2893; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2895 = 4'h7 == index ? ram_0_7 : _GEN_2894; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2896 = 4'h8 == index ? ram_0_8 : _GEN_2895; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2897 = 4'h9 == index ? ram_0_9 : _GEN_2896; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2898 = 4'ha == index ? ram_0_10 : _GEN_2897; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2899 = 4'hb == index ? ram_0_11 : _GEN_2898; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2900 = 4'hc == index ? ram_0_12 : _GEN_2899; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2901 = 4'hd == index ? ram_0_13 : _GEN_2900; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2902 = 4'he == index ? ram_0_14 : _GEN_2901; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2903 = 4'hf == index ? ram_0_15 : _GEN_2902; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _io_to_ifu_rdata_T = _GEN_2903 >> shift_bit; // @[i_cache.scala 153:55]
  wire [511:0] _GEN_2905 = 4'h1 == index ? ram_1_1 : ram_1_0; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2906 = 4'h2 == index ? ram_1_2 : _GEN_2905; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2907 = 4'h3 == index ? ram_1_3 : _GEN_2906; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2908 = 4'h4 == index ? ram_1_4 : _GEN_2907; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2909 = 4'h5 == index ? ram_1_5 : _GEN_2908; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2910 = 4'h6 == index ? ram_1_6 : _GEN_2909; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2911 = 4'h7 == index ? ram_1_7 : _GEN_2910; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2912 = 4'h8 == index ? ram_1_8 : _GEN_2911; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2913 = 4'h9 == index ? ram_1_9 : _GEN_2912; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2914 = 4'ha == index ? ram_1_10 : _GEN_2913; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2915 = 4'hb == index ? ram_1_11 : _GEN_2914; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2916 = 4'hc == index ? ram_1_12 : _GEN_2915; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2917 = 4'hd == index ? ram_1_13 : _GEN_2916; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2918 = 4'he == index ? ram_1_14 : _GEN_2917; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2919 = 4'hf == index ? ram_1_15 : _GEN_2918; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _io_to_ifu_rdata_T_1 = _GEN_2919 >> shift_bit; // @[i_cache.scala 153:95]
  wire [511:0] _GEN_2921 = 4'h1 == index ? ram_2_1 : ram_2_0; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2922 = 4'h2 == index ? ram_2_2 : _GEN_2921; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2923 = 4'h3 == index ? ram_2_3 : _GEN_2922; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2924 = 4'h4 == index ? ram_2_4 : _GEN_2923; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2925 = 4'h5 == index ? ram_2_5 : _GEN_2924; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2926 = 4'h6 == index ? ram_2_6 : _GEN_2925; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2927 = 4'h7 == index ? ram_2_7 : _GEN_2926; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2928 = 4'h8 == index ? ram_2_8 : _GEN_2927; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2929 = 4'h9 == index ? ram_2_9 : _GEN_2928; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2930 = 4'ha == index ? ram_2_10 : _GEN_2929; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2931 = 4'hb == index ? ram_2_11 : _GEN_2930; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2932 = 4'hc == index ? ram_2_12 : _GEN_2931; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2933 = 4'hd == index ? ram_2_13 : _GEN_2932; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2934 = 4'he == index ? ram_2_14 : _GEN_2933; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2935 = 4'hf == index ? ram_2_15 : _GEN_2934; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _io_to_ifu_rdata_T_2 = _GEN_2935 >> shift_bit; // @[i_cache.scala 153:135]
  wire [511:0] _GEN_2937 = 4'h1 == index ? ram_3_1 : ram_3_0; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2938 = 4'h2 == index ? ram_3_2 : _GEN_2937; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2939 = 4'h3 == index ? ram_3_3 : _GEN_2938; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2940 = 4'h4 == index ? ram_3_4 : _GEN_2939; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2941 = 4'h5 == index ? ram_3_5 : _GEN_2940; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2942 = 4'h6 == index ? ram_3_6 : _GEN_2941; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2943 = 4'h7 == index ? ram_3_7 : _GEN_2942; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2944 = 4'h8 == index ? ram_3_8 : _GEN_2943; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2945 = 4'h9 == index ? ram_3_9 : _GEN_2944; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2946 = 4'ha == index ? ram_3_10 : _GEN_2945; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2947 = 4'hb == index ? ram_3_11 : _GEN_2946; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2948 = 4'hc == index ? ram_3_12 : _GEN_2947; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2949 = 4'hd == index ? ram_3_13 : _GEN_2948; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2950 = 4'he == index ? ram_3_14 : _GEN_2949; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2951 = 4'hf == index ? ram_3_15 : _GEN_2950; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _io_to_ifu_rdata_T_3 = _GEN_2951 >> shift_bit; // @[i_cache.scala 153:162]
  wire [511:0] _io_to_ifu_rdata_T_4 = way2_hit ? _io_to_ifu_rdata_T_2 : _io_to_ifu_rdata_T_3; // @[i_cache.scala 153:112]
  wire [511:0] _io_to_ifu_rdata_T_5 = way1_hit ? _io_to_ifu_rdata_T_1 : _io_to_ifu_rdata_T_4; // @[i_cache.scala 153:72]
  wire [511:0] _io_to_ifu_rdata_T_6 = way0_hit ? _io_to_ifu_rdata_T : _io_to_ifu_rdata_T_5; // @[i_cache.scala 153:32]
  wire  _T_19 = state == 3'h2; // @[i_cache.scala 160:21]
  wire [63:0] _GEN_3105 = {{32'd0}, io_from_ifu_araddr}; // @[i_cache.scala 169:49]
  wire [63:0] _io_to_axi_araddr_T = _GEN_3105 & 64'hffffffffffffffc0; // @[i_cache.scala 169:49]
  wire [63:0] _GEN_2954 = state == 3'h2 ? _io_to_axi_araddr_T : {{32'd0}, io_from_ifu_araddr}; // @[i_cache.scala 160:29 169:26 193:26]
  wire [2:0] _GEN_2955 = state == 3'h2 ? 3'h7 : 3'h0; // @[i_cache.scala 160:29 170:25 195:25]
  wire [63:0] _GEN_2959 = state == 3'h1 ? {{32'd0}, io_from_ifu_araddr} : _GEN_2954; // @[i_cache.scala 136:25 138:26]
  wire [2:0] _GEN_2960 = state == 3'h1 ? 3'h0 : _GEN_2955; // @[i_cache.scala 136:25 139:25]
  wire [511:0] _GEN_2964 = state == 3'h1 ? _io_to_ifu_rdata_T_6 : 512'h0; // @[i_cache.scala 136:25 153:25]
  assign io_to_ifu_rdata = _GEN_2964[63:0];
  assign io_to_ifu_rlast = state == 3'h1 & _T_4; // @[i_cache.scala 136:25 156:25]
  assign io_to_ifu_rvalid = state == 3'h1 & _T_4; // @[i_cache.scala 136:25 155:26]
  assign io_to_axi_araddr = _GEN_2959[31:0];
  assign io_to_axi_arlen = {{5'd0}, _GEN_2960};
  assign io_to_axi_arvalid = state == 3'h1 ? 1'h0 : _T_19; // @[i_cache.scala 136:25 137:27]
  assign io_to_axi_rready = state == 3'h1 ? 1'h0 : io_from_ifu_rready; // @[i_cache.scala 136:25 142:26]
  assign io_cache_init = state == 3'h4; // @[i_cache.scala 209:27]
  always @(posedge clock) begin
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_0 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_0 <= _GEN_2026;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_1 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_1 <= _GEN_2027;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_2 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_2 <= _GEN_2028;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_3 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_3 <= _GEN_2029;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_4 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_4 <= _GEN_2030;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_5 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_5 <= _GEN_2031;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_6 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_6 <= _GEN_2032;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_7 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_7 <= _GEN_2033;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_8 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_8 <= _GEN_2034;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_9 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_9 <= _GEN_2035;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_10 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_10 <= _GEN_2036;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_11 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_11 <= _GEN_2037;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_12 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_12 <= _GEN_2038;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_13 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_13 <= _GEN_2039;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_14 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_14 <= _GEN_2040;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_15 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_15 <= _GEN_2041;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_0 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_0 <= _GEN_2090;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_1 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_1 <= _GEN_2091;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_2 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_2 <= _GEN_2092;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_3 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_3 <= _GEN_2093;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_4 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_4 <= _GEN_2094;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_5 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_5 <= _GEN_2095;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_6 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_6 <= _GEN_2096;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_7 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_7 <= _GEN_2097;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_8 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_8 <= _GEN_2098;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_9 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_9 <= _GEN_2099;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_10 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_10 <= _GEN_2100;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_11 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_11 <= _GEN_2101;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_12 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_12 <= _GEN_2102;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_13 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_13 <= _GEN_2103;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_14 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_14 <= _GEN_2104;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_15 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_15 <= _GEN_2105;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_0 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_0 <= _GEN_2138;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_1 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_1 <= _GEN_2139;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_2 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_2 <= _GEN_2140;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_3 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_3 <= _GEN_2141;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_4 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_4 <= _GEN_2142;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_5 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_5 <= _GEN_2143;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_6 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_6 <= _GEN_2144;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_7 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_7 <= _GEN_2145;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_8 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_8 <= _GEN_2146;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_9 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_9 <= _GEN_2147;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_10 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_10 <= _GEN_2148;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_11 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_11 <= _GEN_2149;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_12 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_12 <= _GEN_2150;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_13 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_13 <= _GEN_2151;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_14 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_14 <= _GEN_2152;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_15 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_15 <= _GEN_2153;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_0 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_0 <= _GEN_2186;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_1 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_1 <= _GEN_2187;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_2 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_2 <= _GEN_2188;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_3 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_3 <= _GEN_2189;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_4 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_4 <= _GEN_2190;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_5 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_5 <= _GEN_2191;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_6 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_6 <= _GEN_2192;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_7 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_7 <= _GEN_2193;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_8 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_8 <= _GEN_2194;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_9 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_9 <= _GEN_2195;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_10 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_10 <= _GEN_2196;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_11 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_11 <= _GEN_2197;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_12 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_12 <= _GEN_2198;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_13 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_13 <= _GEN_2199;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_14 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_14 <= _GEN_2200;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_15 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_15 <= _GEN_2201;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_0 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_0 <= _GEN_2042;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_1 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_1 <= _GEN_2043;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_2 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_2 <= _GEN_2044;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_3 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_3 <= _GEN_2045;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_4 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_4 <= _GEN_2046;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_5 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_5 <= _GEN_2047;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_6 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_6 <= _GEN_2048;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_7 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_7 <= _GEN_2049;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_8 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_8 <= _GEN_2050;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_9 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_9 <= _GEN_2051;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_10 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_10 <= _GEN_2052;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_11 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_11 <= _GEN_2053;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_12 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_12 <= _GEN_2054;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_13 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_13 <= _GEN_2055;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_14 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_14 <= _GEN_2056;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_15 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_15 <= _GEN_2057;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_0 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_0 <= _GEN_2106;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_1 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_1 <= _GEN_2107;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_2 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_2 <= _GEN_2108;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_3 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_3 <= _GEN_2109;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_4 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_4 <= _GEN_2110;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_5 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_5 <= _GEN_2111;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_6 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_6 <= _GEN_2112;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_7 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_7 <= _GEN_2113;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_8 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_8 <= _GEN_2114;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_9 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_9 <= _GEN_2115;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_10 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_10 <= _GEN_2116;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_11 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_11 <= _GEN_2117;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_12 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_12 <= _GEN_2118;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_13 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_13 <= _GEN_2119;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_14 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_14 <= _GEN_2120;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_15 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_15 <= _GEN_2121;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_0 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_0 <= _GEN_2154;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_1 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_1 <= _GEN_2155;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_2 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_2 <= _GEN_2156;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_3 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_3 <= _GEN_2157;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_4 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_4 <= _GEN_2158;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_5 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_5 <= _GEN_2159;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_6 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_6 <= _GEN_2160;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_7 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_7 <= _GEN_2161;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_8 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_8 <= _GEN_2162;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_9 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_9 <= _GEN_2163;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_10 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_10 <= _GEN_2164;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_11 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_11 <= _GEN_2165;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_12 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_12 <= _GEN_2166;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_13 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_13 <= _GEN_2167;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_14 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_14 <= _GEN_2168;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_15 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_15 <= _GEN_2169;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_0 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_0 <= _GEN_2202;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_1 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_1 <= _GEN_2203;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_2 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_2 <= _GEN_2204;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_3 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_3 <= _GEN_2205;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_4 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_4 <= _GEN_2206;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_5 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_5 <= _GEN_2207;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_6 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_6 <= _GEN_2208;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_7 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_7 <= _GEN_2209;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_8 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_8 <= _GEN_2210;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_9 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_9 <= _GEN_2211;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_10 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_10 <= _GEN_2212;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_11 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_11 <= _GEN_2213;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_12 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_12 <= _GEN_2214;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_13 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_13 <= _GEN_2215;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_14 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_14 <= _GEN_2216;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_15 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_15 <= _GEN_2217;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_0 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_0 <= _GEN_2058;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_1 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_1 <= _GEN_2059;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_2 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_2 <= _GEN_2060;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_3 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_3 <= _GEN_2061;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_4 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_4 <= _GEN_2062;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_5 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_5 <= _GEN_2063;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_6 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_6 <= _GEN_2064;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_7 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_7 <= _GEN_2065;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_8 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_8 <= _GEN_2066;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_9 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_9 <= _GEN_2067;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_10 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_10 <= _GEN_2068;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_11 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_11 <= _GEN_2069;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_12 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_12 <= _GEN_2070;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_13 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_13 <= _GEN_2071;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_14 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_14 <= _GEN_2072;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_15 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_15 <= _GEN_2073;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_0 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_0 <= _GEN_2122;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_1 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_1 <= _GEN_2123;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_2 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_2 <= _GEN_2124;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_3 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_3 <= _GEN_2125;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_4 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_4 <= _GEN_2126;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_5 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_5 <= _GEN_2127;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_6 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_6 <= _GEN_2128;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_7 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_7 <= _GEN_2129;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_8 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_8 <= _GEN_2130;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_9 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_9 <= _GEN_2131;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_10 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_10 <= _GEN_2132;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_11 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_11 <= _GEN_2133;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_12 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_12 <= _GEN_2134;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_13 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_13 <= _GEN_2135;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_14 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_14 <= _GEN_2136;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_15 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_15 <= _GEN_2137;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_0 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_0 <= _GEN_2170;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_1 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_1 <= _GEN_2171;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_2 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_2 <= _GEN_2172;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_3 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_3 <= _GEN_2173;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_4 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_4 <= _GEN_2174;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_5 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_5 <= _GEN_2175;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_6 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_6 <= _GEN_2176;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_7 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_7 <= _GEN_2177;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_8 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_8 <= _GEN_2178;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_9 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_9 <= _GEN_2179;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_10 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_10 <= _GEN_2180;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_11 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_11 <= _GEN_2181;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_12 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_12 <= _GEN_2182;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_13 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_13 <= _GEN_2183;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_14 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_14 <= _GEN_2184;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_15 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_15 <= _GEN_2185;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_0 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_0 <= _GEN_2218;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_1 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_1 <= _GEN_2219;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_2 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_2 <= _GEN_2220;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_3 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_3 <= _GEN_2221;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_4 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_4 <= _GEN_2222;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_5 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_5 <= _GEN_2223;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_6 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_6 <= _GEN_2224;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_7 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_7 <= _GEN_2225;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_8 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_8 <= _GEN_2226;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_9 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_9 <= _GEN_2227;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_10 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_10 <= _GEN_2228;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_11 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_11 <= _GEN_2229;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_12 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_12 <= _GEN_2230;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_13 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_13 <= _GEN_2231;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_14 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_14 <= _GEN_2232;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_15 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_15 <= _GEN_2233;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_0 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_0 <= _GEN_142;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_1 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_1 <= _GEN_143;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_2 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_2 <= _GEN_144;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_3 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_3 <= _GEN_145;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_4 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_4 <= _GEN_146;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_5 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_5 <= _GEN_147;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_6 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_6 <= _GEN_148;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_7 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_7 <= _GEN_149;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 39:30]
      receive_num <= 3'h0; // @[i_cache.scala 39:30]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (3'h1 == state) begin // @[i_cache.scala 56:18]
        if (!(way0_hit | way1_hit | way2_hit | way3_hit)) begin // @[i_cache.scala 65:57]
          receive_num <= 3'h0; // @[i_cache.scala 71:29]
        end
      end else if (3'h2 == state) begin // @[i_cache.scala 56:18]
        receive_num <= _GEN_150;
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_0 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_0 <= _GEN_2074;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_1 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_1 <= _GEN_2075;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_2 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_2 <= _GEN_2076;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_3 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_3 <= _GEN_2077;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_4 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_4 <= _GEN_2078;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_5 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_5 <= _GEN_2079;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_6 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_6 <= _GEN_2080;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_7 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_7 <= _GEN_2081;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_8 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_8 <= _GEN_2082;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_9 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_9 <= _GEN_2083;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_10 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_10 <= _GEN_2084;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_11 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_11 <= _GEN_2085;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_12 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_12 <= _GEN_2086;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_13 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_13 <= _GEN_2087;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_14 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_14 <= _GEN_2088;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_15 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_15 <= _GEN_2089;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 54:24]
      state <= 3'h0; // @[i_cache.scala 54:24]
    end else if (3'h0 == state) begin // @[i_cache.scala 56:18]
      if (io_clear_cache) begin // @[i_cache.scala 58:33]
        state <= 3'h4; // @[i_cache.scala 59:23]
      end else if (io_from_ifu_arvalid) begin // @[i_cache.scala 60:44]
        state <= 3'h1; // @[i_cache.scala 61:23]
      end
    end else if (3'h1 == state) begin // @[i_cache.scala 56:18]
      if (way0_hit | way1_hit | way2_hit | way3_hit) begin // @[i_cache.scala 65:57]
        state <= _GEN_130;
      end else begin
        state <= 3'h2; // @[i_cache.scala 70:23]
      end
    end else if (3'h2 == state) begin // @[i_cache.scala 56:18]
      state <= _GEN_151;
    end else begin
      state <= _GEN_2025;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  ram_0_0 = _RAND_0[511:0];
  _RAND_1 = {16{`RANDOM}};
  ram_0_1 = _RAND_1[511:0];
  _RAND_2 = {16{`RANDOM}};
  ram_0_2 = _RAND_2[511:0];
  _RAND_3 = {16{`RANDOM}};
  ram_0_3 = _RAND_3[511:0];
  _RAND_4 = {16{`RANDOM}};
  ram_0_4 = _RAND_4[511:0];
  _RAND_5 = {16{`RANDOM}};
  ram_0_5 = _RAND_5[511:0];
  _RAND_6 = {16{`RANDOM}};
  ram_0_6 = _RAND_6[511:0];
  _RAND_7 = {16{`RANDOM}};
  ram_0_7 = _RAND_7[511:0];
  _RAND_8 = {16{`RANDOM}};
  ram_0_8 = _RAND_8[511:0];
  _RAND_9 = {16{`RANDOM}};
  ram_0_9 = _RAND_9[511:0];
  _RAND_10 = {16{`RANDOM}};
  ram_0_10 = _RAND_10[511:0];
  _RAND_11 = {16{`RANDOM}};
  ram_0_11 = _RAND_11[511:0];
  _RAND_12 = {16{`RANDOM}};
  ram_0_12 = _RAND_12[511:0];
  _RAND_13 = {16{`RANDOM}};
  ram_0_13 = _RAND_13[511:0];
  _RAND_14 = {16{`RANDOM}};
  ram_0_14 = _RAND_14[511:0];
  _RAND_15 = {16{`RANDOM}};
  ram_0_15 = _RAND_15[511:0];
  _RAND_16 = {16{`RANDOM}};
  ram_1_0 = _RAND_16[511:0];
  _RAND_17 = {16{`RANDOM}};
  ram_1_1 = _RAND_17[511:0];
  _RAND_18 = {16{`RANDOM}};
  ram_1_2 = _RAND_18[511:0];
  _RAND_19 = {16{`RANDOM}};
  ram_1_3 = _RAND_19[511:0];
  _RAND_20 = {16{`RANDOM}};
  ram_1_4 = _RAND_20[511:0];
  _RAND_21 = {16{`RANDOM}};
  ram_1_5 = _RAND_21[511:0];
  _RAND_22 = {16{`RANDOM}};
  ram_1_6 = _RAND_22[511:0];
  _RAND_23 = {16{`RANDOM}};
  ram_1_7 = _RAND_23[511:0];
  _RAND_24 = {16{`RANDOM}};
  ram_1_8 = _RAND_24[511:0];
  _RAND_25 = {16{`RANDOM}};
  ram_1_9 = _RAND_25[511:0];
  _RAND_26 = {16{`RANDOM}};
  ram_1_10 = _RAND_26[511:0];
  _RAND_27 = {16{`RANDOM}};
  ram_1_11 = _RAND_27[511:0];
  _RAND_28 = {16{`RANDOM}};
  ram_1_12 = _RAND_28[511:0];
  _RAND_29 = {16{`RANDOM}};
  ram_1_13 = _RAND_29[511:0];
  _RAND_30 = {16{`RANDOM}};
  ram_1_14 = _RAND_30[511:0];
  _RAND_31 = {16{`RANDOM}};
  ram_1_15 = _RAND_31[511:0];
  _RAND_32 = {16{`RANDOM}};
  ram_2_0 = _RAND_32[511:0];
  _RAND_33 = {16{`RANDOM}};
  ram_2_1 = _RAND_33[511:0];
  _RAND_34 = {16{`RANDOM}};
  ram_2_2 = _RAND_34[511:0];
  _RAND_35 = {16{`RANDOM}};
  ram_2_3 = _RAND_35[511:0];
  _RAND_36 = {16{`RANDOM}};
  ram_2_4 = _RAND_36[511:0];
  _RAND_37 = {16{`RANDOM}};
  ram_2_5 = _RAND_37[511:0];
  _RAND_38 = {16{`RANDOM}};
  ram_2_6 = _RAND_38[511:0];
  _RAND_39 = {16{`RANDOM}};
  ram_2_7 = _RAND_39[511:0];
  _RAND_40 = {16{`RANDOM}};
  ram_2_8 = _RAND_40[511:0];
  _RAND_41 = {16{`RANDOM}};
  ram_2_9 = _RAND_41[511:0];
  _RAND_42 = {16{`RANDOM}};
  ram_2_10 = _RAND_42[511:0];
  _RAND_43 = {16{`RANDOM}};
  ram_2_11 = _RAND_43[511:0];
  _RAND_44 = {16{`RANDOM}};
  ram_2_12 = _RAND_44[511:0];
  _RAND_45 = {16{`RANDOM}};
  ram_2_13 = _RAND_45[511:0];
  _RAND_46 = {16{`RANDOM}};
  ram_2_14 = _RAND_46[511:0];
  _RAND_47 = {16{`RANDOM}};
  ram_2_15 = _RAND_47[511:0];
  _RAND_48 = {16{`RANDOM}};
  ram_3_0 = _RAND_48[511:0];
  _RAND_49 = {16{`RANDOM}};
  ram_3_1 = _RAND_49[511:0];
  _RAND_50 = {16{`RANDOM}};
  ram_3_2 = _RAND_50[511:0];
  _RAND_51 = {16{`RANDOM}};
  ram_3_3 = _RAND_51[511:0];
  _RAND_52 = {16{`RANDOM}};
  ram_3_4 = _RAND_52[511:0];
  _RAND_53 = {16{`RANDOM}};
  ram_3_5 = _RAND_53[511:0];
  _RAND_54 = {16{`RANDOM}};
  ram_3_6 = _RAND_54[511:0];
  _RAND_55 = {16{`RANDOM}};
  ram_3_7 = _RAND_55[511:0];
  _RAND_56 = {16{`RANDOM}};
  ram_3_8 = _RAND_56[511:0];
  _RAND_57 = {16{`RANDOM}};
  ram_3_9 = _RAND_57[511:0];
  _RAND_58 = {16{`RANDOM}};
  ram_3_10 = _RAND_58[511:0];
  _RAND_59 = {16{`RANDOM}};
  ram_3_11 = _RAND_59[511:0];
  _RAND_60 = {16{`RANDOM}};
  ram_3_12 = _RAND_60[511:0];
  _RAND_61 = {16{`RANDOM}};
  ram_3_13 = _RAND_61[511:0];
  _RAND_62 = {16{`RANDOM}};
  ram_3_14 = _RAND_62[511:0];
  _RAND_63 = {16{`RANDOM}};
  ram_3_15 = _RAND_63[511:0];
  _RAND_64 = {1{`RANDOM}};
  tag_0_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  tag_0_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  tag_0_2 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  tag_0_3 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  tag_0_4 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  tag_0_5 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  tag_0_6 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  tag_0_7 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  tag_0_8 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  tag_0_9 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  tag_0_10 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  tag_0_11 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  tag_0_12 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  tag_0_13 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  tag_0_14 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  tag_0_15 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  tag_1_0 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  tag_1_1 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  tag_1_2 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  tag_1_3 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  tag_1_4 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  tag_1_5 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  tag_1_6 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  tag_1_7 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  tag_1_8 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  tag_1_9 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  tag_1_10 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  tag_1_11 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  tag_1_12 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  tag_1_13 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  tag_1_14 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  tag_1_15 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  tag_2_0 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  tag_2_1 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  tag_2_2 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  tag_2_3 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  tag_2_4 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  tag_2_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  tag_2_6 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  tag_2_7 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  tag_2_8 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  tag_2_9 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  tag_2_10 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  tag_2_11 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  tag_2_12 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  tag_2_13 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  tag_2_14 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  tag_2_15 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  tag_3_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  tag_3_1 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  tag_3_2 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  tag_3_3 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  tag_3_4 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  tag_3_5 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  tag_3_6 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  tag_3_7 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  tag_3_8 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  tag_3_9 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  tag_3_10 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  tag_3_11 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  tag_3_12 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  tag_3_13 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  tag_3_14 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  tag_3_15 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  valid_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_0_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_0_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_0_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_0_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_0_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_0_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_0_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_0_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_0_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_0_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_0_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_0_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_0_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_0_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_1_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_1_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_1_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_1_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_1_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_1_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_1_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_1_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_1_8 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_1_9 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_1_10 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_1_11 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_1_12 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_1_13 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_1_14 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_1_15 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_2_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_2_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_2_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_2_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_2_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_2_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_2_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_2_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_2_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_2_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_2_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_2_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_2_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_2_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_2_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_2_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_3_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_3_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_3_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_3_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_3_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_3_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_3_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_3_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_3_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_3_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_3_10 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_3_11 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_3_12 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_3_13 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_3_14 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_3_15 = _RAND_191[0:0];
  _RAND_192 = {2{`RANDOM}};
  receive_data_0 = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  receive_data_1 = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  receive_data_2 = _RAND_194[63:0];
  _RAND_195 = {2{`RANDOM}};
  receive_data_3 = _RAND_195[63:0];
  _RAND_196 = {2{`RANDOM}};
  receive_data_4 = _RAND_196[63:0];
  _RAND_197 = {2{`RANDOM}};
  receive_data_5 = _RAND_197[63:0];
  _RAND_198 = {2{`RANDOM}};
  receive_data_6 = _RAND_198[63:0];
  _RAND_199 = {2{`RANDOM}};
  receive_data_7 = _RAND_199[63:0];
  _RAND_200 = {1{`RANDOM}};
  receive_num = _RAND_200[2:0];
  _RAND_201 = {1{`RANDOM}};
  quene_0 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  quene_1 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  quene_2 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  quene_3 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  quene_4 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  quene_5 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  quene_6 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  quene_7 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  quene_8 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  quene_9 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  quene_10 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  quene_11 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  quene_12 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  quene_13 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  quene_14 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  quene_15 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  state = _RAND_217[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
