module AXI(
  input         clock,
  input         reset,
  input  [31:0] io_axi_in_araddr,
  input         io_axi_in_arvalid,
  input         io_axi_in_rready,
  input  [31:0] io_axi_in_awaddr,
  input         io_axi_in_awvalid,
  input  [31:0] io_axi_in_wdata,
  input  [7:0]  io_axi_in_wstrb,
  input         io_axi_in_wvalid,
  input         io_axi_in_bready,
  output        io_axi_out_arready,
  output [63:0] io_axi_out_rdata,
  output        io_axi_out_rvalid,
  output        io_axi_out_awready,
  output        io_axi_out_wready,
  output        io_axi_out_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] Mem_modle_Raddr; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Rdata; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Waddr; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Wdata; // @[AXI.scala 26:27]
  wire [7:0] Mem_modle_Wmask; // @[AXI.scala 26:27]
  wire  Mem_modle_Write_en; // @[AXI.scala 26:27]
  wire  Mem_modle_Read_en; // @[AXI.scala 26:27]
  reg  axi_awready; // @[AXI.scala 13:30]
  reg  axi_wready; // @[AXI.scala 14:29]
  reg  axi_bvalid; // @[AXI.scala 17:29]
  reg  axi_arready; // @[AXI.scala 19:30]
  reg  axi_rvalid; // @[AXI.scala 21:29]
  reg [2:0] state; // @[AXI.scala 24:24]
  wire  _GEN_1 = io_axi_in_arvalid ? 1'h0 : axi_arready; // @[AXI.scala 49:42 51:29 19:30]
  wire  _GEN_2 = io_axi_in_arvalid | axi_rvalid; // @[AXI.scala 49:42 52:28 21:29]
  wire  _GEN_4 = io_axi_in_awvalid & io_axi_in_wvalid ? 1'h0 : axi_awready; // @[AXI.scala 39:56 41:29 13:30]
  wire  _GEN_5 = io_axi_in_awvalid & io_axi_in_wvalid ? 1'h0 : axi_wready; // @[AXI.scala 39:56 42:28 14:29]
  wire  _GEN_6 = io_axi_in_awvalid & io_axi_in_wvalid | axi_bvalid; // @[AXI.scala 39:56 43:28 17:29]
  wire  _GEN_7 = io_axi_in_awvalid & io_axi_in_wvalid ? axi_arready : _GEN_1; // @[AXI.scala 19:30 39:56]
  wire  _GEN_11 = io_axi_in_bready | axi_awready; // @[AXI.scala 56:35 59:29 13:30]
  wire  _GEN_12 = io_axi_in_bready | axi_wready; // @[AXI.scala 56:35 60:28 14:29]
  wire [2:0] _GEN_13 = io_axi_in_rready ? 3'h0 : state; // @[AXI.scala 64:35 65:23 24:24]
  wire  _GEN_14 = io_axi_in_rready | axi_arready; // @[AXI.scala 64:35 66:29 19:30]
  wire  _GEN_15 = io_axi_in_rready ? 1'h0 : axi_rvalid; // @[AXI.scala 64:35 67:28 21:29]
  wire  _GEN_17 = 3'h4 == state ? _GEN_14 : axi_arready; // @[AXI.scala 37:18 19:30]
  wire  _GEN_21 = 3'h3 == state ? _GEN_11 : axi_awready; // @[AXI.scala 37:18 13:30]
  wire  _GEN_22 = 3'h3 == state ? _GEN_12 : axi_wready; // @[AXI.scala 37:18 14:29]
  wire  _GEN_23 = 3'h3 == state ? axi_arready : _GEN_17; // @[AXI.scala 37:18 19:30]
  wire  _GEN_26 = 3'h0 == state ? _GEN_4 : _GEN_21; // @[AXI.scala 37:18]
  wire  _GEN_27 = 3'h0 == state ? _GEN_5 : _GEN_22; // @[AXI.scala 37:18]
  wire  _GEN_29 = 3'h0 == state ? _GEN_7 : _GEN_23; // @[AXI.scala 37:18]
  MEM Mem_modle ( // @[AXI.scala 26:27]
    .Raddr(Mem_modle_Raddr),
    .Rdata(Mem_modle_Rdata),
    .Waddr(Mem_modle_Waddr),
    .Wdata(Mem_modle_Wdata),
    .Wmask(Mem_modle_Wmask),
    .Write_en(Mem_modle_Write_en),
    .Read_en(Mem_modle_Read_en)
  );
  assign io_axi_out_arready = axi_arready; // @[AXI.scala 71:24]
  assign io_axi_out_rdata = Mem_modle_Rdata; // @[AXI.scala 72:22]
  assign io_axi_out_rvalid = axi_rvalid; // @[AXI.scala 73:23]
  assign io_axi_out_awready = axi_awready; // @[AXI.scala 74:24]
  assign io_axi_out_wready = axi_wready; // @[AXI.scala 75:23]
  assign io_axi_out_bvalid = axi_bvalid; // @[AXI.scala 76:23]
  assign Mem_modle_Raddr = {32'h0,io_axi_in_araddr}; // @[Cat.scala 31:58]
  assign Mem_modle_Waddr = {{32'd0}, io_axi_in_awaddr}; // @[AXI.scala 28:24]
  assign Mem_modle_Wdata = {{32'd0}, io_axi_in_wdata}; // @[AXI.scala 29:24]
  assign Mem_modle_Wmask = io_axi_in_wstrb; // @[AXI.scala 30:24]
  assign Mem_modle_Write_en = axi_wready & io_axi_in_wvalid; // @[AXI.scala 31:48]
  assign Mem_modle_Read_en = axi_arready & io_axi_in_arvalid; // @[AXI.scala 32:48]
  always @(posedge clock) begin
    axi_awready <= reset | _GEN_26; // @[AXI.scala 13:{30,30}]
    axi_wready <= reset | _GEN_27; // @[AXI.scala 14:{29,29}]
    if (reset) begin // @[AXI.scala 17:29]
      axi_bvalid <= 1'h0; // @[AXI.scala 17:29]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      axi_bvalid <= _GEN_6;
    end else if (3'h3 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_bready) begin // @[AXI.scala 56:35]
        axi_bvalid <= 1'h0; // @[AXI.scala 58:28]
      end
    end
    axi_arready <= reset | _GEN_29; // @[AXI.scala 19:{30,30}]
    if (reset) begin // @[AXI.scala 21:29]
      axi_rvalid <= 1'h0; // @[AXI.scala 21:29]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      if (!(io_axi_in_awvalid & io_axi_in_wvalid)) begin // @[AXI.scala 39:56]
        axi_rvalid <= _GEN_2;
      end
    end else if (!(3'h3 == state)) begin // @[AXI.scala 37:18]
      if (3'h4 == state) begin // @[AXI.scala 37:18]
        axi_rvalid <= _GEN_15;
      end
    end
    if (reset) begin // @[AXI.scala 24:24]
      state <= 3'h0; // @[AXI.scala 24:24]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_awvalid & io_axi_in_wvalid) begin // @[AXI.scala 39:56]
        state <= 3'h3; // @[AXI.scala 40:23]
      end else if (io_axi_in_arvalid) begin // @[AXI.scala 49:42]
        state <= 3'h4; // @[AXI.scala 50:23]
      end
    end else if (3'h3 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_bready) begin // @[AXI.scala 56:35]
        state <= 3'h0; // @[AXI.scala 57:23]
      end
    end else if (3'h4 == state) begin // @[AXI.scala 37:18]
      state <= _GEN_13;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_awready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  axi_wready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  axi_bvalid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  axi_arready = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  axi_rvalid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSU(
  input         clock,
  input         reset,
  input         io_inst_store,
  input         io_inst_load,
  input  [31:0] io_mem_addr,
  input  [63:0] io_mem_wdata,
  input  [7:0]  io_mem_wstrb,
  output [63:0] io_mem_rdata,
  input         io_axi_in_arready,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  input         io_axi_in_awready,
  input         io_axi_in_wready,
  input         io_axi_in_bvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  output [31:0] io_axi_out_awaddr,
  output        io_axi_out_awvalid,
  output [31:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid,
  output        io_axi_out_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  axi_arvalid; // @[LSU.scala 19:30]
  reg  axi_rready; // @[LSU.scala 22:29]
  reg  axi_awvalid; // @[LSU.scala 23:30]
  reg  axi_wvalid; // @[LSU.scala 24:29]
  reg  axi_bready; // @[LSU.scala 25:29]
  reg [1:0] state; // @[LSU.scala 28:24]
  wire  _GEN_1 = io_inst_store | axi_awvalid; // @[LSU.scala 36:38 38:29 23:30]
  wire  _GEN_2 = io_inst_store | axi_wvalid; // @[LSU.scala 36:38 39:28 24:29]
  wire  _GEN_3 = io_inst_store | axi_bready; // @[LSU.scala 36:38 40:28 25:29]
  wire  _GEN_5 = io_inst_load | axi_arvalid; // @[LSU.scala 32:31 34:29 19:30]
  wire  _GEN_6 = io_inst_load | axi_rready; // @[LSU.scala 32:31 35:28 22:29]
  wire  _GEN_9 = io_inst_load ? axi_bready : _GEN_3; // @[LSU.scala 25:29 32:31]
  wire  _GEN_11 = io_axi_in_bvalid ? 1'h0 : axi_bready; // @[LSU.scala 44:35 46:28 25:29]
  wire  _GEN_14 = io_axi_in_arready ? 1'h0 : axi_arvalid; // @[LSU.scala 56:36 57:29 19:30]
  wire [1:0] _GEN_15 = io_axi_in_rvalid ? 2'h0 : state; // @[LSU.scala 59:35 60:23 28:24]
  wire  _GEN_16 = io_axi_in_rvalid ? 1'h0 : axi_rready; // @[LSU.scala 59:35 61:28 22:29]
  wire  _GEN_19 = 2'h2 == state ? _GEN_16 : axi_rready; // @[LSU.scala 30:18 22:29]
  wire  _GEN_21 = 2'h1 == state ? _GEN_11 : axi_bready; // @[LSU.scala 30:18 25:29]
  wire  _GEN_25 = 2'h1 == state ? axi_rready : _GEN_19; // @[LSU.scala 30:18 22:29]
  wire  _GEN_28 = 2'h0 == state ? _GEN_6 : _GEN_25; // @[LSU.scala 30:18]
  wire  _GEN_31 = 2'h0 == state ? _GEN_9 : _GEN_21; // @[LSU.scala 30:18]
  assign io_mem_rdata = io_axi_in_rdata; // @[LSU.scala 72:18]
  assign io_axi_out_araddr = io_mem_addr; // @[LSU.scala 73:23]
  assign io_axi_out_arvalid = axi_arvalid; // @[LSU.scala 74:24]
  assign io_axi_out_rready = axi_rready; // @[LSU.scala 75:23]
  assign io_axi_out_awaddr = io_mem_addr; // @[LSU.scala 76:23]
  assign io_axi_out_awvalid = axi_awvalid; // @[LSU.scala 77:24]
  assign io_axi_out_wdata = io_mem_wdata[31:0]; // @[LSU.scala 78:22]
  assign io_axi_out_wstrb = io_mem_wstrb; // @[LSU.scala 79:22]
  assign io_axi_out_wvalid = axi_wvalid; // @[LSU.scala 80:23]
  assign io_axi_out_bready = axi_bready; // @[LSU.scala 81:23]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 19:30]
      axi_arvalid <= 1'h0; // @[LSU.scala 19:30]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      axi_arvalid <= _GEN_5;
    end else if (!(2'h1 == state)) begin // @[LSU.scala 30:18]
      if (2'h2 == state) begin // @[LSU.scala 30:18]
        axi_arvalid <= _GEN_14;
      end
    end
    axi_rready <= reset | _GEN_28; // @[LSU.scala 22:{29,29}]
    if (reset) begin // @[LSU.scala 23:30]
      axi_awvalid <= 1'h0; // @[LSU.scala 23:30]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (!(io_inst_load)) begin // @[LSU.scala 32:31]
        axi_awvalid <= _GEN_1;
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_awready) begin // @[LSU.scala 51:36]
        axi_awvalid <= 1'h0; // @[LSU.scala 52:29]
      end
    end
    if (reset) begin // @[LSU.scala 24:29]
      axi_wvalid <= 1'h0; // @[LSU.scala 24:29]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (!(io_inst_load)) begin // @[LSU.scala 32:31]
        axi_wvalid <= _GEN_2;
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_wready) begin // @[LSU.scala 48:35]
        axi_wvalid <= 1'h0; // @[LSU.scala 49:28]
      end
    end
    axi_bready <= reset | _GEN_31; // @[LSU.scala 25:{29,29}]
    if (reset) begin // @[LSU.scala 28:24]
      state <= 2'h0; // @[LSU.scala 28:24]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (io_inst_load) begin // @[LSU.scala 32:31]
        state <= 2'h2; // @[LSU.scala 33:23]
      end else if (io_inst_store) begin // @[LSU.scala 36:38]
        state <= 2'h1; // @[LSU.scala 37:23]
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_bvalid) begin // @[LSU.scala 44:35]
        state <= 2'h0; // @[LSU.scala 45:23]
      end
    end else if (2'h2 == state) begin // @[LSU.scala 30:18]
      state <= _GEN_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_arvalid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  axi_rready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  axi_awvalid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  axi_wvalid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  axi_bready = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI_ARBITER(
  input         clock,
  input         reset,
  input  [31:0] io_ifu_axi_in_araddr,
  input         io_ifu_axi_in_arvalid,
  input         io_ifu_axi_in_rready,
  output [63:0] io_ifu_axi_out_rdata,
  output        io_ifu_axi_out_rvalid,
  input  [31:0] io_lsu_axi_in_araddr,
  input         io_lsu_axi_in_arvalid,
  input         io_lsu_axi_in_rready,
  input  [31:0] io_lsu_axi_in_awaddr,
  input         io_lsu_axi_in_awvalid,
  input  [31:0] io_lsu_axi_in_wdata,
  input  [7:0]  io_lsu_axi_in_wstrb,
  input         io_lsu_axi_in_wvalid,
  input         io_lsu_axi_in_bready,
  output        io_lsu_axi_out_arready,
  output [63:0] io_lsu_axi_out_rdata,
  output        io_lsu_axi_out_rvalid,
  output        io_lsu_axi_out_awready,
  output        io_lsu_axi_out_wready,
  output        io_lsu_axi_out_bvalid,
  input         io_axi_in_arready,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  input         io_axi_in_awready,
  input         io_axi_in_wready,
  input         io_axi_in_bvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  output [31:0] io_axi_out_awaddr,
  output        io_axi_out_awvalid,
  output [31:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid,
  output        io_axi_out_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[axi_arbiter.scala 18:24]
  wire [1:0] _GEN_0 = io_ifu_axi_in_arvalid ? 2'h1 : state; // @[axi_arbiter.scala 51:46 52:23 18:24]
  wire [31:0] _GEN_1 = io_ifu_axi_in_arvalid ? io_ifu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 51:46 53:28 57:28]
  wire  _GEN_3 = io_ifu_axi_in_arvalid & io_ifu_axi_in_rready; // @[axi_arbiter.scala 51:46 53:28 57:28]
  wire [63:0] _GEN_11 = io_ifu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 51:46 54:32 59:32]
  wire  _GEN_12 = io_ifu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 51:46 54:32 59:32]
  wire [31:0] _GEN_23 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_araddr : _GEN_1; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_24 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_arvalid : io_ifu_axi_in_arvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_25 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_rready : _GEN_3; // @[axi_arbiter.scala 46:46 48:28]
  wire [31:0] _GEN_26 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_27 = io_lsu_axi_in_arvalid & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire [31:0] _GEN_28 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wdata : 32'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire [7:0] _GEN_29 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_30 = io_lsu_axi_in_arvalid & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_31 = io_lsu_axi_in_arvalid & io_lsu_axi_in_bready; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_32 = io_lsu_axi_in_arvalid & io_axi_in_arready; // @[axi_arbiter.scala 46:46 49:32]
  wire [63:0] _GEN_33 = io_lsu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_34 = io_lsu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_35 = io_lsu_axi_in_arvalid & io_axi_in_awready; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_36 = io_lsu_axi_in_arvalid & io_axi_in_wready; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_37 = io_lsu_axi_in_arvalid & io_axi_in_bvalid; // @[axi_arbiter.scala 46:46 49:32]
  wire [63:0] _GEN_39 = io_lsu_axi_in_arvalid ? 64'h0 : _GEN_11; // @[axi_arbiter.scala 46:46 50:32]
  wire  _GEN_40 = io_lsu_axi_in_arvalid ? 1'h0 : _GEN_12; // @[axi_arbiter.scala 46:46 50:32]
  wire [31:0] _GEN_45 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_araddr : _GEN_23; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_46 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_arvalid : _GEN_24; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_47 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_rready : _GEN_25; // @[axi_arbiter.scala 41:40 43:28]
  wire [31:0] _GEN_48 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awaddr : _GEN_26; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_49 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awvalid : _GEN_27; // @[axi_arbiter.scala 41:40 43:28]
  wire [31:0] _GEN_50 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wdata : _GEN_28; // @[axi_arbiter.scala 41:40 43:28]
  wire [7:0] _GEN_51 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wstrb : _GEN_29; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_52 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wvalid : _GEN_30; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_53 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_bready : _GEN_31; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_54 = io_lsu_axi_in_awvalid ? io_axi_in_arready : _GEN_32; // @[axi_arbiter.scala 41:40 44:32]
  wire [63:0] _GEN_55 = io_lsu_axi_in_awvalid ? io_axi_in_rdata : _GEN_33; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_56 = io_lsu_axi_in_awvalid ? io_axi_in_rvalid : _GEN_34; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_57 = io_lsu_axi_in_awvalid ? io_axi_in_awready : _GEN_35; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_58 = io_lsu_axi_in_awvalid ? io_axi_in_wready : _GEN_36; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_59 = io_lsu_axi_in_awvalid ? io_axi_in_bvalid : _GEN_37; // @[axi_arbiter.scala 41:40 44:32]
  wire [63:0] _GEN_61 = io_lsu_axi_in_awvalid ? 64'h0 : _GEN_39; // @[axi_arbiter.scala 41:40 45:32]
  wire  _GEN_62 = io_lsu_axi_in_awvalid ? 1'h0 : _GEN_40; // @[axi_arbiter.scala 41:40 45:32]
  wire [1:0] _GEN_67 = io_lsu_axi_out_rvalid & io_lsu_axi_in_rready ? 2'h0 : state; // @[axi_arbiter.scala 74:64 75:23 18:24]
  wire [1:0] _GEN_68 = io_lsu_axi_out_bvalid & io_lsu_axi_in_bready ? 2'h0 : state; // @[axi_arbiter.scala 82:64 83:23 18:24]
  wire [31:0] _GEN_69 = state == 2'h3 ? io_lsu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_70 = state == 2'h3 & io_lsu_axi_in_arvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_71 = state == 2'h3 & io_lsu_axi_in_rready; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [31:0] _GEN_72 = state == 2'h3 ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_73 = state == 2'h3 & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [31:0] _GEN_74 = state == 2'h3 ? io_lsu_axi_in_wdata : 32'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [7:0] _GEN_75 = state == 2'h3 ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_76 = state == 2'h3 & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_77 = state == 2'h3 & io_lsu_axi_in_bready; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_78 = state == 2'h3 & io_axi_in_arready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire [63:0] _GEN_79 = state == 2'h3 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_80 = state == 2'h3 & io_axi_in_rvalid; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_81 = state == 2'h3 & io_axi_in_awready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_82 = state == 2'h3 & io_axi_in_wready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_83 = state == 2'h3 & io_axi_in_bvalid; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire [1:0] _GEN_90 = state == 2'h3 ? _GEN_68 : state; // @[axi_arbiter.scala 18:24 78:39]
  wire [31:0] _GEN_91 = state == 2'h2 ? io_lsu_axi_in_araddr : _GEN_69; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_92 = state == 2'h2 ? io_lsu_axi_in_arvalid : _GEN_70; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_93 = state == 2'h2 ? io_lsu_axi_in_rready : _GEN_71; // @[axi_arbiter.scala 70:39 71:24]
  wire [31:0] _GEN_94 = state == 2'h2 ? io_lsu_axi_in_awaddr : _GEN_72; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_95 = state == 2'h2 ? io_lsu_axi_in_awvalid : _GEN_73; // @[axi_arbiter.scala 70:39 71:24]
  wire [31:0] _GEN_96 = state == 2'h2 ? io_lsu_axi_in_wdata : _GEN_74; // @[axi_arbiter.scala 70:39 71:24]
  wire [7:0] _GEN_97 = state == 2'h2 ? io_lsu_axi_in_wstrb : _GEN_75; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_98 = state == 2'h2 ? io_lsu_axi_in_wvalid : _GEN_76; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_99 = state == 2'h2 ? io_lsu_axi_in_bready : _GEN_77; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_100 = state == 2'h2 ? io_axi_in_arready : _GEN_78; // @[axi_arbiter.scala 70:39 72:28]
  wire [63:0] _GEN_101 = state == 2'h2 ? io_axi_in_rdata : _GEN_79; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_102 = state == 2'h2 ? io_axi_in_rvalid : _GEN_80; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_103 = state == 2'h2 ? io_axi_in_awready : _GEN_81; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_104 = state == 2'h2 ? io_axi_in_wready : _GEN_82; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_105 = state == 2'h2 ? io_axi_in_bvalid : _GEN_83; // @[axi_arbiter.scala 70:39 72:28]
  wire [31:0] _GEN_113 = state == 2'h1 ? io_ifu_axi_in_araddr : _GEN_91; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_114 = state == 2'h1 ? io_ifu_axi_in_arvalid : _GEN_92; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_115 = state == 2'h1 ? io_ifu_axi_in_rready : _GEN_93; // @[axi_arbiter.scala 62:39 63:24]
  wire [31:0] _GEN_116 = state == 2'h1 ? 32'h0 : _GEN_94; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_117 = state == 2'h1 ? 1'h0 : _GEN_95; // @[axi_arbiter.scala 62:39 63:24]
  wire [31:0] _GEN_118 = state == 2'h1 ? 32'h0 : _GEN_96; // @[axi_arbiter.scala 62:39 63:24]
  wire [7:0] _GEN_119 = state == 2'h1 ? 8'h0 : _GEN_97; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_120 = state == 2'h1 ? 1'h0 : _GEN_98; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_121 = state == 2'h1 ? 1'h0 : _GEN_99; // @[axi_arbiter.scala 62:39 63:24]
  wire [63:0] _GEN_123 = state == 2'h1 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 62:39 64:28]
  wire  _GEN_124 = state == 2'h1 & io_axi_in_rvalid; // @[axi_arbiter.scala 62:39 64:28]
  wire  _GEN_128 = state == 2'h1 ? 1'h0 : _GEN_100; // @[axi_arbiter.scala 62:39 65:28]
  wire [63:0] _GEN_129 = state == 2'h1 ? 64'h0 : _GEN_101; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_130 = state == 2'h1 ? 1'h0 : _GEN_102; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_131 = state == 2'h1 ? 1'h0 : _GEN_103; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_132 = state == 2'h1 ? 1'h0 : _GEN_104; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_133 = state == 2'h1 ? 1'h0 : _GEN_105; // @[axi_arbiter.scala 62:39 65:28]
  assign io_ifu_axi_out_rdata = state == 2'h0 ? _GEN_61 : _GEN_123; // @[axi_arbiter.scala 40:27]
  assign io_ifu_axi_out_rvalid = state == 2'h0 ? _GEN_62 : _GEN_124; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_arready = state == 2'h0 ? _GEN_54 : _GEN_128; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_rdata = state == 2'h0 ? _GEN_55 : _GEN_129; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_rvalid = state == 2'h0 ? _GEN_56 : _GEN_130; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_awready = state == 2'h0 ? _GEN_57 : _GEN_131; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_wready = state == 2'h0 ? _GEN_58 : _GEN_132; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_bvalid = state == 2'h0 ? _GEN_59 : _GEN_133; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_araddr = state == 2'h0 ? _GEN_45 : _GEN_113; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_arvalid = state == 2'h0 ? _GEN_46 : _GEN_114; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_rready = state == 2'h0 ? _GEN_47 : _GEN_115; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_awaddr = state == 2'h0 ? _GEN_48 : _GEN_116; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_awvalid = state == 2'h0 ? _GEN_49 : _GEN_117; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wdata = state == 2'h0 ? _GEN_50 : _GEN_118; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wstrb = state == 2'h0 ? _GEN_51 : _GEN_119; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wvalid = state == 2'h0 ? _GEN_52 : _GEN_120; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_bready = state == 2'h0 ? _GEN_53 : _GEN_121; // @[axi_arbiter.scala 40:27]
  always @(posedge clock) begin
    if (reset) begin // @[axi_arbiter.scala 18:24]
      state <= 2'h0; // @[axi_arbiter.scala 18:24]
    end else if (state == 2'h0) begin // @[axi_arbiter.scala 40:27]
      if (io_lsu_axi_in_awvalid) begin // @[axi_arbiter.scala 41:40]
        state <= 2'h3; // @[axi_arbiter.scala 42:23]
      end else if (io_lsu_axi_in_arvalid) begin // @[axi_arbiter.scala 46:46]
        state <= 2'h2; // @[axi_arbiter.scala 47:23]
      end else begin
        state <= _GEN_0;
      end
    end else if (state == 2'h1) begin // @[axi_arbiter.scala 62:39]
      if (io_ifu_axi_out_rvalid & io_ifu_axi_in_rready) begin // @[axi_arbiter.scala 66:64]
        state <= 2'h0; // @[axi_arbiter.scala 67:23]
      end
    end else if (state == 2'h2) begin // @[axi_arbiter.scala 70:39]
      state <= _GEN_67;
    end else begin
      state <= _GEN_90;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU_AXI(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_pc_valid,
  output        io_inst_valid,
  output [31:0] io_inst,
  output [31:0] io_inst_reg,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  inst_ready; // @[IFU_AXI.scala 19:29]
  wire  _GEN_0 = io_axi_in_rvalid & inst_ready ? 1'h0 : 1'h1; // @[IFU_AXI.scala 20:41 21:20 23:20]
  reg [31:0] inst_reg; // @[IFU_AXI.scala 25:27]
  assign io_inst_valid = io_axi_in_rvalid; // @[IFU_AXI.scala 43:19]
  assign io_inst = io_axi_in_rdata[31:0]; // @[IFU_AXI.scala 41:31]
  assign io_inst_reg = inst_reg; // @[IFU_AXI.scala 42:17]
  assign io_axi_out_araddr = io_pc[31:0]; // @[IFU_AXI.scala 31:31]
  assign io_axi_out_arvalid = io_pc_valid; // @[IFU_AXI.scala 32:24]
  assign io_axi_out_rready = inst_ready; // @[IFU_AXI.scala 33:23]
  always @(posedge clock) begin
    inst_ready <= reset | _GEN_0; // @[IFU_AXI.scala 19:{29,29}]
    if (reset) begin // @[IFU_AXI.scala 25:27]
      inst_reg <= 32'h0; // @[IFU_AXI.scala 25:27]
    end else if (io_axi_in_rvalid) begin // @[IFU_AXI.scala 26:27]
      inst_reg <= io_axi_in_rdata[31:0]; // @[IFU_AXI.scala 27:18]
    end else if (io_pc_valid) begin // @[IFU_AXI.scala 28:28]
      inst_reg <= 32'h0; // @[IFU_AXI.scala 29:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst_ready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  inst_reg = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module I_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_ifu_araddr,
  input         io_from_ifu_arvalid,
  input         io_from_ifu_rready,
  output [63:0] io_to_ifu_rdata,
  output        io_to_ifu_rvalid,
  output [31:0] io_to_axi_araddr,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [63:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_0_0; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_1; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_2; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_3; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_4; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_5; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_6; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_7; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_8; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_9; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_10; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_11; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_12; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_13; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_14; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_15; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_16; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_17; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_18; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_19; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_20; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_21; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_22; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_23; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_24; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_25; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_26; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_27; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_28; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_29; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_30; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_31; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_32; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_33; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_34; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_35; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_36; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_37; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_38; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_39; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_40; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_41; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_42; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_43; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_44; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_45; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_46; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_47; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_48; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_49; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_50; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_51; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_52; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_53; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_54; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_55; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_56; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_57; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_58; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_59; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_60; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_61; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_62; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_63; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_64; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_65; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_66; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_67; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_68; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_69; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_70; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_71; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_72; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_73; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_74; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_75; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_76; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_77; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_78; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_79; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_80; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_81; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_82; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_83; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_84; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_85; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_86; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_87; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_88; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_89; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_90; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_91; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_92; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_93; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_94; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_95; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_96; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_97; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_98; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_99; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_100; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_101; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_102; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_103; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_104; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_105; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_106; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_107; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_108; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_109; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_110; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_111; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_112; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_113; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_114; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_115; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_116; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_117; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_118; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_119; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_120; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_121; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_122; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_123; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_124; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_125; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_126; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_127; // @[i_cache.scala 17:24]
  reg [63:0] ram_1_0; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_1; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_2; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_3; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_4; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_5; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_6; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_7; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_8; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_9; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_10; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_11; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_12; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_13; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_14; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_15; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_16; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_17; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_18; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_19; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_20; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_21; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_22; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_23; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_24; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_25; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_26; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_27; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_28; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_29; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_30; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_31; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_32; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_33; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_34; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_35; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_36; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_37; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_38; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_39; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_40; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_41; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_42; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_43; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_44; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_45; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_46; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_47; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_48; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_49; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_50; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_51; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_52; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_53; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_54; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_55; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_56; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_57; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_58; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_59; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_60; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_61; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_62; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_63; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_64; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_65; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_66; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_67; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_68; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_69; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_70; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_71; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_72; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_73; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_74; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_75; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_76; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_77; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_78; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_79; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_80; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_81; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_82; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_83; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_84; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_85; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_86; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_87; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_88; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_89; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_90; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_91; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_92; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_93; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_94; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_95; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_96; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_97; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_98; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_99; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_100; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_101; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_102; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_103; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_104; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_105; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_106; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_107; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_108; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_109; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_110; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_111; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_112; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_113; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_114; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_115; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_116; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_117; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_118; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_119; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_120; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_121; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_122; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_123; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_124; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_125; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_126; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_127; // @[i_cache.scala 18:24]
  reg [31:0] tag_0_0; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_1; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_2; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_3; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_4; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_5; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_6; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_7; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_8; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_9; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_10; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_11; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_12; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_13; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_14; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_15; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_16; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_17; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_18; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_19; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_20; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_21; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_22; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_23; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_24; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_25; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_26; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_27; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_28; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_29; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_30; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_31; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_32; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_33; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_34; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_35; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_36; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_37; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_38; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_39; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_40; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_41; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_42; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_43; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_44; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_45; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_46; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_47; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_48; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_49; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_50; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_51; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_52; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_53; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_54; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_55; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_56; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_57; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_58; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_59; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_60; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_61; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_62; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_63; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_64; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_65; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_66; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_67; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_68; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_69; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_70; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_71; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_72; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_73; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_74; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_75; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_76; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_77; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_78; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_79; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_80; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_81; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_82; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_83; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_84; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_85; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_86; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_87; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_88; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_89; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_90; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_91; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_92; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_93; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_94; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_95; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_96; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_97; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_98; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_99; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_100; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_101; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_102; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_103; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_104; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_105; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_106; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_107; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_108; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_109; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_110; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_111; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_112; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_113; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_114; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_115; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_116; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_117; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_118; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_119; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_120; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_121; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_122; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_123; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_124; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_125; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_126; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_127; // @[i_cache.scala 19:24]
  reg [31:0] tag_1_0; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_1; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_2; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_3; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_4; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_5; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_6; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_7; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_8; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_9; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_10; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_11; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_12; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_13; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_14; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_15; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_16; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_17; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_18; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_19; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_20; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_21; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_22; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_23; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_24; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_25; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_26; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_27; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_28; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_29; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_30; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_31; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_32; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_33; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_34; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_35; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_36; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_37; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_38; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_39; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_40; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_41; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_42; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_43; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_44; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_45; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_46; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_47; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_48; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_49; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_50; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_51; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_52; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_53; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_54; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_55; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_56; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_57; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_58; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_59; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_60; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_61; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_62; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_63; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_64; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_65; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_66; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_67; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_68; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_69; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_70; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_71; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_72; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_73; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_74; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_75; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_76; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_77; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_78; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_79; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_80; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_81; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_82; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_83; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_84; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_85; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_86; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_87; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_88; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_89; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_90; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_91; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_92; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_93; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_94; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_95; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_96; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_97; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_98; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_99; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_100; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_101; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_102; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_103; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_104; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_105; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_106; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_107; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_108; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_109; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_110; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_111; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_112; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_113; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_114; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_115; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_116; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_117; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_118; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_119; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_120; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_121; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_122; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_123; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_124; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_125; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_126; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_127; // @[i_cache.scala 20:24]
  reg  valid_0_0; // @[i_cache.scala 21:26]
  reg  valid_0_1; // @[i_cache.scala 21:26]
  reg  valid_0_2; // @[i_cache.scala 21:26]
  reg  valid_0_3; // @[i_cache.scala 21:26]
  reg  valid_0_4; // @[i_cache.scala 21:26]
  reg  valid_0_5; // @[i_cache.scala 21:26]
  reg  valid_0_6; // @[i_cache.scala 21:26]
  reg  valid_0_7; // @[i_cache.scala 21:26]
  reg  valid_0_8; // @[i_cache.scala 21:26]
  reg  valid_0_9; // @[i_cache.scala 21:26]
  reg  valid_0_10; // @[i_cache.scala 21:26]
  reg  valid_0_11; // @[i_cache.scala 21:26]
  reg  valid_0_12; // @[i_cache.scala 21:26]
  reg  valid_0_13; // @[i_cache.scala 21:26]
  reg  valid_0_14; // @[i_cache.scala 21:26]
  reg  valid_0_15; // @[i_cache.scala 21:26]
  reg  valid_0_16; // @[i_cache.scala 21:26]
  reg  valid_0_17; // @[i_cache.scala 21:26]
  reg  valid_0_18; // @[i_cache.scala 21:26]
  reg  valid_0_19; // @[i_cache.scala 21:26]
  reg  valid_0_20; // @[i_cache.scala 21:26]
  reg  valid_0_21; // @[i_cache.scala 21:26]
  reg  valid_0_22; // @[i_cache.scala 21:26]
  reg  valid_0_23; // @[i_cache.scala 21:26]
  reg  valid_0_24; // @[i_cache.scala 21:26]
  reg  valid_0_25; // @[i_cache.scala 21:26]
  reg  valid_0_26; // @[i_cache.scala 21:26]
  reg  valid_0_27; // @[i_cache.scala 21:26]
  reg  valid_0_28; // @[i_cache.scala 21:26]
  reg  valid_0_29; // @[i_cache.scala 21:26]
  reg  valid_0_30; // @[i_cache.scala 21:26]
  reg  valid_0_31; // @[i_cache.scala 21:26]
  reg  valid_0_32; // @[i_cache.scala 21:26]
  reg  valid_0_33; // @[i_cache.scala 21:26]
  reg  valid_0_34; // @[i_cache.scala 21:26]
  reg  valid_0_35; // @[i_cache.scala 21:26]
  reg  valid_0_36; // @[i_cache.scala 21:26]
  reg  valid_0_37; // @[i_cache.scala 21:26]
  reg  valid_0_38; // @[i_cache.scala 21:26]
  reg  valid_0_39; // @[i_cache.scala 21:26]
  reg  valid_0_40; // @[i_cache.scala 21:26]
  reg  valid_0_41; // @[i_cache.scala 21:26]
  reg  valid_0_42; // @[i_cache.scala 21:26]
  reg  valid_0_43; // @[i_cache.scala 21:26]
  reg  valid_0_44; // @[i_cache.scala 21:26]
  reg  valid_0_45; // @[i_cache.scala 21:26]
  reg  valid_0_46; // @[i_cache.scala 21:26]
  reg  valid_0_47; // @[i_cache.scala 21:26]
  reg  valid_0_48; // @[i_cache.scala 21:26]
  reg  valid_0_49; // @[i_cache.scala 21:26]
  reg  valid_0_50; // @[i_cache.scala 21:26]
  reg  valid_0_51; // @[i_cache.scala 21:26]
  reg  valid_0_52; // @[i_cache.scala 21:26]
  reg  valid_0_53; // @[i_cache.scala 21:26]
  reg  valid_0_54; // @[i_cache.scala 21:26]
  reg  valid_0_55; // @[i_cache.scala 21:26]
  reg  valid_0_56; // @[i_cache.scala 21:26]
  reg  valid_0_57; // @[i_cache.scala 21:26]
  reg  valid_0_58; // @[i_cache.scala 21:26]
  reg  valid_0_59; // @[i_cache.scala 21:26]
  reg  valid_0_60; // @[i_cache.scala 21:26]
  reg  valid_0_61; // @[i_cache.scala 21:26]
  reg  valid_0_62; // @[i_cache.scala 21:26]
  reg  valid_0_63; // @[i_cache.scala 21:26]
  reg  valid_0_64; // @[i_cache.scala 21:26]
  reg  valid_0_65; // @[i_cache.scala 21:26]
  reg  valid_0_66; // @[i_cache.scala 21:26]
  reg  valid_0_67; // @[i_cache.scala 21:26]
  reg  valid_0_68; // @[i_cache.scala 21:26]
  reg  valid_0_69; // @[i_cache.scala 21:26]
  reg  valid_0_70; // @[i_cache.scala 21:26]
  reg  valid_0_71; // @[i_cache.scala 21:26]
  reg  valid_0_72; // @[i_cache.scala 21:26]
  reg  valid_0_73; // @[i_cache.scala 21:26]
  reg  valid_0_74; // @[i_cache.scala 21:26]
  reg  valid_0_75; // @[i_cache.scala 21:26]
  reg  valid_0_76; // @[i_cache.scala 21:26]
  reg  valid_0_77; // @[i_cache.scala 21:26]
  reg  valid_0_78; // @[i_cache.scala 21:26]
  reg  valid_0_79; // @[i_cache.scala 21:26]
  reg  valid_0_80; // @[i_cache.scala 21:26]
  reg  valid_0_81; // @[i_cache.scala 21:26]
  reg  valid_0_82; // @[i_cache.scala 21:26]
  reg  valid_0_83; // @[i_cache.scala 21:26]
  reg  valid_0_84; // @[i_cache.scala 21:26]
  reg  valid_0_85; // @[i_cache.scala 21:26]
  reg  valid_0_86; // @[i_cache.scala 21:26]
  reg  valid_0_87; // @[i_cache.scala 21:26]
  reg  valid_0_88; // @[i_cache.scala 21:26]
  reg  valid_0_89; // @[i_cache.scala 21:26]
  reg  valid_0_90; // @[i_cache.scala 21:26]
  reg  valid_0_91; // @[i_cache.scala 21:26]
  reg  valid_0_92; // @[i_cache.scala 21:26]
  reg  valid_0_93; // @[i_cache.scala 21:26]
  reg  valid_0_94; // @[i_cache.scala 21:26]
  reg  valid_0_95; // @[i_cache.scala 21:26]
  reg  valid_0_96; // @[i_cache.scala 21:26]
  reg  valid_0_97; // @[i_cache.scala 21:26]
  reg  valid_0_98; // @[i_cache.scala 21:26]
  reg  valid_0_99; // @[i_cache.scala 21:26]
  reg  valid_0_100; // @[i_cache.scala 21:26]
  reg  valid_0_101; // @[i_cache.scala 21:26]
  reg  valid_0_102; // @[i_cache.scala 21:26]
  reg  valid_0_103; // @[i_cache.scala 21:26]
  reg  valid_0_104; // @[i_cache.scala 21:26]
  reg  valid_0_105; // @[i_cache.scala 21:26]
  reg  valid_0_106; // @[i_cache.scala 21:26]
  reg  valid_0_107; // @[i_cache.scala 21:26]
  reg  valid_0_108; // @[i_cache.scala 21:26]
  reg  valid_0_109; // @[i_cache.scala 21:26]
  reg  valid_0_110; // @[i_cache.scala 21:26]
  reg  valid_0_111; // @[i_cache.scala 21:26]
  reg  valid_0_112; // @[i_cache.scala 21:26]
  reg  valid_0_113; // @[i_cache.scala 21:26]
  reg  valid_0_114; // @[i_cache.scala 21:26]
  reg  valid_0_115; // @[i_cache.scala 21:26]
  reg  valid_0_116; // @[i_cache.scala 21:26]
  reg  valid_0_117; // @[i_cache.scala 21:26]
  reg  valid_0_118; // @[i_cache.scala 21:26]
  reg  valid_0_119; // @[i_cache.scala 21:26]
  reg  valid_0_120; // @[i_cache.scala 21:26]
  reg  valid_0_121; // @[i_cache.scala 21:26]
  reg  valid_0_122; // @[i_cache.scala 21:26]
  reg  valid_0_123; // @[i_cache.scala 21:26]
  reg  valid_0_124; // @[i_cache.scala 21:26]
  reg  valid_0_125; // @[i_cache.scala 21:26]
  reg  valid_0_126; // @[i_cache.scala 21:26]
  reg  valid_0_127; // @[i_cache.scala 21:26]
  reg  valid_1_0; // @[i_cache.scala 22:26]
  reg  valid_1_1; // @[i_cache.scala 22:26]
  reg  valid_1_2; // @[i_cache.scala 22:26]
  reg  valid_1_3; // @[i_cache.scala 22:26]
  reg  valid_1_4; // @[i_cache.scala 22:26]
  reg  valid_1_5; // @[i_cache.scala 22:26]
  reg  valid_1_6; // @[i_cache.scala 22:26]
  reg  valid_1_7; // @[i_cache.scala 22:26]
  reg  valid_1_8; // @[i_cache.scala 22:26]
  reg  valid_1_9; // @[i_cache.scala 22:26]
  reg  valid_1_10; // @[i_cache.scala 22:26]
  reg  valid_1_11; // @[i_cache.scala 22:26]
  reg  valid_1_12; // @[i_cache.scala 22:26]
  reg  valid_1_13; // @[i_cache.scala 22:26]
  reg  valid_1_14; // @[i_cache.scala 22:26]
  reg  valid_1_15; // @[i_cache.scala 22:26]
  reg  valid_1_16; // @[i_cache.scala 22:26]
  reg  valid_1_17; // @[i_cache.scala 22:26]
  reg  valid_1_18; // @[i_cache.scala 22:26]
  reg  valid_1_19; // @[i_cache.scala 22:26]
  reg  valid_1_20; // @[i_cache.scala 22:26]
  reg  valid_1_21; // @[i_cache.scala 22:26]
  reg  valid_1_22; // @[i_cache.scala 22:26]
  reg  valid_1_23; // @[i_cache.scala 22:26]
  reg  valid_1_24; // @[i_cache.scala 22:26]
  reg  valid_1_25; // @[i_cache.scala 22:26]
  reg  valid_1_26; // @[i_cache.scala 22:26]
  reg  valid_1_27; // @[i_cache.scala 22:26]
  reg  valid_1_28; // @[i_cache.scala 22:26]
  reg  valid_1_29; // @[i_cache.scala 22:26]
  reg  valid_1_30; // @[i_cache.scala 22:26]
  reg  valid_1_31; // @[i_cache.scala 22:26]
  reg  valid_1_32; // @[i_cache.scala 22:26]
  reg  valid_1_33; // @[i_cache.scala 22:26]
  reg  valid_1_34; // @[i_cache.scala 22:26]
  reg  valid_1_35; // @[i_cache.scala 22:26]
  reg  valid_1_36; // @[i_cache.scala 22:26]
  reg  valid_1_37; // @[i_cache.scala 22:26]
  reg  valid_1_38; // @[i_cache.scala 22:26]
  reg  valid_1_39; // @[i_cache.scala 22:26]
  reg  valid_1_40; // @[i_cache.scala 22:26]
  reg  valid_1_41; // @[i_cache.scala 22:26]
  reg  valid_1_42; // @[i_cache.scala 22:26]
  reg  valid_1_43; // @[i_cache.scala 22:26]
  reg  valid_1_44; // @[i_cache.scala 22:26]
  reg  valid_1_45; // @[i_cache.scala 22:26]
  reg  valid_1_46; // @[i_cache.scala 22:26]
  reg  valid_1_47; // @[i_cache.scala 22:26]
  reg  valid_1_48; // @[i_cache.scala 22:26]
  reg  valid_1_49; // @[i_cache.scala 22:26]
  reg  valid_1_50; // @[i_cache.scala 22:26]
  reg  valid_1_51; // @[i_cache.scala 22:26]
  reg  valid_1_52; // @[i_cache.scala 22:26]
  reg  valid_1_53; // @[i_cache.scala 22:26]
  reg  valid_1_54; // @[i_cache.scala 22:26]
  reg  valid_1_55; // @[i_cache.scala 22:26]
  reg  valid_1_56; // @[i_cache.scala 22:26]
  reg  valid_1_57; // @[i_cache.scala 22:26]
  reg  valid_1_58; // @[i_cache.scala 22:26]
  reg  valid_1_59; // @[i_cache.scala 22:26]
  reg  valid_1_60; // @[i_cache.scala 22:26]
  reg  valid_1_61; // @[i_cache.scala 22:26]
  reg  valid_1_62; // @[i_cache.scala 22:26]
  reg  valid_1_63; // @[i_cache.scala 22:26]
  reg  valid_1_64; // @[i_cache.scala 22:26]
  reg  valid_1_65; // @[i_cache.scala 22:26]
  reg  valid_1_66; // @[i_cache.scala 22:26]
  reg  valid_1_67; // @[i_cache.scala 22:26]
  reg  valid_1_68; // @[i_cache.scala 22:26]
  reg  valid_1_69; // @[i_cache.scala 22:26]
  reg  valid_1_70; // @[i_cache.scala 22:26]
  reg  valid_1_71; // @[i_cache.scala 22:26]
  reg  valid_1_72; // @[i_cache.scala 22:26]
  reg  valid_1_73; // @[i_cache.scala 22:26]
  reg  valid_1_74; // @[i_cache.scala 22:26]
  reg  valid_1_75; // @[i_cache.scala 22:26]
  reg  valid_1_76; // @[i_cache.scala 22:26]
  reg  valid_1_77; // @[i_cache.scala 22:26]
  reg  valid_1_78; // @[i_cache.scala 22:26]
  reg  valid_1_79; // @[i_cache.scala 22:26]
  reg  valid_1_80; // @[i_cache.scala 22:26]
  reg  valid_1_81; // @[i_cache.scala 22:26]
  reg  valid_1_82; // @[i_cache.scala 22:26]
  reg  valid_1_83; // @[i_cache.scala 22:26]
  reg  valid_1_84; // @[i_cache.scala 22:26]
  reg  valid_1_85; // @[i_cache.scala 22:26]
  reg  valid_1_86; // @[i_cache.scala 22:26]
  reg  valid_1_87; // @[i_cache.scala 22:26]
  reg  valid_1_88; // @[i_cache.scala 22:26]
  reg  valid_1_89; // @[i_cache.scala 22:26]
  reg  valid_1_90; // @[i_cache.scala 22:26]
  reg  valid_1_91; // @[i_cache.scala 22:26]
  reg  valid_1_92; // @[i_cache.scala 22:26]
  reg  valid_1_93; // @[i_cache.scala 22:26]
  reg  valid_1_94; // @[i_cache.scala 22:26]
  reg  valid_1_95; // @[i_cache.scala 22:26]
  reg  valid_1_96; // @[i_cache.scala 22:26]
  reg  valid_1_97; // @[i_cache.scala 22:26]
  reg  valid_1_98; // @[i_cache.scala 22:26]
  reg  valid_1_99; // @[i_cache.scala 22:26]
  reg  valid_1_100; // @[i_cache.scala 22:26]
  reg  valid_1_101; // @[i_cache.scala 22:26]
  reg  valid_1_102; // @[i_cache.scala 22:26]
  reg  valid_1_103; // @[i_cache.scala 22:26]
  reg  valid_1_104; // @[i_cache.scala 22:26]
  reg  valid_1_105; // @[i_cache.scala 22:26]
  reg  valid_1_106; // @[i_cache.scala 22:26]
  reg  valid_1_107; // @[i_cache.scala 22:26]
  reg  valid_1_108; // @[i_cache.scala 22:26]
  reg  valid_1_109; // @[i_cache.scala 22:26]
  reg  valid_1_110; // @[i_cache.scala 22:26]
  reg  valid_1_111; // @[i_cache.scala 22:26]
  reg  valid_1_112; // @[i_cache.scala 22:26]
  reg  valid_1_113; // @[i_cache.scala 22:26]
  reg  valid_1_114; // @[i_cache.scala 22:26]
  reg  valid_1_115; // @[i_cache.scala 22:26]
  reg  valid_1_116; // @[i_cache.scala 22:26]
  reg  valid_1_117; // @[i_cache.scala 22:26]
  reg  valid_1_118; // @[i_cache.scala 22:26]
  reg  valid_1_119; // @[i_cache.scala 22:26]
  reg  valid_1_120; // @[i_cache.scala 22:26]
  reg  valid_1_121; // @[i_cache.scala 22:26]
  reg  valid_1_122; // @[i_cache.scala 22:26]
  reg  valid_1_123; // @[i_cache.scala 22:26]
  reg  valid_1_124; // @[i_cache.scala 22:26]
  reg  valid_1_125; // @[i_cache.scala 22:26]
  reg  valid_1_126; // @[i_cache.scala 22:26]
  reg  valid_1_127; // @[i_cache.scala 22:26]
  reg  way0_hit; // @[i_cache.scala 23:27]
  reg  way1_hit; // @[i_cache.scala 24:27]
  reg [1:0] unuse_way; // @[i_cache.scala 26:28]
  reg [63:0] receive_data; // @[i_cache.scala 27:31]
  reg  quene; // @[i_cache.scala 28:24]
  wire [6:0] index = io_from_ifu_araddr[6:0]; // @[i_cache.scala 31:35]
  wire [24:0] tag = io_from_ifu_araddr[31:7]; // @[i_cache.scala 32:33]
  wire [31:0] _GEN_1 = 7'h1 == index ? tag_0_1 : tag_0_0; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_2 = 7'h2 == index ? tag_0_2 : _GEN_1; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_3 = 7'h3 == index ? tag_0_3 : _GEN_2; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_4 = 7'h4 == index ? tag_0_4 : _GEN_3; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_5 = 7'h5 == index ? tag_0_5 : _GEN_4; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_6 = 7'h6 == index ? tag_0_6 : _GEN_5; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_7 = 7'h7 == index ? tag_0_7 : _GEN_6; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_8 = 7'h8 == index ? tag_0_8 : _GEN_7; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_9 = 7'h9 == index ? tag_0_9 : _GEN_8; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_10 = 7'ha == index ? tag_0_10 : _GEN_9; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_11 = 7'hb == index ? tag_0_11 : _GEN_10; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_12 = 7'hc == index ? tag_0_12 : _GEN_11; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_13 = 7'hd == index ? tag_0_13 : _GEN_12; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_14 = 7'he == index ? tag_0_14 : _GEN_13; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_15 = 7'hf == index ? tag_0_15 : _GEN_14; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_16 = 7'h10 == index ? tag_0_16 : _GEN_15; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_17 = 7'h11 == index ? tag_0_17 : _GEN_16; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_18 = 7'h12 == index ? tag_0_18 : _GEN_17; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_19 = 7'h13 == index ? tag_0_19 : _GEN_18; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_20 = 7'h14 == index ? tag_0_20 : _GEN_19; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_21 = 7'h15 == index ? tag_0_21 : _GEN_20; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_22 = 7'h16 == index ? tag_0_22 : _GEN_21; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_23 = 7'h17 == index ? tag_0_23 : _GEN_22; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_24 = 7'h18 == index ? tag_0_24 : _GEN_23; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_25 = 7'h19 == index ? tag_0_25 : _GEN_24; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_26 = 7'h1a == index ? tag_0_26 : _GEN_25; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_27 = 7'h1b == index ? tag_0_27 : _GEN_26; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_28 = 7'h1c == index ? tag_0_28 : _GEN_27; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_29 = 7'h1d == index ? tag_0_29 : _GEN_28; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_30 = 7'h1e == index ? tag_0_30 : _GEN_29; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_31 = 7'h1f == index ? tag_0_31 : _GEN_30; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_32 = 7'h20 == index ? tag_0_32 : _GEN_31; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_33 = 7'h21 == index ? tag_0_33 : _GEN_32; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_34 = 7'h22 == index ? tag_0_34 : _GEN_33; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_35 = 7'h23 == index ? tag_0_35 : _GEN_34; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_36 = 7'h24 == index ? tag_0_36 : _GEN_35; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_37 = 7'h25 == index ? tag_0_37 : _GEN_36; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_38 = 7'h26 == index ? tag_0_38 : _GEN_37; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_39 = 7'h27 == index ? tag_0_39 : _GEN_38; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_40 = 7'h28 == index ? tag_0_40 : _GEN_39; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_41 = 7'h29 == index ? tag_0_41 : _GEN_40; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_42 = 7'h2a == index ? tag_0_42 : _GEN_41; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_43 = 7'h2b == index ? tag_0_43 : _GEN_42; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_44 = 7'h2c == index ? tag_0_44 : _GEN_43; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_45 = 7'h2d == index ? tag_0_45 : _GEN_44; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_46 = 7'h2e == index ? tag_0_46 : _GEN_45; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_47 = 7'h2f == index ? tag_0_47 : _GEN_46; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_48 = 7'h30 == index ? tag_0_48 : _GEN_47; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_49 = 7'h31 == index ? tag_0_49 : _GEN_48; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_50 = 7'h32 == index ? tag_0_50 : _GEN_49; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_51 = 7'h33 == index ? tag_0_51 : _GEN_50; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_52 = 7'h34 == index ? tag_0_52 : _GEN_51; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_53 = 7'h35 == index ? tag_0_53 : _GEN_52; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_54 = 7'h36 == index ? tag_0_54 : _GEN_53; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_55 = 7'h37 == index ? tag_0_55 : _GEN_54; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_56 = 7'h38 == index ? tag_0_56 : _GEN_55; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_57 = 7'h39 == index ? tag_0_57 : _GEN_56; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_58 = 7'h3a == index ? tag_0_58 : _GEN_57; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_59 = 7'h3b == index ? tag_0_59 : _GEN_58; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_60 = 7'h3c == index ? tag_0_60 : _GEN_59; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_61 = 7'h3d == index ? tag_0_61 : _GEN_60; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_62 = 7'h3e == index ? tag_0_62 : _GEN_61; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_63 = 7'h3f == index ? tag_0_63 : _GEN_62; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_64 = 7'h40 == index ? tag_0_64 : _GEN_63; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_65 = 7'h41 == index ? tag_0_65 : _GEN_64; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_66 = 7'h42 == index ? tag_0_66 : _GEN_65; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_67 = 7'h43 == index ? tag_0_67 : _GEN_66; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_68 = 7'h44 == index ? tag_0_68 : _GEN_67; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_69 = 7'h45 == index ? tag_0_69 : _GEN_68; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_70 = 7'h46 == index ? tag_0_70 : _GEN_69; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_71 = 7'h47 == index ? tag_0_71 : _GEN_70; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_72 = 7'h48 == index ? tag_0_72 : _GEN_71; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_73 = 7'h49 == index ? tag_0_73 : _GEN_72; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_74 = 7'h4a == index ? tag_0_74 : _GEN_73; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_75 = 7'h4b == index ? tag_0_75 : _GEN_74; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_76 = 7'h4c == index ? tag_0_76 : _GEN_75; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_77 = 7'h4d == index ? tag_0_77 : _GEN_76; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_78 = 7'h4e == index ? tag_0_78 : _GEN_77; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_79 = 7'h4f == index ? tag_0_79 : _GEN_78; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_80 = 7'h50 == index ? tag_0_80 : _GEN_79; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_81 = 7'h51 == index ? tag_0_81 : _GEN_80; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_82 = 7'h52 == index ? tag_0_82 : _GEN_81; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_83 = 7'h53 == index ? tag_0_83 : _GEN_82; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_84 = 7'h54 == index ? tag_0_84 : _GEN_83; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_85 = 7'h55 == index ? tag_0_85 : _GEN_84; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_86 = 7'h56 == index ? tag_0_86 : _GEN_85; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_87 = 7'h57 == index ? tag_0_87 : _GEN_86; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_88 = 7'h58 == index ? tag_0_88 : _GEN_87; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_89 = 7'h59 == index ? tag_0_89 : _GEN_88; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_90 = 7'h5a == index ? tag_0_90 : _GEN_89; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_91 = 7'h5b == index ? tag_0_91 : _GEN_90; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_92 = 7'h5c == index ? tag_0_92 : _GEN_91; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_93 = 7'h5d == index ? tag_0_93 : _GEN_92; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_94 = 7'h5e == index ? tag_0_94 : _GEN_93; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_95 = 7'h5f == index ? tag_0_95 : _GEN_94; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_96 = 7'h60 == index ? tag_0_96 : _GEN_95; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_97 = 7'h61 == index ? tag_0_97 : _GEN_96; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_98 = 7'h62 == index ? tag_0_98 : _GEN_97; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_99 = 7'h63 == index ? tag_0_99 : _GEN_98; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_100 = 7'h64 == index ? tag_0_100 : _GEN_99; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_101 = 7'h65 == index ? tag_0_101 : _GEN_100; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_102 = 7'h66 == index ? tag_0_102 : _GEN_101; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_103 = 7'h67 == index ? tag_0_103 : _GEN_102; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_104 = 7'h68 == index ? tag_0_104 : _GEN_103; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_105 = 7'h69 == index ? tag_0_105 : _GEN_104; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_106 = 7'h6a == index ? tag_0_106 : _GEN_105; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_107 = 7'h6b == index ? tag_0_107 : _GEN_106; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_108 = 7'h6c == index ? tag_0_108 : _GEN_107; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_109 = 7'h6d == index ? tag_0_109 : _GEN_108; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_110 = 7'h6e == index ? tag_0_110 : _GEN_109; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_111 = 7'h6f == index ? tag_0_111 : _GEN_110; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_112 = 7'h70 == index ? tag_0_112 : _GEN_111; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_113 = 7'h71 == index ? tag_0_113 : _GEN_112; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_114 = 7'h72 == index ? tag_0_114 : _GEN_113; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_115 = 7'h73 == index ? tag_0_115 : _GEN_114; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_116 = 7'h74 == index ? tag_0_116 : _GEN_115; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_117 = 7'h75 == index ? tag_0_117 : _GEN_116; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_118 = 7'h76 == index ? tag_0_118 : _GEN_117; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_119 = 7'h77 == index ? tag_0_119 : _GEN_118; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_120 = 7'h78 == index ? tag_0_120 : _GEN_119; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_121 = 7'h79 == index ? tag_0_121 : _GEN_120; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_122 = 7'h7a == index ? tag_0_122 : _GEN_121; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_123 = 7'h7b == index ? tag_0_123 : _GEN_122; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_124 = 7'h7c == index ? tag_0_124 : _GEN_123; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_125 = 7'h7d == index ? tag_0_125 : _GEN_124; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_126 = 7'h7e == index ? tag_0_126 : _GEN_125; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_127 = 7'h7f == index ? tag_0_127 : _GEN_126; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_7706 = {{7'd0}, tag}; // @[i_cache.scala 34:24]
  wire  _GEN_129 = 7'h1 == index ? valid_0_1 : valid_0_0; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_130 = 7'h2 == index ? valid_0_2 : _GEN_129; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_131 = 7'h3 == index ? valid_0_3 : _GEN_130; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_132 = 7'h4 == index ? valid_0_4 : _GEN_131; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_133 = 7'h5 == index ? valid_0_5 : _GEN_132; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_134 = 7'h6 == index ? valid_0_6 : _GEN_133; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_135 = 7'h7 == index ? valid_0_7 : _GEN_134; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_136 = 7'h8 == index ? valid_0_8 : _GEN_135; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_137 = 7'h9 == index ? valid_0_9 : _GEN_136; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_138 = 7'ha == index ? valid_0_10 : _GEN_137; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_139 = 7'hb == index ? valid_0_11 : _GEN_138; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_140 = 7'hc == index ? valid_0_12 : _GEN_139; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_141 = 7'hd == index ? valid_0_13 : _GEN_140; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_142 = 7'he == index ? valid_0_14 : _GEN_141; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_143 = 7'hf == index ? valid_0_15 : _GEN_142; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_144 = 7'h10 == index ? valid_0_16 : _GEN_143; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_145 = 7'h11 == index ? valid_0_17 : _GEN_144; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_146 = 7'h12 == index ? valid_0_18 : _GEN_145; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_147 = 7'h13 == index ? valid_0_19 : _GEN_146; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_148 = 7'h14 == index ? valid_0_20 : _GEN_147; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_149 = 7'h15 == index ? valid_0_21 : _GEN_148; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_150 = 7'h16 == index ? valid_0_22 : _GEN_149; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_151 = 7'h17 == index ? valid_0_23 : _GEN_150; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_152 = 7'h18 == index ? valid_0_24 : _GEN_151; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_153 = 7'h19 == index ? valid_0_25 : _GEN_152; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_154 = 7'h1a == index ? valid_0_26 : _GEN_153; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_155 = 7'h1b == index ? valid_0_27 : _GEN_154; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_156 = 7'h1c == index ? valid_0_28 : _GEN_155; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_157 = 7'h1d == index ? valid_0_29 : _GEN_156; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_158 = 7'h1e == index ? valid_0_30 : _GEN_157; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_159 = 7'h1f == index ? valid_0_31 : _GEN_158; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_160 = 7'h20 == index ? valid_0_32 : _GEN_159; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_161 = 7'h21 == index ? valid_0_33 : _GEN_160; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_162 = 7'h22 == index ? valid_0_34 : _GEN_161; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_163 = 7'h23 == index ? valid_0_35 : _GEN_162; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_164 = 7'h24 == index ? valid_0_36 : _GEN_163; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_165 = 7'h25 == index ? valid_0_37 : _GEN_164; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_166 = 7'h26 == index ? valid_0_38 : _GEN_165; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_167 = 7'h27 == index ? valid_0_39 : _GEN_166; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_168 = 7'h28 == index ? valid_0_40 : _GEN_167; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_169 = 7'h29 == index ? valid_0_41 : _GEN_168; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_170 = 7'h2a == index ? valid_0_42 : _GEN_169; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_171 = 7'h2b == index ? valid_0_43 : _GEN_170; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_172 = 7'h2c == index ? valid_0_44 : _GEN_171; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_173 = 7'h2d == index ? valid_0_45 : _GEN_172; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_174 = 7'h2e == index ? valid_0_46 : _GEN_173; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_175 = 7'h2f == index ? valid_0_47 : _GEN_174; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_176 = 7'h30 == index ? valid_0_48 : _GEN_175; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_177 = 7'h31 == index ? valid_0_49 : _GEN_176; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_178 = 7'h32 == index ? valid_0_50 : _GEN_177; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_179 = 7'h33 == index ? valid_0_51 : _GEN_178; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_180 = 7'h34 == index ? valid_0_52 : _GEN_179; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_181 = 7'h35 == index ? valid_0_53 : _GEN_180; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_182 = 7'h36 == index ? valid_0_54 : _GEN_181; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_183 = 7'h37 == index ? valid_0_55 : _GEN_182; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_184 = 7'h38 == index ? valid_0_56 : _GEN_183; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_185 = 7'h39 == index ? valid_0_57 : _GEN_184; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_186 = 7'h3a == index ? valid_0_58 : _GEN_185; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_187 = 7'h3b == index ? valid_0_59 : _GEN_186; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_188 = 7'h3c == index ? valid_0_60 : _GEN_187; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_189 = 7'h3d == index ? valid_0_61 : _GEN_188; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_190 = 7'h3e == index ? valid_0_62 : _GEN_189; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_191 = 7'h3f == index ? valid_0_63 : _GEN_190; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_192 = 7'h40 == index ? valid_0_64 : _GEN_191; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_193 = 7'h41 == index ? valid_0_65 : _GEN_192; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_194 = 7'h42 == index ? valid_0_66 : _GEN_193; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_195 = 7'h43 == index ? valid_0_67 : _GEN_194; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_196 = 7'h44 == index ? valid_0_68 : _GEN_195; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_197 = 7'h45 == index ? valid_0_69 : _GEN_196; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_198 = 7'h46 == index ? valid_0_70 : _GEN_197; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_199 = 7'h47 == index ? valid_0_71 : _GEN_198; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_200 = 7'h48 == index ? valid_0_72 : _GEN_199; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_201 = 7'h49 == index ? valid_0_73 : _GEN_200; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_202 = 7'h4a == index ? valid_0_74 : _GEN_201; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_203 = 7'h4b == index ? valid_0_75 : _GEN_202; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_204 = 7'h4c == index ? valid_0_76 : _GEN_203; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_205 = 7'h4d == index ? valid_0_77 : _GEN_204; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_206 = 7'h4e == index ? valid_0_78 : _GEN_205; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_207 = 7'h4f == index ? valid_0_79 : _GEN_206; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_208 = 7'h50 == index ? valid_0_80 : _GEN_207; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_209 = 7'h51 == index ? valid_0_81 : _GEN_208; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_210 = 7'h52 == index ? valid_0_82 : _GEN_209; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_211 = 7'h53 == index ? valid_0_83 : _GEN_210; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_212 = 7'h54 == index ? valid_0_84 : _GEN_211; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_213 = 7'h55 == index ? valid_0_85 : _GEN_212; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_214 = 7'h56 == index ? valid_0_86 : _GEN_213; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_215 = 7'h57 == index ? valid_0_87 : _GEN_214; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_216 = 7'h58 == index ? valid_0_88 : _GEN_215; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_217 = 7'h59 == index ? valid_0_89 : _GEN_216; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_218 = 7'h5a == index ? valid_0_90 : _GEN_217; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_219 = 7'h5b == index ? valid_0_91 : _GEN_218; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_220 = 7'h5c == index ? valid_0_92 : _GEN_219; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_221 = 7'h5d == index ? valid_0_93 : _GEN_220; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_222 = 7'h5e == index ? valid_0_94 : _GEN_221; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_223 = 7'h5f == index ? valid_0_95 : _GEN_222; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_224 = 7'h60 == index ? valid_0_96 : _GEN_223; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_225 = 7'h61 == index ? valid_0_97 : _GEN_224; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_226 = 7'h62 == index ? valid_0_98 : _GEN_225; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_227 = 7'h63 == index ? valid_0_99 : _GEN_226; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_228 = 7'h64 == index ? valid_0_100 : _GEN_227; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_229 = 7'h65 == index ? valid_0_101 : _GEN_228; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_230 = 7'h66 == index ? valid_0_102 : _GEN_229; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_231 = 7'h67 == index ? valid_0_103 : _GEN_230; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_232 = 7'h68 == index ? valid_0_104 : _GEN_231; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_233 = 7'h69 == index ? valid_0_105 : _GEN_232; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_234 = 7'h6a == index ? valid_0_106 : _GEN_233; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_235 = 7'h6b == index ? valid_0_107 : _GEN_234; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_236 = 7'h6c == index ? valid_0_108 : _GEN_235; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_237 = 7'h6d == index ? valid_0_109 : _GEN_236; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_238 = 7'h6e == index ? valid_0_110 : _GEN_237; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_239 = 7'h6f == index ? valid_0_111 : _GEN_238; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_240 = 7'h70 == index ? valid_0_112 : _GEN_239; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_241 = 7'h71 == index ? valid_0_113 : _GEN_240; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_242 = 7'h72 == index ? valid_0_114 : _GEN_241; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_243 = 7'h73 == index ? valid_0_115 : _GEN_242; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_244 = 7'h74 == index ? valid_0_116 : _GEN_243; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_245 = 7'h75 == index ? valid_0_117 : _GEN_244; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_246 = 7'h76 == index ? valid_0_118 : _GEN_245; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_247 = 7'h77 == index ? valid_0_119 : _GEN_246; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_248 = 7'h78 == index ? valid_0_120 : _GEN_247; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_249 = 7'h79 == index ? valid_0_121 : _GEN_248; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_250 = 7'h7a == index ? valid_0_122 : _GEN_249; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_251 = 7'h7b == index ? valid_0_123 : _GEN_250; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_252 = 7'h7c == index ? valid_0_124 : _GEN_251; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_253 = 7'h7d == index ? valid_0_125 : _GEN_252; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_254 = 7'h7e == index ? valid_0_126 : _GEN_253; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_255 = 7'h7f == index ? valid_0_127 : _GEN_254; // @[i_cache.scala 34:{50,50}]
  wire  _T_2 = _GEN_127 == _GEN_7706 & _GEN_255; // @[i_cache.scala 34:33]
  wire [31:0] _GEN_258 = 7'h1 == index ? tag_1_1 : tag_1_0; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_259 = 7'h2 == index ? tag_1_2 : _GEN_258; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_260 = 7'h3 == index ? tag_1_3 : _GEN_259; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_261 = 7'h4 == index ? tag_1_4 : _GEN_260; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_262 = 7'h5 == index ? tag_1_5 : _GEN_261; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_263 = 7'h6 == index ? tag_1_6 : _GEN_262; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_264 = 7'h7 == index ? tag_1_7 : _GEN_263; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_265 = 7'h8 == index ? tag_1_8 : _GEN_264; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_266 = 7'h9 == index ? tag_1_9 : _GEN_265; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_267 = 7'ha == index ? tag_1_10 : _GEN_266; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_268 = 7'hb == index ? tag_1_11 : _GEN_267; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_269 = 7'hc == index ? tag_1_12 : _GEN_268; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_270 = 7'hd == index ? tag_1_13 : _GEN_269; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_271 = 7'he == index ? tag_1_14 : _GEN_270; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_272 = 7'hf == index ? tag_1_15 : _GEN_271; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_273 = 7'h10 == index ? tag_1_16 : _GEN_272; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_274 = 7'h11 == index ? tag_1_17 : _GEN_273; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_275 = 7'h12 == index ? tag_1_18 : _GEN_274; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_276 = 7'h13 == index ? tag_1_19 : _GEN_275; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_277 = 7'h14 == index ? tag_1_20 : _GEN_276; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_278 = 7'h15 == index ? tag_1_21 : _GEN_277; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_279 = 7'h16 == index ? tag_1_22 : _GEN_278; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_280 = 7'h17 == index ? tag_1_23 : _GEN_279; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_281 = 7'h18 == index ? tag_1_24 : _GEN_280; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_282 = 7'h19 == index ? tag_1_25 : _GEN_281; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_283 = 7'h1a == index ? tag_1_26 : _GEN_282; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_284 = 7'h1b == index ? tag_1_27 : _GEN_283; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_285 = 7'h1c == index ? tag_1_28 : _GEN_284; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_286 = 7'h1d == index ? tag_1_29 : _GEN_285; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_287 = 7'h1e == index ? tag_1_30 : _GEN_286; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_288 = 7'h1f == index ? tag_1_31 : _GEN_287; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_289 = 7'h20 == index ? tag_1_32 : _GEN_288; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_290 = 7'h21 == index ? tag_1_33 : _GEN_289; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_291 = 7'h22 == index ? tag_1_34 : _GEN_290; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_292 = 7'h23 == index ? tag_1_35 : _GEN_291; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_293 = 7'h24 == index ? tag_1_36 : _GEN_292; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_294 = 7'h25 == index ? tag_1_37 : _GEN_293; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_295 = 7'h26 == index ? tag_1_38 : _GEN_294; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_296 = 7'h27 == index ? tag_1_39 : _GEN_295; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_297 = 7'h28 == index ? tag_1_40 : _GEN_296; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_298 = 7'h29 == index ? tag_1_41 : _GEN_297; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_299 = 7'h2a == index ? tag_1_42 : _GEN_298; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_300 = 7'h2b == index ? tag_1_43 : _GEN_299; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_301 = 7'h2c == index ? tag_1_44 : _GEN_300; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_302 = 7'h2d == index ? tag_1_45 : _GEN_301; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_303 = 7'h2e == index ? tag_1_46 : _GEN_302; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_304 = 7'h2f == index ? tag_1_47 : _GEN_303; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_305 = 7'h30 == index ? tag_1_48 : _GEN_304; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_306 = 7'h31 == index ? tag_1_49 : _GEN_305; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_307 = 7'h32 == index ? tag_1_50 : _GEN_306; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_308 = 7'h33 == index ? tag_1_51 : _GEN_307; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_309 = 7'h34 == index ? tag_1_52 : _GEN_308; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_310 = 7'h35 == index ? tag_1_53 : _GEN_309; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_311 = 7'h36 == index ? tag_1_54 : _GEN_310; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_312 = 7'h37 == index ? tag_1_55 : _GEN_311; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_313 = 7'h38 == index ? tag_1_56 : _GEN_312; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_314 = 7'h39 == index ? tag_1_57 : _GEN_313; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_315 = 7'h3a == index ? tag_1_58 : _GEN_314; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_316 = 7'h3b == index ? tag_1_59 : _GEN_315; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_317 = 7'h3c == index ? tag_1_60 : _GEN_316; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_318 = 7'h3d == index ? tag_1_61 : _GEN_317; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_319 = 7'h3e == index ? tag_1_62 : _GEN_318; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_320 = 7'h3f == index ? tag_1_63 : _GEN_319; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_321 = 7'h40 == index ? tag_1_64 : _GEN_320; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_322 = 7'h41 == index ? tag_1_65 : _GEN_321; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_323 = 7'h42 == index ? tag_1_66 : _GEN_322; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_324 = 7'h43 == index ? tag_1_67 : _GEN_323; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_325 = 7'h44 == index ? tag_1_68 : _GEN_324; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_326 = 7'h45 == index ? tag_1_69 : _GEN_325; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_327 = 7'h46 == index ? tag_1_70 : _GEN_326; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_328 = 7'h47 == index ? tag_1_71 : _GEN_327; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_329 = 7'h48 == index ? tag_1_72 : _GEN_328; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_330 = 7'h49 == index ? tag_1_73 : _GEN_329; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_331 = 7'h4a == index ? tag_1_74 : _GEN_330; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_332 = 7'h4b == index ? tag_1_75 : _GEN_331; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_333 = 7'h4c == index ? tag_1_76 : _GEN_332; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_334 = 7'h4d == index ? tag_1_77 : _GEN_333; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_335 = 7'h4e == index ? tag_1_78 : _GEN_334; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_336 = 7'h4f == index ? tag_1_79 : _GEN_335; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_337 = 7'h50 == index ? tag_1_80 : _GEN_336; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_338 = 7'h51 == index ? tag_1_81 : _GEN_337; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_339 = 7'h52 == index ? tag_1_82 : _GEN_338; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_340 = 7'h53 == index ? tag_1_83 : _GEN_339; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_341 = 7'h54 == index ? tag_1_84 : _GEN_340; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_342 = 7'h55 == index ? tag_1_85 : _GEN_341; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_343 = 7'h56 == index ? tag_1_86 : _GEN_342; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_344 = 7'h57 == index ? tag_1_87 : _GEN_343; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_345 = 7'h58 == index ? tag_1_88 : _GEN_344; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_346 = 7'h59 == index ? tag_1_89 : _GEN_345; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_347 = 7'h5a == index ? tag_1_90 : _GEN_346; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_348 = 7'h5b == index ? tag_1_91 : _GEN_347; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_349 = 7'h5c == index ? tag_1_92 : _GEN_348; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_350 = 7'h5d == index ? tag_1_93 : _GEN_349; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_351 = 7'h5e == index ? tag_1_94 : _GEN_350; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_352 = 7'h5f == index ? tag_1_95 : _GEN_351; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_353 = 7'h60 == index ? tag_1_96 : _GEN_352; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_354 = 7'h61 == index ? tag_1_97 : _GEN_353; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_355 = 7'h62 == index ? tag_1_98 : _GEN_354; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_356 = 7'h63 == index ? tag_1_99 : _GEN_355; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_357 = 7'h64 == index ? tag_1_100 : _GEN_356; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_358 = 7'h65 == index ? tag_1_101 : _GEN_357; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_359 = 7'h66 == index ? tag_1_102 : _GEN_358; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_360 = 7'h67 == index ? tag_1_103 : _GEN_359; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_361 = 7'h68 == index ? tag_1_104 : _GEN_360; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_362 = 7'h69 == index ? tag_1_105 : _GEN_361; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_363 = 7'h6a == index ? tag_1_106 : _GEN_362; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_364 = 7'h6b == index ? tag_1_107 : _GEN_363; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_365 = 7'h6c == index ? tag_1_108 : _GEN_364; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_366 = 7'h6d == index ? tag_1_109 : _GEN_365; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_367 = 7'h6e == index ? tag_1_110 : _GEN_366; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_368 = 7'h6f == index ? tag_1_111 : _GEN_367; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_369 = 7'h70 == index ? tag_1_112 : _GEN_368; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_370 = 7'h71 == index ? tag_1_113 : _GEN_369; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_371 = 7'h72 == index ? tag_1_114 : _GEN_370; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_372 = 7'h73 == index ? tag_1_115 : _GEN_371; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_373 = 7'h74 == index ? tag_1_116 : _GEN_372; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_374 = 7'h75 == index ? tag_1_117 : _GEN_373; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_375 = 7'h76 == index ? tag_1_118 : _GEN_374; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_376 = 7'h77 == index ? tag_1_119 : _GEN_375; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_377 = 7'h78 == index ? tag_1_120 : _GEN_376; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_378 = 7'h79 == index ? tag_1_121 : _GEN_377; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_379 = 7'h7a == index ? tag_1_122 : _GEN_378; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_380 = 7'h7b == index ? tag_1_123 : _GEN_379; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_381 = 7'h7c == index ? tag_1_124 : _GEN_380; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_382 = 7'h7d == index ? tag_1_125 : _GEN_381; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_383 = 7'h7e == index ? tag_1_126 : _GEN_382; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_384 = 7'h7f == index ? tag_1_127 : _GEN_383; // @[i_cache.scala 39:{24,24}]
  wire  _GEN_386 = 7'h1 == index ? valid_1_1 : valid_1_0; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_387 = 7'h2 == index ? valid_1_2 : _GEN_386; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_388 = 7'h3 == index ? valid_1_3 : _GEN_387; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_389 = 7'h4 == index ? valid_1_4 : _GEN_388; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_390 = 7'h5 == index ? valid_1_5 : _GEN_389; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_391 = 7'h6 == index ? valid_1_6 : _GEN_390; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_392 = 7'h7 == index ? valid_1_7 : _GEN_391; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_393 = 7'h8 == index ? valid_1_8 : _GEN_392; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_394 = 7'h9 == index ? valid_1_9 : _GEN_393; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_395 = 7'ha == index ? valid_1_10 : _GEN_394; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_396 = 7'hb == index ? valid_1_11 : _GEN_395; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_397 = 7'hc == index ? valid_1_12 : _GEN_396; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_398 = 7'hd == index ? valid_1_13 : _GEN_397; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_399 = 7'he == index ? valid_1_14 : _GEN_398; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_400 = 7'hf == index ? valid_1_15 : _GEN_399; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_401 = 7'h10 == index ? valid_1_16 : _GEN_400; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_402 = 7'h11 == index ? valid_1_17 : _GEN_401; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_403 = 7'h12 == index ? valid_1_18 : _GEN_402; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_404 = 7'h13 == index ? valid_1_19 : _GEN_403; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_405 = 7'h14 == index ? valid_1_20 : _GEN_404; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_406 = 7'h15 == index ? valid_1_21 : _GEN_405; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_407 = 7'h16 == index ? valid_1_22 : _GEN_406; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_408 = 7'h17 == index ? valid_1_23 : _GEN_407; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_409 = 7'h18 == index ? valid_1_24 : _GEN_408; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_410 = 7'h19 == index ? valid_1_25 : _GEN_409; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_411 = 7'h1a == index ? valid_1_26 : _GEN_410; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_412 = 7'h1b == index ? valid_1_27 : _GEN_411; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_413 = 7'h1c == index ? valid_1_28 : _GEN_412; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_414 = 7'h1d == index ? valid_1_29 : _GEN_413; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_415 = 7'h1e == index ? valid_1_30 : _GEN_414; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_416 = 7'h1f == index ? valid_1_31 : _GEN_415; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_417 = 7'h20 == index ? valid_1_32 : _GEN_416; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_418 = 7'h21 == index ? valid_1_33 : _GEN_417; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_419 = 7'h22 == index ? valid_1_34 : _GEN_418; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_420 = 7'h23 == index ? valid_1_35 : _GEN_419; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_421 = 7'h24 == index ? valid_1_36 : _GEN_420; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_422 = 7'h25 == index ? valid_1_37 : _GEN_421; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_423 = 7'h26 == index ? valid_1_38 : _GEN_422; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_424 = 7'h27 == index ? valid_1_39 : _GEN_423; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_425 = 7'h28 == index ? valid_1_40 : _GEN_424; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_426 = 7'h29 == index ? valid_1_41 : _GEN_425; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_427 = 7'h2a == index ? valid_1_42 : _GEN_426; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_428 = 7'h2b == index ? valid_1_43 : _GEN_427; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_429 = 7'h2c == index ? valid_1_44 : _GEN_428; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_430 = 7'h2d == index ? valid_1_45 : _GEN_429; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_431 = 7'h2e == index ? valid_1_46 : _GEN_430; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_432 = 7'h2f == index ? valid_1_47 : _GEN_431; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_433 = 7'h30 == index ? valid_1_48 : _GEN_432; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_434 = 7'h31 == index ? valid_1_49 : _GEN_433; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_435 = 7'h32 == index ? valid_1_50 : _GEN_434; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_436 = 7'h33 == index ? valid_1_51 : _GEN_435; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_437 = 7'h34 == index ? valid_1_52 : _GEN_436; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_438 = 7'h35 == index ? valid_1_53 : _GEN_437; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_439 = 7'h36 == index ? valid_1_54 : _GEN_438; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_440 = 7'h37 == index ? valid_1_55 : _GEN_439; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_441 = 7'h38 == index ? valid_1_56 : _GEN_440; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_442 = 7'h39 == index ? valid_1_57 : _GEN_441; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_443 = 7'h3a == index ? valid_1_58 : _GEN_442; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_444 = 7'h3b == index ? valid_1_59 : _GEN_443; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_445 = 7'h3c == index ? valid_1_60 : _GEN_444; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_446 = 7'h3d == index ? valid_1_61 : _GEN_445; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_447 = 7'h3e == index ? valid_1_62 : _GEN_446; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_448 = 7'h3f == index ? valid_1_63 : _GEN_447; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_449 = 7'h40 == index ? valid_1_64 : _GEN_448; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_450 = 7'h41 == index ? valid_1_65 : _GEN_449; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_451 = 7'h42 == index ? valid_1_66 : _GEN_450; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_452 = 7'h43 == index ? valid_1_67 : _GEN_451; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_453 = 7'h44 == index ? valid_1_68 : _GEN_452; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_454 = 7'h45 == index ? valid_1_69 : _GEN_453; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_455 = 7'h46 == index ? valid_1_70 : _GEN_454; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_456 = 7'h47 == index ? valid_1_71 : _GEN_455; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_457 = 7'h48 == index ? valid_1_72 : _GEN_456; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_458 = 7'h49 == index ? valid_1_73 : _GEN_457; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_459 = 7'h4a == index ? valid_1_74 : _GEN_458; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_460 = 7'h4b == index ? valid_1_75 : _GEN_459; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_461 = 7'h4c == index ? valid_1_76 : _GEN_460; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_462 = 7'h4d == index ? valid_1_77 : _GEN_461; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_463 = 7'h4e == index ? valid_1_78 : _GEN_462; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_464 = 7'h4f == index ? valid_1_79 : _GEN_463; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_465 = 7'h50 == index ? valid_1_80 : _GEN_464; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_466 = 7'h51 == index ? valid_1_81 : _GEN_465; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_467 = 7'h52 == index ? valid_1_82 : _GEN_466; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_468 = 7'h53 == index ? valid_1_83 : _GEN_467; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_469 = 7'h54 == index ? valid_1_84 : _GEN_468; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_470 = 7'h55 == index ? valid_1_85 : _GEN_469; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_471 = 7'h56 == index ? valid_1_86 : _GEN_470; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_472 = 7'h57 == index ? valid_1_87 : _GEN_471; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_473 = 7'h58 == index ? valid_1_88 : _GEN_472; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_474 = 7'h59 == index ? valid_1_89 : _GEN_473; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_475 = 7'h5a == index ? valid_1_90 : _GEN_474; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_476 = 7'h5b == index ? valid_1_91 : _GEN_475; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_477 = 7'h5c == index ? valid_1_92 : _GEN_476; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_478 = 7'h5d == index ? valid_1_93 : _GEN_477; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_479 = 7'h5e == index ? valid_1_94 : _GEN_478; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_480 = 7'h5f == index ? valid_1_95 : _GEN_479; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_481 = 7'h60 == index ? valid_1_96 : _GEN_480; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_482 = 7'h61 == index ? valid_1_97 : _GEN_481; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_483 = 7'h62 == index ? valid_1_98 : _GEN_482; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_484 = 7'h63 == index ? valid_1_99 : _GEN_483; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_485 = 7'h64 == index ? valid_1_100 : _GEN_484; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_486 = 7'h65 == index ? valid_1_101 : _GEN_485; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_487 = 7'h66 == index ? valid_1_102 : _GEN_486; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_488 = 7'h67 == index ? valid_1_103 : _GEN_487; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_489 = 7'h68 == index ? valid_1_104 : _GEN_488; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_490 = 7'h69 == index ? valid_1_105 : _GEN_489; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_491 = 7'h6a == index ? valid_1_106 : _GEN_490; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_492 = 7'h6b == index ? valid_1_107 : _GEN_491; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_493 = 7'h6c == index ? valid_1_108 : _GEN_492; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_494 = 7'h6d == index ? valid_1_109 : _GEN_493; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_495 = 7'h6e == index ? valid_1_110 : _GEN_494; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_496 = 7'h6f == index ? valid_1_111 : _GEN_495; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_497 = 7'h70 == index ? valid_1_112 : _GEN_496; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_498 = 7'h71 == index ? valid_1_113 : _GEN_497; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_499 = 7'h72 == index ? valid_1_114 : _GEN_498; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_500 = 7'h73 == index ? valid_1_115 : _GEN_499; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_501 = 7'h74 == index ? valid_1_116 : _GEN_500; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_502 = 7'h75 == index ? valid_1_117 : _GEN_501; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_503 = 7'h76 == index ? valid_1_118 : _GEN_502; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_504 = 7'h77 == index ? valid_1_119 : _GEN_503; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_505 = 7'h78 == index ? valid_1_120 : _GEN_504; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_506 = 7'h79 == index ? valid_1_121 : _GEN_505; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_507 = 7'h7a == index ? valid_1_122 : _GEN_506; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_508 = 7'h7b == index ? valid_1_123 : _GEN_507; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_509 = 7'h7c == index ? valid_1_124 : _GEN_508; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_510 = 7'h7d == index ? valid_1_125 : _GEN_509; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_511 = 7'h7e == index ? valid_1_126 : _GEN_510; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_512 = 7'h7f == index ? valid_1_127 : _GEN_511; // @[i_cache.scala 39:{50,50}]
  wire  _T_5 = _GEN_384 == _GEN_7706 & _GEN_512; // @[i_cache.scala 39:33]
  reg [2:0] state; // @[i_cache.scala 53:24]
  wire [2:0] _GEN_517 = io_from_ifu_rready ? 3'h0 : state; // @[i_cache.scala 53:24 64:41 65:27]
  wire [2:0] _GEN_518 = way1_hit ? _GEN_517 : 3'h2; // @[i_cache.scala 68:33 73:23]
  wire [2:0] _GEN_520 = io_from_axi_rvalid ? 3'h3 : state; // @[i_cache.scala 77:37 78:23 53:24]
  wire [63:0] _GEN_521 = io_from_axi_rvalid ? io_from_axi_rdata : receive_data; // @[i_cache.scala 80:37 81:30 27:31]
  wire [63:0] _GEN_522 = 7'h0 == index ? receive_data : ram_0_0; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_523 = 7'h1 == index ? receive_data : ram_0_1; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_524 = 7'h2 == index ? receive_data : ram_0_2; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_525 = 7'h3 == index ? receive_data : ram_0_3; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_526 = 7'h4 == index ? receive_data : ram_0_4; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_527 = 7'h5 == index ? receive_data : ram_0_5; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_528 = 7'h6 == index ? receive_data : ram_0_6; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_529 = 7'h7 == index ? receive_data : ram_0_7; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_530 = 7'h8 == index ? receive_data : ram_0_8; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_531 = 7'h9 == index ? receive_data : ram_0_9; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_532 = 7'ha == index ? receive_data : ram_0_10; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_533 = 7'hb == index ? receive_data : ram_0_11; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_534 = 7'hc == index ? receive_data : ram_0_12; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_535 = 7'hd == index ? receive_data : ram_0_13; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_536 = 7'he == index ? receive_data : ram_0_14; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_537 = 7'hf == index ? receive_data : ram_0_15; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_538 = 7'h10 == index ? receive_data : ram_0_16; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_539 = 7'h11 == index ? receive_data : ram_0_17; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_540 = 7'h12 == index ? receive_data : ram_0_18; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_541 = 7'h13 == index ? receive_data : ram_0_19; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_542 = 7'h14 == index ? receive_data : ram_0_20; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_543 = 7'h15 == index ? receive_data : ram_0_21; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_544 = 7'h16 == index ? receive_data : ram_0_22; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_545 = 7'h17 == index ? receive_data : ram_0_23; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_546 = 7'h18 == index ? receive_data : ram_0_24; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_547 = 7'h19 == index ? receive_data : ram_0_25; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_548 = 7'h1a == index ? receive_data : ram_0_26; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_549 = 7'h1b == index ? receive_data : ram_0_27; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_550 = 7'h1c == index ? receive_data : ram_0_28; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_551 = 7'h1d == index ? receive_data : ram_0_29; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_552 = 7'h1e == index ? receive_data : ram_0_30; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_553 = 7'h1f == index ? receive_data : ram_0_31; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_554 = 7'h20 == index ? receive_data : ram_0_32; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_555 = 7'h21 == index ? receive_data : ram_0_33; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_556 = 7'h22 == index ? receive_data : ram_0_34; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_557 = 7'h23 == index ? receive_data : ram_0_35; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_558 = 7'h24 == index ? receive_data : ram_0_36; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_559 = 7'h25 == index ? receive_data : ram_0_37; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_560 = 7'h26 == index ? receive_data : ram_0_38; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_561 = 7'h27 == index ? receive_data : ram_0_39; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_562 = 7'h28 == index ? receive_data : ram_0_40; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_563 = 7'h29 == index ? receive_data : ram_0_41; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_564 = 7'h2a == index ? receive_data : ram_0_42; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_565 = 7'h2b == index ? receive_data : ram_0_43; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_566 = 7'h2c == index ? receive_data : ram_0_44; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_567 = 7'h2d == index ? receive_data : ram_0_45; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_568 = 7'h2e == index ? receive_data : ram_0_46; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_569 = 7'h2f == index ? receive_data : ram_0_47; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_570 = 7'h30 == index ? receive_data : ram_0_48; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_571 = 7'h31 == index ? receive_data : ram_0_49; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_572 = 7'h32 == index ? receive_data : ram_0_50; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_573 = 7'h33 == index ? receive_data : ram_0_51; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_574 = 7'h34 == index ? receive_data : ram_0_52; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_575 = 7'h35 == index ? receive_data : ram_0_53; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_576 = 7'h36 == index ? receive_data : ram_0_54; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_577 = 7'h37 == index ? receive_data : ram_0_55; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_578 = 7'h38 == index ? receive_data : ram_0_56; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_579 = 7'h39 == index ? receive_data : ram_0_57; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_580 = 7'h3a == index ? receive_data : ram_0_58; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_581 = 7'h3b == index ? receive_data : ram_0_59; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_582 = 7'h3c == index ? receive_data : ram_0_60; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_583 = 7'h3d == index ? receive_data : ram_0_61; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_584 = 7'h3e == index ? receive_data : ram_0_62; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_585 = 7'h3f == index ? receive_data : ram_0_63; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_586 = 7'h40 == index ? receive_data : ram_0_64; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_587 = 7'h41 == index ? receive_data : ram_0_65; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_588 = 7'h42 == index ? receive_data : ram_0_66; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_589 = 7'h43 == index ? receive_data : ram_0_67; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_590 = 7'h44 == index ? receive_data : ram_0_68; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_591 = 7'h45 == index ? receive_data : ram_0_69; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_592 = 7'h46 == index ? receive_data : ram_0_70; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_593 = 7'h47 == index ? receive_data : ram_0_71; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_594 = 7'h48 == index ? receive_data : ram_0_72; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_595 = 7'h49 == index ? receive_data : ram_0_73; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_596 = 7'h4a == index ? receive_data : ram_0_74; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_597 = 7'h4b == index ? receive_data : ram_0_75; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_598 = 7'h4c == index ? receive_data : ram_0_76; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_599 = 7'h4d == index ? receive_data : ram_0_77; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_600 = 7'h4e == index ? receive_data : ram_0_78; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_601 = 7'h4f == index ? receive_data : ram_0_79; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_602 = 7'h50 == index ? receive_data : ram_0_80; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_603 = 7'h51 == index ? receive_data : ram_0_81; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_604 = 7'h52 == index ? receive_data : ram_0_82; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_605 = 7'h53 == index ? receive_data : ram_0_83; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_606 = 7'h54 == index ? receive_data : ram_0_84; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_607 = 7'h55 == index ? receive_data : ram_0_85; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_608 = 7'h56 == index ? receive_data : ram_0_86; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_609 = 7'h57 == index ? receive_data : ram_0_87; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_610 = 7'h58 == index ? receive_data : ram_0_88; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_611 = 7'h59 == index ? receive_data : ram_0_89; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_612 = 7'h5a == index ? receive_data : ram_0_90; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_613 = 7'h5b == index ? receive_data : ram_0_91; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_614 = 7'h5c == index ? receive_data : ram_0_92; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_615 = 7'h5d == index ? receive_data : ram_0_93; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_616 = 7'h5e == index ? receive_data : ram_0_94; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_617 = 7'h5f == index ? receive_data : ram_0_95; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_618 = 7'h60 == index ? receive_data : ram_0_96; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_619 = 7'h61 == index ? receive_data : ram_0_97; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_620 = 7'h62 == index ? receive_data : ram_0_98; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_621 = 7'h63 == index ? receive_data : ram_0_99; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_622 = 7'h64 == index ? receive_data : ram_0_100; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_623 = 7'h65 == index ? receive_data : ram_0_101; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_624 = 7'h66 == index ? receive_data : ram_0_102; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_625 = 7'h67 == index ? receive_data : ram_0_103; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_626 = 7'h68 == index ? receive_data : ram_0_104; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_627 = 7'h69 == index ? receive_data : ram_0_105; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_628 = 7'h6a == index ? receive_data : ram_0_106; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_629 = 7'h6b == index ? receive_data : ram_0_107; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_630 = 7'h6c == index ? receive_data : ram_0_108; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_631 = 7'h6d == index ? receive_data : ram_0_109; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_632 = 7'h6e == index ? receive_data : ram_0_110; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_633 = 7'h6f == index ? receive_data : ram_0_111; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_634 = 7'h70 == index ? receive_data : ram_0_112; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_635 = 7'h71 == index ? receive_data : ram_0_113; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_636 = 7'h72 == index ? receive_data : ram_0_114; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_637 = 7'h73 == index ? receive_data : ram_0_115; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_638 = 7'h74 == index ? receive_data : ram_0_116; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_639 = 7'h75 == index ? receive_data : ram_0_117; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_640 = 7'h76 == index ? receive_data : ram_0_118; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_641 = 7'h77 == index ? receive_data : ram_0_119; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_642 = 7'h78 == index ? receive_data : ram_0_120; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_643 = 7'h79 == index ? receive_data : ram_0_121; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_644 = 7'h7a == index ? receive_data : ram_0_122; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_645 = 7'h7b == index ? receive_data : ram_0_123; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_646 = 7'h7c == index ? receive_data : ram_0_124; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_647 = 7'h7d == index ? receive_data : ram_0_125; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_648 = 7'h7e == index ? receive_data : ram_0_126; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_649 = 7'h7f == index ? receive_data : ram_0_127; // @[i_cache.scala 17:24 87:{30,30}]
  wire [31:0] _GEN_650 = 7'h0 == index ? _GEN_7706 : tag_0_0; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_651 = 7'h1 == index ? _GEN_7706 : tag_0_1; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_652 = 7'h2 == index ? _GEN_7706 : tag_0_2; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_653 = 7'h3 == index ? _GEN_7706 : tag_0_3; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_654 = 7'h4 == index ? _GEN_7706 : tag_0_4; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_655 = 7'h5 == index ? _GEN_7706 : tag_0_5; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_656 = 7'h6 == index ? _GEN_7706 : tag_0_6; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_657 = 7'h7 == index ? _GEN_7706 : tag_0_7; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_658 = 7'h8 == index ? _GEN_7706 : tag_0_8; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_659 = 7'h9 == index ? _GEN_7706 : tag_0_9; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_660 = 7'ha == index ? _GEN_7706 : tag_0_10; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_661 = 7'hb == index ? _GEN_7706 : tag_0_11; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_662 = 7'hc == index ? _GEN_7706 : tag_0_12; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_663 = 7'hd == index ? _GEN_7706 : tag_0_13; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_664 = 7'he == index ? _GEN_7706 : tag_0_14; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_665 = 7'hf == index ? _GEN_7706 : tag_0_15; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_666 = 7'h10 == index ? _GEN_7706 : tag_0_16; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_667 = 7'h11 == index ? _GEN_7706 : tag_0_17; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_668 = 7'h12 == index ? _GEN_7706 : tag_0_18; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_669 = 7'h13 == index ? _GEN_7706 : tag_0_19; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_670 = 7'h14 == index ? _GEN_7706 : tag_0_20; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_671 = 7'h15 == index ? _GEN_7706 : tag_0_21; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_672 = 7'h16 == index ? _GEN_7706 : tag_0_22; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_673 = 7'h17 == index ? _GEN_7706 : tag_0_23; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_674 = 7'h18 == index ? _GEN_7706 : tag_0_24; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_675 = 7'h19 == index ? _GEN_7706 : tag_0_25; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_676 = 7'h1a == index ? _GEN_7706 : tag_0_26; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_677 = 7'h1b == index ? _GEN_7706 : tag_0_27; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_678 = 7'h1c == index ? _GEN_7706 : tag_0_28; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_679 = 7'h1d == index ? _GEN_7706 : tag_0_29; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_680 = 7'h1e == index ? _GEN_7706 : tag_0_30; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_681 = 7'h1f == index ? _GEN_7706 : tag_0_31; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_682 = 7'h20 == index ? _GEN_7706 : tag_0_32; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_683 = 7'h21 == index ? _GEN_7706 : tag_0_33; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_684 = 7'h22 == index ? _GEN_7706 : tag_0_34; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_685 = 7'h23 == index ? _GEN_7706 : tag_0_35; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_686 = 7'h24 == index ? _GEN_7706 : tag_0_36; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_687 = 7'h25 == index ? _GEN_7706 : tag_0_37; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_688 = 7'h26 == index ? _GEN_7706 : tag_0_38; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_689 = 7'h27 == index ? _GEN_7706 : tag_0_39; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_690 = 7'h28 == index ? _GEN_7706 : tag_0_40; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_691 = 7'h29 == index ? _GEN_7706 : tag_0_41; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_692 = 7'h2a == index ? _GEN_7706 : tag_0_42; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_693 = 7'h2b == index ? _GEN_7706 : tag_0_43; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_694 = 7'h2c == index ? _GEN_7706 : tag_0_44; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_695 = 7'h2d == index ? _GEN_7706 : tag_0_45; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_696 = 7'h2e == index ? _GEN_7706 : tag_0_46; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_697 = 7'h2f == index ? _GEN_7706 : tag_0_47; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_698 = 7'h30 == index ? _GEN_7706 : tag_0_48; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_699 = 7'h31 == index ? _GEN_7706 : tag_0_49; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_700 = 7'h32 == index ? _GEN_7706 : tag_0_50; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_701 = 7'h33 == index ? _GEN_7706 : tag_0_51; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_702 = 7'h34 == index ? _GEN_7706 : tag_0_52; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_703 = 7'h35 == index ? _GEN_7706 : tag_0_53; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_704 = 7'h36 == index ? _GEN_7706 : tag_0_54; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_705 = 7'h37 == index ? _GEN_7706 : tag_0_55; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_706 = 7'h38 == index ? _GEN_7706 : tag_0_56; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_707 = 7'h39 == index ? _GEN_7706 : tag_0_57; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_708 = 7'h3a == index ? _GEN_7706 : tag_0_58; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_709 = 7'h3b == index ? _GEN_7706 : tag_0_59; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_710 = 7'h3c == index ? _GEN_7706 : tag_0_60; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_711 = 7'h3d == index ? _GEN_7706 : tag_0_61; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_712 = 7'h3e == index ? _GEN_7706 : tag_0_62; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_713 = 7'h3f == index ? _GEN_7706 : tag_0_63; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_714 = 7'h40 == index ? _GEN_7706 : tag_0_64; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_715 = 7'h41 == index ? _GEN_7706 : tag_0_65; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_716 = 7'h42 == index ? _GEN_7706 : tag_0_66; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_717 = 7'h43 == index ? _GEN_7706 : tag_0_67; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_718 = 7'h44 == index ? _GEN_7706 : tag_0_68; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_719 = 7'h45 == index ? _GEN_7706 : tag_0_69; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_720 = 7'h46 == index ? _GEN_7706 : tag_0_70; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_721 = 7'h47 == index ? _GEN_7706 : tag_0_71; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_722 = 7'h48 == index ? _GEN_7706 : tag_0_72; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_723 = 7'h49 == index ? _GEN_7706 : tag_0_73; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_724 = 7'h4a == index ? _GEN_7706 : tag_0_74; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_725 = 7'h4b == index ? _GEN_7706 : tag_0_75; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_726 = 7'h4c == index ? _GEN_7706 : tag_0_76; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_727 = 7'h4d == index ? _GEN_7706 : tag_0_77; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_728 = 7'h4e == index ? _GEN_7706 : tag_0_78; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_729 = 7'h4f == index ? _GEN_7706 : tag_0_79; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_730 = 7'h50 == index ? _GEN_7706 : tag_0_80; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_731 = 7'h51 == index ? _GEN_7706 : tag_0_81; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_732 = 7'h52 == index ? _GEN_7706 : tag_0_82; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_733 = 7'h53 == index ? _GEN_7706 : tag_0_83; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_734 = 7'h54 == index ? _GEN_7706 : tag_0_84; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_735 = 7'h55 == index ? _GEN_7706 : tag_0_85; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_736 = 7'h56 == index ? _GEN_7706 : tag_0_86; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_737 = 7'h57 == index ? _GEN_7706 : tag_0_87; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_738 = 7'h58 == index ? _GEN_7706 : tag_0_88; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_739 = 7'h59 == index ? _GEN_7706 : tag_0_89; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_740 = 7'h5a == index ? _GEN_7706 : tag_0_90; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_741 = 7'h5b == index ? _GEN_7706 : tag_0_91; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_742 = 7'h5c == index ? _GEN_7706 : tag_0_92; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_743 = 7'h5d == index ? _GEN_7706 : tag_0_93; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_744 = 7'h5e == index ? _GEN_7706 : tag_0_94; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_745 = 7'h5f == index ? _GEN_7706 : tag_0_95; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_746 = 7'h60 == index ? _GEN_7706 : tag_0_96; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_747 = 7'h61 == index ? _GEN_7706 : tag_0_97; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_748 = 7'h62 == index ? _GEN_7706 : tag_0_98; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_749 = 7'h63 == index ? _GEN_7706 : tag_0_99; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_750 = 7'h64 == index ? _GEN_7706 : tag_0_100; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_751 = 7'h65 == index ? _GEN_7706 : tag_0_101; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_752 = 7'h66 == index ? _GEN_7706 : tag_0_102; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_753 = 7'h67 == index ? _GEN_7706 : tag_0_103; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_754 = 7'h68 == index ? _GEN_7706 : tag_0_104; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_755 = 7'h69 == index ? _GEN_7706 : tag_0_105; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_756 = 7'h6a == index ? _GEN_7706 : tag_0_106; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_757 = 7'h6b == index ? _GEN_7706 : tag_0_107; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_758 = 7'h6c == index ? _GEN_7706 : tag_0_108; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_759 = 7'h6d == index ? _GEN_7706 : tag_0_109; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_760 = 7'h6e == index ? _GEN_7706 : tag_0_110; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_761 = 7'h6f == index ? _GEN_7706 : tag_0_111; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_762 = 7'h70 == index ? _GEN_7706 : tag_0_112; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_763 = 7'h71 == index ? _GEN_7706 : tag_0_113; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_764 = 7'h72 == index ? _GEN_7706 : tag_0_114; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_765 = 7'h73 == index ? _GEN_7706 : tag_0_115; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_766 = 7'h74 == index ? _GEN_7706 : tag_0_116; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_767 = 7'h75 == index ? _GEN_7706 : tag_0_117; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_768 = 7'h76 == index ? _GEN_7706 : tag_0_118; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_769 = 7'h77 == index ? _GEN_7706 : tag_0_119; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_770 = 7'h78 == index ? _GEN_7706 : tag_0_120; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_771 = 7'h79 == index ? _GEN_7706 : tag_0_121; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_772 = 7'h7a == index ? _GEN_7706 : tag_0_122; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_773 = 7'h7b == index ? _GEN_7706 : tag_0_123; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_774 = 7'h7c == index ? _GEN_7706 : tag_0_124; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_775 = 7'h7d == index ? _GEN_7706 : tag_0_125; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_776 = 7'h7e == index ? _GEN_7706 : tag_0_126; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_777 = 7'h7f == index ? _GEN_7706 : tag_0_127; // @[i_cache.scala 19:24 88:{30,30}]
  wire  _GEN_7710 = 7'h0 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_778 = 7'h0 == index | valid_0_0; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7712 = 7'h1 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_779 = 7'h1 == index | valid_0_1; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7714 = 7'h2 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_780 = 7'h2 == index | valid_0_2; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7718 = 7'h3 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_781 = 7'h3 == index | valid_0_3; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7727 = 7'h4 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_782 = 7'h4 == index | valid_0_4; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7729 = 7'h5 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_783 = 7'h5 == index | valid_0_5; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7731 = 7'h6 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_784 = 7'h6 == index | valid_0_6; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7733 = 7'h7 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_785 = 7'h7 == index | valid_0_7; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7738 = 7'h8 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_786 = 7'h8 == index | valid_0_8; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7739 = 7'h9 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_787 = 7'h9 == index | valid_0_9; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7740 = 7'ha == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_788 = 7'ha == index | valid_0_10; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7741 = 7'hb == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_789 = 7'hb == index | valid_0_11; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7742 = 7'hc == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_790 = 7'hc == index | valid_0_12; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7743 = 7'hd == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_791 = 7'hd == index | valid_0_13; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7744 = 7'he == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_792 = 7'he == index | valid_0_14; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7745 = 7'hf == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_793 = 7'hf == index | valid_0_15; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7746 = 7'h10 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_794 = 7'h10 == index | valid_0_16; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7747 = 7'h11 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_795 = 7'h11 == index | valid_0_17; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7748 = 7'h12 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_796 = 7'h12 == index | valid_0_18; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7749 = 7'h13 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_797 = 7'h13 == index | valid_0_19; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7750 = 7'h14 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_798 = 7'h14 == index | valid_0_20; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7751 = 7'h15 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_799 = 7'h15 == index | valid_0_21; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7752 = 7'h16 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_800 = 7'h16 == index | valid_0_22; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7753 = 7'h17 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_801 = 7'h17 == index | valid_0_23; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7754 = 7'h18 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_802 = 7'h18 == index | valid_0_24; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7755 = 7'h19 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_803 = 7'h19 == index | valid_0_25; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7756 = 7'h1a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_804 = 7'h1a == index | valid_0_26; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7757 = 7'h1b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_805 = 7'h1b == index | valid_0_27; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7758 = 7'h1c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_806 = 7'h1c == index | valid_0_28; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7759 = 7'h1d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_807 = 7'h1d == index | valid_0_29; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7760 = 7'h1e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_808 = 7'h1e == index | valid_0_30; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7761 = 7'h1f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_809 = 7'h1f == index | valid_0_31; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7762 = 7'h20 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_810 = 7'h20 == index | valid_0_32; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7763 = 7'h21 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_811 = 7'h21 == index | valid_0_33; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7764 = 7'h22 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_812 = 7'h22 == index | valid_0_34; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7765 = 7'h23 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_813 = 7'h23 == index | valid_0_35; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7766 = 7'h24 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_814 = 7'h24 == index | valid_0_36; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7767 = 7'h25 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_815 = 7'h25 == index | valid_0_37; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7768 = 7'h26 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_816 = 7'h26 == index | valid_0_38; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7769 = 7'h27 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_817 = 7'h27 == index | valid_0_39; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7770 = 7'h28 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_818 = 7'h28 == index | valid_0_40; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7771 = 7'h29 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_819 = 7'h29 == index | valid_0_41; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7772 = 7'h2a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_820 = 7'h2a == index | valid_0_42; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7773 = 7'h2b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_821 = 7'h2b == index | valid_0_43; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7774 = 7'h2c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_822 = 7'h2c == index | valid_0_44; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7775 = 7'h2d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_823 = 7'h2d == index | valid_0_45; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7776 = 7'h2e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_824 = 7'h2e == index | valid_0_46; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7777 = 7'h2f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_825 = 7'h2f == index | valid_0_47; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7778 = 7'h30 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_826 = 7'h30 == index | valid_0_48; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7779 = 7'h31 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_827 = 7'h31 == index | valid_0_49; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7780 = 7'h32 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_828 = 7'h32 == index | valid_0_50; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7781 = 7'h33 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_829 = 7'h33 == index | valid_0_51; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7782 = 7'h34 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_830 = 7'h34 == index | valid_0_52; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7783 = 7'h35 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_831 = 7'h35 == index | valid_0_53; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7784 = 7'h36 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_832 = 7'h36 == index | valid_0_54; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7785 = 7'h37 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_833 = 7'h37 == index | valid_0_55; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7786 = 7'h38 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_834 = 7'h38 == index | valid_0_56; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7787 = 7'h39 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_835 = 7'h39 == index | valid_0_57; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7788 = 7'h3a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_836 = 7'h3a == index | valid_0_58; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7789 = 7'h3b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_837 = 7'h3b == index | valid_0_59; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7790 = 7'h3c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_838 = 7'h3c == index | valid_0_60; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7791 = 7'h3d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_839 = 7'h3d == index | valid_0_61; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7792 = 7'h3e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_840 = 7'h3e == index | valid_0_62; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7793 = 7'h3f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_841 = 7'h3f == index | valid_0_63; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7794 = 7'h40 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_842 = 7'h40 == index | valid_0_64; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7795 = 7'h41 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_843 = 7'h41 == index | valid_0_65; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7796 = 7'h42 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_844 = 7'h42 == index | valid_0_66; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7797 = 7'h43 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_845 = 7'h43 == index | valid_0_67; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7798 = 7'h44 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_846 = 7'h44 == index | valid_0_68; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7799 = 7'h45 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_847 = 7'h45 == index | valid_0_69; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7800 = 7'h46 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_848 = 7'h46 == index | valid_0_70; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7801 = 7'h47 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_849 = 7'h47 == index | valid_0_71; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7802 = 7'h48 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_850 = 7'h48 == index | valid_0_72; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7803 = 7'h49 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_851 = 7'h49 == index | valid_0_73; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7804 = 7'h4a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_852 = 7'h4a == index | valid_0_74; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7805 = 7'h4b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_853 = 7'h4b == index | valid_0_75; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7806 = 7'h4c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_854 = 7'h4c == index | valid_0_76; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7807 = 7'h4d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_855 = 7'h4d == index | valid_0_77; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7808 = 7'h4e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_856 = 7'h4e == index | valid_0_78; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7809 = 7'h4f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_857 = 7'h4f == index | valid_0_79; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7810 = 7'h50 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_858 = 7'h50 == index | valid_0_80; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7811 = 7'h51 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_859 = 7'h51 == index | valid_0_81; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7812 = 7'h52 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_860 = 7'h52 == index | valid_0_82; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7813 = 7'h53 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_861 = 7'h53 == index | valid_0_83; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7814 = 7'h54 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_862 = 7'h54 == index | valid_0_84; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7815 = 7'h55 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_863 = 7'h55 == index | valid_0_85; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7816 = 7'h56 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_864 = 7'h56 == index | valid_0_86; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7817 = 7'h57 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_865 = 7'h57 == index | valid_0_87; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7818 = 7'h58 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_866 = 7'h58 == index | valid_0_88; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7819 = 7'h59 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_867 = 7'h59 == index | valid_0_89; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7820 = 7'h5a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_868 = 7'h5a == index | valid_0_90; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7821 = 7'h5b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_869 = 7'h5b == index | valid_0_91; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7822 = 7'h5c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_870 = 7'h5c == index | valid_0_92; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7823 = 7'h5d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_871 = 7'h5d == index | valid_0_93; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7824 = 7'h5e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_872 = 7'h5e == index | valid_0_94; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7825 = 7'h5f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_873 = 7'h5f == index | valid_0_95; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7826 = 7'h60 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_874 = 7'h60 == index | valid_0_96; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7827 = 7'h61 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_875 = 7'h61 == index | valid_0_97; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7828 = 7'h62 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_876 = 7'h62 == index | valid_0_98; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7829 = 7'h63 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_877 = 7'h63 == index | valid_0_99; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7830 = 7'h64 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_878 = 7'h64 == index | valid_0_100; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7831 = 7'h65 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_879 = 7'h65 == index | valid_0_101; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7832 = 7'h66 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_880 = 7'h66 == index | valid_0_102; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7833 = 7'h67 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_881 = 7'h67 == index | valid_0_103; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7834 = 7'h68 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_882 = 7'h68 == index | valid_0_104; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7835 = 7'h69 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_883 = 7'h69 == index | valid_0_105; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7836 = 7'h6a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_884 = 7'h6a == index | valid_0_106; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7837 = 7'h6b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_885 = 7'h6b == index | valid_0_107; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7838 = 7'h6c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_886 = 7'h6c == index | valid_0_108; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7839 = 7'h6d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_887 = 7'h6d == index | valid_0_109; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7840 = 7'h6e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_888 = 7'h6e == index | valid_0_110; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7841 = 7'h6f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_889 = 7'h6f == index | valid_0_111; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7842 = 7'h70 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_890 = 7'h70 == index | valid_0_112; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7843 = 7'h71 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_891 = 7'h71 == index | valid_0_113; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7844 = 7'h72 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_892 = 7'h72 == index | valid_0_114; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7845 = 7'h73 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_893 = 7'h73 == index | valid_0_115; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7846 = 7'h74 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_894 = 7'h74 == index | valid_0_116; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7847 = 7'h75 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_895 = 7'h75 == index | valid_0_117; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7848 = 7'h76 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_896 = 7'h76 == index | valid_0_118; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7849 = 7'h77 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_897 = 7'h77 == index | valid_0_119; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7850 = 7'h78 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_898 = 7'h78 == index | valid_0_120; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7851 = 7'h79 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_899 = 7'h79 == index | valid_0_121; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7852 = 7'h7a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_900 = 7'h7a == index | valid_0_122; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7853 = 7'h7b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_901 = 7'h7b == index | valid_0_123; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7854 = 7'h7c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_902 = 7'h7c == index | valid_0_124; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7855 = 7'h7d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_903 = 7'h7d == index | valid_0_125; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7856 = 7'h7e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_904 = 7'h7e == index | valid_0_126; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7857 = 7'h7f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_905 = 7'h7f == index | valid_0_127; // @[i_cache.scala 21:26 89:{32,32}]
  wire [63:0] _GEN_906 = 7'h0 == index ? receive_data : ram_1_0; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_907 = 7'h1 == index ? receive_data : ram_1_1; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_908 = 7'h2 == index ? receive_data : ram_1_2; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_909 = 7'h3 == index ? receive_data : ram_1_3; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_910 = 7'h4 == index ? receive_data : ram_1_4; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_911 = 7'h5 == index ? receive_data : ram_1_5; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_912 = 7'h6 == index ? receive_data : ram_1_6; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_913 = 7'h7 == index ? receive_data : ram_1_7; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_914 = 7'h8 == index ? receive_data : ram_1_8; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_915 = 7'h9 == index ? receive_data : ram_1_9; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_916 = 7'ha == index ? receive_data : ram_1_10; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_917 = 7'hb == index ? receive_data : ram_1_11; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_918 = 7'hc == index ? receive_data : ram_1_12; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_919 = 7'hd == index ? receive_data : ram_1_13; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_920 = 7'he == index ? receive_data : ram_1_14; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_921 = 7'hf == index ? receive_data : ram_1_15; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_922 = 7'h10 == index ? receive_data : ram_1_16; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_923 = 7'h11 == index ? receive_data : ram_1_17; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_924 = 7'h12 == index ? receive_data : ram_1_18; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_925 = 7'h13 == index ? receive_data : ram_1_19; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_926 = 7'h14 == index ? receive_data : ram_1_20; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_927 = 7'h15 == index ? receive_data : ram_1_21; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_928 = 7'h16 == index ? receive_data : ram_1_22; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_929 = 7'h17 == index ? receive_data : ram_1_23; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_930 = 7'h18 == index ? receive_data : ram_1_24; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_931 = 7'h19 == index ? receive_data : ram_1_25; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_932 = 7'h1a == index ? receive_data : ram_1_26; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_933 = 7'h1b == index ? receive_data : ram_1_27; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_934 = 7'h1c == index ? receive_data : ram_1_28; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_935 = 7'h1d == index ? receive_data : ram_1_29; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_936 = 7'h1e == index ? receive_data : ram_1_30; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_937 = 7'h1f == index ? receive_data : ram_1_31; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_938 = 7'h20 == index ? receive_data : ram_1_32; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_939 = 7'h21 == index ? receive_data : ram_1_33; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_940 = 7'h22 == index ? receive_data : ram_1_34; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_941 = 7'h23 == index ? receive_data : ram_1_35; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_942 = 7'h24 == index ? receive_data : ram_1_36; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_943 = 7'h25 == index ? receive_data : ram_1_37; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_944 = 7'h26 == index ? receive_data : ram_1_38; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_945 = 7'h27 == index ? receive_data : ram_1_39; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_946 = 7'h28 == index ? receive_data : ram_1_40; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_947 = 7'h29 == index ? receive_data : ram_1_41; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_948 = 7'h2a == index ? receive_data : ram_1_42; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_949 = 7'h2b == index ? receive_data : ram_1_43; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_950 = 7'h2c == index ? receive_data : ram_1_44; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_951 = 7'h2d == index ? receive_data : ram_1_45; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_952 = 7'h2e == index ? receive_data : ram_1_46; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_953 = 7'h2f == index ? receive_data : ram_1_47; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_954 = 7'h30 == index ? receive_data : ram_1_48; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_955 = 7'h31 == index ? receive_data : ram_1_49; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_956 = 7'h32 == index ? receive_data : ram_1_50; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_957 = 7'h33 == index ? receive_data : ram_1_51; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_958 = 7'h34 == index ? receive_data : ram_1_52; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_959 = 7'h35 == index ? receive_data : ram_1_53; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_960 = 7'h36 == index ? receive_data : ram_1_54; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_961 = 7'h37 == index ? receive_data : ram_1_55; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_962 = 7'h38 == index ? receive_data : ram_1_56; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_963 = 7'h39 == index ? receive_data : ram_1_57; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_964 = 7'h3a == index ? receive_data : ram_1_58; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_965 = 7'h3b == index ? receive_data : ram_1_59; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_966 = 7'h3c == index ? receive_data : ram_1_60; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_967 = 7'h3d == index ? receive_data : ram_1_61; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_968 = 7'h3e == index ? receive_data : ram_1_62; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_969 = 7'h3f == index ? receive_data : ram_1_63; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_970 = 7'h40 == index ? receive_data : ram_1_64; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_971 = 7'h41 == index ? receive_data : ram_1_65; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_972 = 7'h42 == index ? receive_data : ram_1_66; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_973 = 7'h43 == index ? receive_data : ram_1_67; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_974 = 7'h44 == index ? receive_data : ram_1_68; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_975 = 7'h45 == index ? receive_data : ram_1_69; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_976 = 7'h46 == index ? receive_data : ram_1_70; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_977 = 7'h47 == index ? receive_data : ram_1_71; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_978 = 7'h48 == index ? receive_data : ram_1_72; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_979 = 7'h49 == index ? receive_data : ram_1_73; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_980 = 7'h4a == index ? receive_data : ram_1_74; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_981 = 7'h4b == index ? receive_data : ram_1_75; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_982 = 7'h4c == index ? receive_data : ram_1_76; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_983 = 7'h4d == index ? receive_data : ram_1_77; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_984 = 7'h4e == index ? receive_data : ram_1_78; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_985 = 7'h4f == index ? receive_data : ram_1_79; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_986 = 7'h50 == index ? receive_data : ram_1_80; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_987 = 7'h51 == index ? receive_data : ram_1_81; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_988 = 7'h52 == index ? receive_data : ram_1_82; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_989 = 7'h53 == index ? receive_data : ram_1_83; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_990 = 7'h54 == index ? receive_data : ram_1_84; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_991 = 7'h55 == index ? receive_data : ram_1_85; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_992 = 7'h56 == index ? receive_data : ram_1_86; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_993 = 7'h57 == index ? receive_data : ram_1_87; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_994 = 7'h58 == index ? receive_data : ram_1_88; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_995 = 7'h59 == index ? receive_data : ram_1_89; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_996 = 7'h5a == index ? receive_data : ram_1_90; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_997 = 7'h5b == index ? receive_data : ram_1_91; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_998 = 7'h5c == index ? receive_data : ram_1_92; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_999 = 7'h5d == index ? receive_data : ram_1_93; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1000 = 7'h5e == index ? receive_data : ram_1_94; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1001 = 7'h5f == index ? receive_data : ram_1_95; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1002 = 7'h60 == index ? receive_data : ram_1_96; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1003 = 7'h61 == index ? receive_data : ram_1_97; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1004 = 7'h62 == index ? receive_data : ram_1_98; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1005 = 7'h63 == index ? receive_data : ram_1_99; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1006 = 7'h64 == index ? receive_data : ram_1_100; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1007 = 7'h65 == index ? receive_data : ram_1_101; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1008 = 7'h66 == index ? receive_data : ram_1_102; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1009 = 7'h67 == index ? receive_data : ram_1_103; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1010 = 7'h68 == index ? receive_data : ram_1_104; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1011 = 7'h69 == index ? receive_data : ram_1_105; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1012 = 7'h6a == index ? receive_data : ram_1_106; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1013 = 7'h6b == index ? receive_data : ram_1_107; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1014 = 7'h6c == index ? receive_data : ram_1_108; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1015 = 7'h6d == index ? receive_data : ram_1_109; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1016 = 7'h6e == index ? receive_data : ram_1_110; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1017 = 7'h6f == index ? receive_data : ram_1_111; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1018 = 7'h70 == index ? receive_data : ram_1_112; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1019 = 7'h71 == index ? receive_data : ram_1_113; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1020 = 7'h72 == index ? receive_data : ram_1_114; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1021 = 7'h73 == index ? receive_data : ram_1_115; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1022 = 7'h74 == index ? receive_data : ram_1_116; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1023 = 7'h75 == index ? receive_data : ram_1_117; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1024 = 7'h76 == index ? receive_data : ram_1_118; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1025 = 7'h77 == index ? receive_data : ram_1_119; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1026 = 7'h78 == index ? receive_data : ram_1_120; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1027 = 7'h79 == index ? receive_data : ram_1_121; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1028 = 7'h7a == index ? receive_data : ram_1_122; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1029 = 7'h7b == index ? receive_data : ram_1_123; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1030 = 7'h7c == index ? receive_data : ram_1_124; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1031 = 7'h7d == index ? receive_data : ram_1_125; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1032 = 7'h7e == index ? receive_data : ram_1_126; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1033 = 7'h7f == index ? receive_data : ram_1_127; // @[i_cache.scala 18:24 92:{30,30}]
  wire [31:0] _GEN_1034 = 7'h0 == index ? _GEN_7706 : tag_1_0; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1035 = 7'h1 == index ? _GEN_7706 : tag_1_1; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1036 = 7'h2 == index ? _GEN_7706 : tag_1_2; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1037 = 7'h3 == index ? _GEN_7706 : tag_1_3; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1038 = 7'h4 == index ? _GEN_7706 : tag_1_4; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1039 = 7'h5 == index ? _GEN_7706 : tag_1_5; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1040 = 7'h6 == index ? _GEN_7706 : tag_1_6; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1041 = 7'h7 == index ? _GEN_7706 : tag_1_7; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1042 = 7'h8 == index ? _GEN_7706 : tag_1_8; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1043 = 7'h9 == index ? _GEN_7706 : tag_1_9; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1044 = 7'ha == index ? _GEN_7706 : tag_1_10; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1045 = 7'hb == index ? _GEN_7706 : tag_1_11; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1046 = 7'hc == index ? _GEN_7706 : tag_1_12; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1047 = 7'hd == index ? _GEN_7706 : tag_1_13; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1048 = 7'he == index ? _GEN_7706 : tag_1_14; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1049 = 7'hf == index ? _GEN_7706 : tag_1_15; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1050 = 7'h10 == index ? _GEN_7706 : tag_1_16; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1051 = 7'h11 == index ? _GEN_7706 : tag_1_17; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1052 = 7'h12 == index ? _GEN_7706 : tag_1_18; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1053 = 7'h13 == index ? _GEN_7706 : tag_1_19; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1054 = 7'h14 == index ? _GEN_7706 : tag_1_20; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1055 = 7'h15 == index ? _GEN_7706 : tag_1_21; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1056 = 7'h16 == index ? _GEN_7706 : tag_1_22; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1057 = 7'h17 == index ? _GEN_7706 : tag_1_23; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1058 = 7'h18 == index ? _GEN_7706 : tag_1_24; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1059 = 7'h19 == index ? _GEN_7706 : tag_1_25; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1060 = 7'h1a == index ? _GEN_7706 : tag_1_26; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1061 = 7'h1b == index ? _GEN_7706 : tag_1_27; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1062 = 7'h1c == index ? _GEN_7706 : tag_1_28; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1063 = 7'h1d == index ? _GEN_7706 : tag_1_29; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1064 = 7'h1e == index ? _GEN_7706 : tag_1_30; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1065 = 7'h1f == index ? _GEN_7706 : tag_1_31; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1066 = 7'h20 == index ? _GEN_7706 : tag_1_32; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1067 = 7'h21 == index ? _GEN_7706 : tag_1_33; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1068 = 7'h22 == index ? _GEN_7706 : tag_1_34; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1069 = 7'h23 == index ? _GEN_7706 : tag_1_35; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1070 = 7'h24 == index ? _GEN_7706 : tag_1_36; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1071 = 7'h25 == index ? _GEN_7706 : tag_1_37; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1072 = 7'h26 == index ? _GEN_7706 : tag_1_38; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1073 = 7'h27 == index ? _GEN_7706 : tag_1_39; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1074 = 7'h28 == index ? _GEN_7706 : tag_1_40; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1075 = 7'h29 == index ? _GEN_7706 : tag_1_41; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1076 = 7'h2a == index ? _GEN_7706 : tag_1_42; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1077 = 7'h2b == index ? _GEN_7706 : tag_1_43; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1078 = 7'h2c == index ? _GEN_7706 : tag_1_44; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1079 = 7'h2d == index ? _GEN_7706 : tag_1_45; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1080 = 7'h2e == index ? _GEN_7706 : tag_1_46; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1081 = 7'h2f == index ? _GEN_7706 : tag_1_47; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1082 = 7'h30 == index ? _GEN_7706 : tag_1_48; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1083 = 7'h31 == index ? _GEN_7706 : tag_1_49; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1084 = 7'h32 == index ? _GEN_7706 : tag_1_50; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1085 = 7'h33 == index ? _GEN_7706 : tag_1_51; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1086 = 7'h34 == index ? _GEN_7706 : tag_1_52; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1087 = 7'h35 == index ? _GEN_7706 : tag_1_53; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1088 = 7'h36 == index ? _GEN_7706 : tag_1_54; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1089 = 7'h37 == index ? _GEN_7706 : tag_1_55; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1090 = 7'h38 == index ? _GEN_7706 : tag_1_56; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1091 = 7'h39 == index ? _GEN_7706 : tag_1_57; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1092 = 7'h3a == index ? _GEN_7706 : tag_1_58; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1093 = 7'h3b == index ? _GEN_7706 : tag_1_59; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1094 = 7'h3c == index ? _GEN_7706 : tag_1_60; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1095 = 7'h3d == index ? _GEN_7706 : tag_1_61; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1096 = 7'h3e == index ? _GEN_7706 : tag_1_62; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1097 = 7'h3f == index ? _GEN_7706 : tag_1_63; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1098 = 7'h40 == index ? _GEN_7706 : tag_1_64; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1099 = 7'h41 == index ? _GEN_7706 : tag_1_65; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1100 = 7'h42 == index ? _GEN_7706 : tag_1_66; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1101 = 7'h43 == index ? _GEN_7706 : tag_1_67; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1102 = 7'h44 == index ? _GEN_7706 : tag_1_68; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1103 = 7'h45 == index ? _GEN_7706 : tag_1_69; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1104 = 7'h46 == index ? _GEN_7706 : tag_1_70; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1105 = 7'h47 == index ? _GEN_7706 : tag_1_71; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1106 = 7'h48 == index ? _GEN_7706 : tag_1_72; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1107 = 7'h49 == index ? _GEN_7706 : tag_1_73; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1108 = 7'h4a == index ? _GEN_7706 : tag_1_74; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1109 = 7'h4b == index ? _GEN_7706 : tag_1_75; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1110 = 7'h4c == index ? _GEN_7706 : tag_1_76; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1111 = 7'h4d == index ? _GEN_7706 : tag_1_77; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1112 = 7'h4e == index ? _GEN_7706 : tag_1_78; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1113 = 7'h4f == index ? _GEN_7706 : tag_1_79; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1114 = 7'h50 == index ? _GEN_7706 : tag_1_80; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1115 = 7'h51 == index ? _GEN_7706 : tag_1_81; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1116 = 7'h52 == index ? _GEN_7706 : tag_1_82; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1117 = 7'h53 == index ? _GEN_7706 : tag_1_83; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1118 = 7'h54 == index ? _GEN_7706 : tag_1_84; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1119 = 7'h55 == index ? _GEN_7706 : tag_1_85; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1120 = 7'h56 == index ? _GEN_7706 : tag_1_86; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1121 = 7'h57 == index ? _GEN_7706 : tag_1_87; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1122 = 7'h58 == index ? _GEN_7706 : tag_1_88; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1123 = 7'h59 == index ? _GEN_7706 : tag_1_89; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1124 = 7'h5a == index ? _GEN_7706 : tag_1_90; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1125 = 7'h5b == index ? _GEN_7706 : tag_1_91; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1126 = 7'h5c == index ? _GEN_7706 : tag_1_92; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1127 = 7'h5d == index ? _GEN_7706 : tag_1_93; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1128 = 7'h5e == index ? _GEN_7706 : tag_1_94; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1129 = 7'h5f == index ? _GEN_7706 : tag_1_95; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1130 = 7'h60 == index ? _GEN_7706 : tag_1_96; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1131 = 7'h61 == index ? _GEN_7706 : tag_1_97; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1132 = 7'h62 == index ? _GEN_7706 : tag_1_98; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1133 = 7'h63 == index ? _GEN_7706 : tag_1_99; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1134 = 7'h64 == index ? _GEN_7706 : tag_1_100; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1135 = 7'h65 == index ? _GEN_7706 : tag_1_101; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1136 = 7'h66 == index ? _GEN_7706 : tag_1_102; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1137 = 7'h67 == index ? _GEN_7706 : tag_1_103; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1138 = 7'h68 == index ? _GEN_7706 : tag_1_104; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1139 = 7'h69 == index ? _GEN_7706 : tag_1_105; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1140 = 7'h6a == index ? _GEN_7706 : tag_1_106; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1141 = 7'h6b == index ? _GEN_7706 : tag_1_107; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1142 = 7'h6c == index ? _GEN_7706 : tag_1_108; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1143 = 7'h6d == index ? _GEN_7706 : tag_1_109; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1144 = 7'h6e == index ? _GEN_7706 : tag_1_110; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1145 = 7'h6f == index ? _GEN_7706 : tag_1_111; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1146 = 7'h70 == index ? _GEN_7706 : tag_1_112; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1147 = 7'h71 == index ? _GEN_7706 : tag_1_113; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1148 = 7'h72 == index ? _GEN_7706 : tag_1_114; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1149 = 7'h73 == index ? _GEN_7706 : tag_1_115; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1150 = 7'h74 == index ? _GEN_7706 : tag_1_116; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1151 = 7'h75 == index ? _GEN_7706 : tag_1_117; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1152 = 7'h76 == index ? _GEN_7706 : tag_1_118; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1153 = 7'h77 == index ? _GEN_7706 : tag_1_119; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1154 = 7'h78 == index ? _GEN_7706 : tag_1_120; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1155 = 7'h79 == index ? _GEN_7706 : tag_1_121; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1156 = 7'h7a == index ? _GEN_7706 : tag_1_122; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1157 = 7'h7b == index ? _GEN_7706 : tag_1_123; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1158 = 7'h7c == index ? _GEN_7706 : tag_1_124; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1159 = 7'h7d == index ? _GEN_7706 : tag_1_125; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1160 = 7'h7e == index ? _GEN_7706 : tag_1_126; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1161 = 7'h7f == index ? _GEN_7706 : tag_1_127; // @[i_cache.scala 20:24 93:{30,30}]
  wire  _GEN_1162 = _GEN_7710 | valid_1_0; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1163 = _GEN_7712 | valid_1_1; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1164 = _GEN_7714 | valid_1_2; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1165 = _GEN_7718 | valid_1_3; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1166 = _GEN_7727 | valid_1_4; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1167 = _GEN_7729 | valid_1_5; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1168 = _GEN_7731 | valid_1_6; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1169 = _GEN_7733 | valid_1_7; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1170 = _GEN_7738 | valid_1_8; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1171 = _GEN_7739 | valid_1_9; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1172 = _GEN_7740 | valid_1_10; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1173 = _GEN_7741 | valid_1_11; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1174 = _GEN_7742 | valid_1_12; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1175 = _GEN_7743 | valid_1_13; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1176 = _GEN_7744 | valid_1_14; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1177 = _GEN_7745 | valid_1_15; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1178 = _GEN_7746 | valid_1_16; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1179 = _GEN_7747 | valid_1_17; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1180 = _GEN_7748 | valid_1_18; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1181 = _GEN_7749 | valid_1_19; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1182 = _GEN_7750 | valid_1_20; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1183 = _GEN_7751 | valid_1_21; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1184 = _GEN_7752 | valid_1_22; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1185 = _GEN_7753 | valid_1_23; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1186 = _GEN_7754 | valid_1_24; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1187 = _GEN_7755 | valid_1_25; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1188 = _GEN_7756 | valid_1_26; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1189 = _GEN_7757 | valid_1_27; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1190 = _GEN_7758 | valid_1_28; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1191 = _GEN_7759 | valid_1_29; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1192 = _GEN_7760 | valid_1_30; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1193 = _GEN_7761 | valid_1_31; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1194 = _GEN_7762 | valid_1_32; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1195 = _GEN_7763 | valid_1_33; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1196 = _GEN_7764 | valid_1_34; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1197 = _GEN_7765 | valid_1_35; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1198 = _GEN_7766 | valid_1_36; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1199 = _GEN_7767 | valid_1_37; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1200 = _GEN_7768 | valid_1_38; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1201 = _GEN_7769 | valid_1_39; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1202 = _GEN_7770 | valid_1_40; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1203 = _GEN_7771 | valid_1_41; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1204 = _GEN_7772 | valid_1_42; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1205 = _GEN_7773 | valid_1_43; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1206 = _GEN_7774 | valid_1_44; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1207 = _GEN_7775 | valid_1_45; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1208 = _GEN_7776 | valid_1_46; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1209 = _GEN_7777 | valid_1_47; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1210 = _GEN_7778 | valid_1_48; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1211 = _GEN_7779 | valid_1_49; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1212 = _GEN_7780 | valid_1_50; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1213 = _GEN_7781 | valid_1_51; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1214 = _GEN_7782 | valid_1_52; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1215 = _GEN_7783 | valid_1_53; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1216 = _GEN_7784 | valid_1_54; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1217 = _GEN_7785 | valid_1_55; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1218 = _GEN_7786 | valid_1_56; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1219 = _GEN_7787 | valid_1_57; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1220 = _GEN_7788 | valid_1_58; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1221 = _GEN_7789 | valid_1_59; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1222 = _GEN_7790 | valid_1_60; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1223 = _GEN_7791 | valid_1_61; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1224 = _GEN_7792 | valid_1_62; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1225 = _GEN_7793 | valid_1_63; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1226 = _GEN_7794 | valid_1_64; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1227 = _GEN_7795 | valid_1_65; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1228 = _GEN_7796 | valid_1_66; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1229 = _GEN_7797 | valid_1_67; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1230 = _GEN_7798 | valid_1_68; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1231 = _GEN_7799 | valid_1_69; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1232 = _GEN_7800 | valid_1_70; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1233 = _GEN_7801 | valid_1_71; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1234 = _GEN_7802 | valid_1_72; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1235 = _GEN_7803 | valid_1_73; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1236 = _GEN_7804 | valid_1_74; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1237 = _GEN_7805 | valid_1_75; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1238 = _GEN_7806 | valid_1_76; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1239 = _GEN_7807 | valid_1_77; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1240 = _GEN_7808 | valid_1_78; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1241 = _GEN_7809 | valid_1_79; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1242 = _GEN_7810 | valid_1_80; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1243 = _GEN_7811 | valid_1_81; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1244 = _GEN_7812 | valid_1_82; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1245 = _GEN_7813 | valid_1_83; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1246 = _GEN_7814 | valid_1_84; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1247 = _GEN_7815 | valid_1_85; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1248 = _GEN_7816 | valid_1_86; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1249 = _GEN_7817 | valid_1_87; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1250 = _GEN_7818 | valid_1_88; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1251 = _GEN_7819 | valid_1_89; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1252 = _GEN_7820 | valid_1_90; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1253 = _GEN_7821 | valid_1_91; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1254 = _GEN_7822 | valid_1_92; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1255 = _GEN_7823 | valid_1_93; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1256 = _GEN_7824 | valid_1_94; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1257 = _GEN_7825 | valid_1_95; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1258 = _GEN_7826 | valid_1_96; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1259 = _GEN_7827 | valid_1_97; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1260 = _GEN_7828 | valid_1_98; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1261 = _GEN_7829 | valid_1_99; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1262 = _GEN_7830 | valid_1_100; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1263 = _GEN_7831 | valid_1_101; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1264 = _GEN_7832 | valid_1_102; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1265 = _GEN_7833 | valid_1_103; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1266 = _GEN_7834 | valid_1_104; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1267 = _GEN_7835 | valid_1_105; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1268 = _GEN_7836 | valid_1_106; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1269 = _GEN_7837 | valid_1_107; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1270 = _GEN_7838 | valid_1_108; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1271 = _GEN_7839 | valid_1_109; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1272 = _GEN_7840 | valid_1_110; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1273 = _GEN_7841 | valid_1_111; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1274 = _GEN_7842 | valid_1_112; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1275 = _GEN_7843 | valid_1_113; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1276 = _GEN_7844 | valid_1_114; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1277 = _GEN_7845 | valid_1_115; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1278 = _GEN_7846 | valid_1_116; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1279 = _GEN_7847 | valid_1_117; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1280 = _GEN_7848 | valid_1_118; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1281 = _GEN_7849 | valid_1_119; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1282 = _GEN_7850 | valid_1_120; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1283 = _GEN_7851 | valid_1_121; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1284 = _GEN_7852 | valid_1_122; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1285 = _GEN_7853 | valid_1_123; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1286 = _GEN_7854 | valid_1_124; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1287 = _GEN_7855 | valid_1_125; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1288 = _GEN_7856 | valid_1_126; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1289 = _GEN_7857 | valid_1_127; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _T_14 = ~quene; // @[i_cache.scala 97:27]
  wire [63:0] _GEN_2058 = ~quene ? _GEN_522 : ram_0_0; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2059 = ~quene ? _GEN_523 : ram_0_1; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2060 = ~quene ? _GEN_524 : ram_0_2; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2061 = ~quene ? _GEN_525 : ram_0_3; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2062 = ~quene ? _GEN_526 : ram_0_4; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2063 = ~quene ? _GEN_527 : ram_0_5; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2064 = ~quene ? _GEN_528 : ram_0_6; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2065 = ~quene ? _GEN_529 : ram_0_7; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2066 = ~quene ? _GEN_530 : ram_0_8; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2067 = ~quene ? _GEN_531 : ram_0_9; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2068 = ~quene ? _GEN_532 : ram_0_10; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2069 = ~quene ? _GEN_533 : ram_0_11; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2070 = ~quene ? _GEN_534 : ram_0_12; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2071 = ~quene ? _GEN_535 : ram_0_13; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2072 = ~quene ? _GEN_536 : ram_0_14; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2073 = ~quene ? _GEN_537 : ram_0_15; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2074 = ~quene ? _GEN_538 : ram_0_16; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2075 = ~quene ? _GEN_539 : ram_0_17; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2076 = ~quene ? _GEN_540 : ram_0_18; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2077 = ~quene ? _GEN_541 : ram_0_19; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2078 = ~quene ? _GEN_542 : ram_0_20; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2079 = ~quene ? _GEN_543 : ram_0_21; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2080 = ~quene ? _GEN_544 : ram_0_22; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2081 = ~quene ? _GEN_545 : ram_0_23; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2082 = ~quene ? _GEN_546 : ram_0_24; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2083 = ~quene ? _GEN_547 : ram_0_25; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2084 = ~quene ? _GEN_548 : ram_0_26; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2085 = ~quene ? _GEN_549 : ram_0_27; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2086 = ~quene ? _GEN_550 : ram_0_28; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2087 = ~quene ? _GEN_551 : ram_0_29; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2088 = ~quene ? _GEN_552 : ram_0_30; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2089 = ~quene ? _GEN_553 : ram_0_31; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2090 = ~quene ? _GEN_554 : ram_0_32; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2091 = ~quene ? _GEN_555 : ram_0_33; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2092 = ~quene ? _GEN_556 : ram_0_34; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2093 = ~quene ? _GEN_557 : ram_0_35; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2094 = ~quene ? _GEN_558 : ram_0_36; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2095 = ~quene ? _GEN_559 : ram_0_37; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2096 = ~quene ? _GEN_560 : ram_0_38; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2097 = ~quene ? _GEN_561 : ram_0_39; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2098 = ~quene ? _GEN_562 : ram_0_40; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2099 = ~quene ? _GEN_563 : ram_0_41; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2100 = ~quene ? _GEN_564 : ram_0_42; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2101 = ~quene ? _GEN_565 : ram_0_43; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2102 = ~quene ? _GEN_566 : ram_0_44; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2103 = ~quene ? _GEN_567 : ram_0_45; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2104 = ~quene ? _GEN_568 : ram_0_46; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2105 = ~quene ? _GEN_569 : ram_0_47; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2106 = ~quene ? _GEN_570 : ram_0_48; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2107 = ~quene ? _GEN_571 : ram_0_49; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2108 = ~quene ? _GEN_572 : ram_0_50; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2109 = ~quene ? _GEN_573 : ram_0_51; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2110 = ~quene ? _GEN_574 : ram_0_52; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2111 = ~quene ? _GEN_575 : ram_0_53; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2112 = ~quene ? _GEN_576 : ram_0_54; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2113 = ~quene ? _GEN_577 : ram_0_55; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2114 = ~quene ? _GEN_578 : ram_0_56; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2115 = ~quene ? _GEN_579 : ram_0_57; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2116 = ~quene ? _GEN_580 : ram_0_58; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2117 = ~quene ? _GEN_581 : ram_0_59; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2118 = ~quene ? _GEN_582 : ram_0_60; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2119 = ~quene ? _GEN_583 : ram_0_61; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2120 = ~quene ? _GEN_584 : ram_0_62; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2121 = ~quene ? _GEN_585 : ram_0_63; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2122 = ~quene ? _GEN_586 : ram_0_64; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2123 = ~quene ? _GEN_587 : ram_0_65; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2124 = ~quene ? _GEN_588 : ram_0_66; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2125 = ~quene ? _GEN_589 : ram_0_67; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2126 = ~quene ? _GEN_590 : ram_0_68; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2127 = ~quene ? _GEN_591 : ram_0_69; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2128 = ~quene ? _GEN_592 : ram_0_70; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2129 = ~quene ? _GEN_593 : ram_0_71; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2130 = ~quene ? _GEN_594 : ram_0_72; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2131 = ~quene ? _GEN_595 : ram_0_73; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2132 = ~quene ? _GEN_596 : ram_0_74; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2133 = ~quene ? _GEN_597 : ram_0_75; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2134 = ~quene ? _GEN_598 : ram_0_76; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2135 = ~quene ? _GEN_599 : ram_0_77; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2136 = ~quene ? _GEN_600 : ram_0_78; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2137 = ~quene ? _GEN_601 : ram_0_79; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2138 = ~quene ? _GEN_602 : ram_0_80; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2139 = ~quene ? _GEN_603 : ram_0_81; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2140 = ~quene ? _GEN_604 : ram_0_82; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2141 = ~quene ? _GEN_605 : ram_0_83; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2142 = ~quene ? _GEN_606 : ram_0_84; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2143 = ~quene ? _GEN_607 : ram_0_85; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2144 = ~quene ? _GEN_608 : ram_0_86; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2145 = ~quene ? _GEN_609 : ram_0_87; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2146 = ~quene ? _GEN_610 : ram_0_88; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2147 = ~quene ? _GEN_611 : ram_0_89; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2148 = ~quene ? _GEN_612 : ram_0_90; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2149 = ~quene ? _GEN_613 : ram_0_91; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2150 = ~quene ? _GEN_614 : ram_0_92; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2151 = ~quene ? _GEN_615 : ram_0_93; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2152 = ~quene ? _GEN_616 : ram_0_94; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2153 = ~quene ? _GEN_617 : ram_0_95; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2154 = ~quene ? _GEN_618 : ram_0_96; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2155 = ~quene ? _GEN_619 : ram_0_97; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2156 = ~quene ? _GEN_620 : ram_0_98; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2157 = ~quene ? _GEN_621 : ram_0_99; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2158 = ~quene ? _GEN_622 : ram_0_100; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2159 = ~quene ? _GEN_623 : ram_0_101; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2160 = ~quene ? _GEN_624 : ram_0_102; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2161 = ~quene ? _GEN_625 : ram_0_103; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2162 = ~quene ? _GEN_626 : ram_0_104; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2163 = ~quene ? _GEN_627 : ram_0_105; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2164 = ~quene ? _GEN_628 : ram_0_106; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2165 = ~quene ? _GEN_629 : ram_0_107; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2166 = ~quene ? _GEN_630 : ram_0_108; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2167 = ~quene ? _GEN_631 : ram_0_109; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2168 = ~quene ? _GEN_632 : ram_0_110; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2169 = ~quene ? _GEN_633 : ram_0_111; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2170 = ~quene ? _GEN_634 : ram_0_112; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2171 = ~quene ? _GEN_635 : ram_0_113; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2172 = ~quene ? _GEN_636 : ram_0_114; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2173 = ~quene ? _GEN_637 : ram_0_115; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2174 = ~quene ? _GEN_638 : ram_0_116; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2175 = ~quene ? _GEN_639 : ram_0_117; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2176 = ~quene ? _GEN_640 : ram_0_118; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2177 = ~quene ? _GEN_641 : ram_0_119; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2178 = ~quene ? _GEN_642 : ram_0_120; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2179 = ~quene ? _GEN_643 : ram_0_121; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2180 = ~quene ? _GEN_644 : ram_0_122; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2181 = ~quene ? _GEN_645 : ram_0_123; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2182 = ~quene ? _GEN_646 : ram_0_124; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2183 = ~quene ? _GEN_647 : ram_0_125; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2184 = ~quene ? _GEN_648 : ram_0_126; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2185 = ~quene ? _GEN_649 : ram_0_127; // @[i_cache.scala 17:24 97:34]
  wire [31:0] _GEN_2186 = ~quene ? _GEN_650 : tag_0_0; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2187 = ~quene ? _GEN_651 : tag_0_1; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2188 = ~quene ? _GEN_652 : tag_0_2; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2189 = ~quene ? _GEN_653 : tag_0_3; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2190 = ~quene ? _GEN_654 : tag_0_4; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2191 = ~quene ? _GEN_655 : tag_0_5; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2192 = ~quene ? _GEN_656 : tag_0_6; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2193 = ~quene ? _GEN_657 : tag_0_7; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2194 = ~quene ? _GEN_658 : tag_0_8; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2195 = ~quene ? _GEN_659 : tag_0_9; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2196 = ~quene ? _GEN_660 : tag_0_10; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2197 = ~quene ? _GEN_661 : tag_0_11; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2198 = ~quene ? _GEN_662 : tag_0_12; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2199 = ~quene ? _GEN_663 : tag_0_13; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2200 = ~quene ? _GEN_664 : tag_0_14; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2201 = ~quene ? _GEN_665 : tag_0_15; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2202 = ~quene ? _GEN_666 : tag_0_16; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2203 = ~quene ? _GEN_667 : tag_0_17; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2204 = ~quene ? _GEN_668 : tag_0_18; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2205 = ~quene ? _GEN_669 : tag_0_19; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2206 = ~quene ? _GEN_670 : tag_0_20; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2207 = ~quene ? _GEN_671 : tag_0_21; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2208 = ~quene ? _GEN_672 : tag_0_22; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2209 = ~quene ? _GEN_673 : tag_0_23; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2210 = ~quene ? _GEN_674 : tag_0_24; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2211 = ~quene ? _GEN_675 : tag_0_25; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2212 = ~quene ? _GEN_676 : tag_0_26; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2213 = ~quene ? _GEN_677 : tag_0_27; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2214 = ~quene ? _GEN_678 : tag_0_28; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2215 = ~quene ? _GEN_679 : tag_0_29; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2216 = ~quene ? _GEN_680 : tag_0_30; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2217 = ~quene ? _GEN_681 : tag_0_31; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2218 = ~quene ? _GEN_682 : tag_0_32; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2219 = ~quene ? _GEN_683 : tag_0_33; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2220 = ~quene ? _GEN_684 : tag_0_34; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2221 = ~quene ? _GEN_685 : tag_0_35; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2222 = ~quene ? _GEN_686 : tag_0_36; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2223 = ~quene ? _GEN_687 : tag_0_37; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2224 = ~quene ? _GEN_688 : tag_0_38; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2225 = ~quene ? _GEN_689 : tag_0_39; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2226 = ~quene ? _GEN_690 : tag_0_40; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2227 = ~quene ? _GEN_691 : tag_0_41; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2228 = ~quene ? _GEN_692 : tag_0_42; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2229 = ~quene ? _GEN_693 : tag_0_43; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2230 = ~quene ? _GEN_694 : tag_0_44; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2231 = ~quene ? _GEN_695 : tag_0_45; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2232 = ~quene ? _GEN_696 : tag_0_46; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2233 = ~quene ? _GEN_697 : tag_0_47; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2234 = ~quene ? _GEN_698 : tag_0_48; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2235 = ~quene ? _GEN_699 : tag_0_49; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2236 = ~quene ? _GEN_700 : tag_0_50; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2237 = ~quene ? _GEN_701 : tag_0_51; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2238 = ~quene ? _GEN_702 : tag_0_52; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2239 = ~quene ? _GEN_703 : tag_0_53; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2240 = ~quene ? _GEN_704 : tag_0_54; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2241 = ~quene ? _GEN_705 : tag_0_55; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2242 = ~quene ? _GEN_706 : tag_0_56; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2243 = ~quene ? _GEN_707 : tag_0_57; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2244 = ~quene ? _GEN_708 : tag_0_58; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2245 = ~quene ? _GEN_709 : tag_0_59; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2246 = ~quene ? _GEN_710 : tag_0_60; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2247 = ~quene ? _GEN_711 : tag_0_61; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2248 = ~quene ? _GEN_712 : tag_0_62; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2249 = ~quene ? _GEN_713 : tag_0_63; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2250 = ~quene ? _GEN_714 : tag_0_64; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2251 = ~quene ? _GEN_715 : tag_0_65; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2252 = ~quene ? _GEN_716 : tag_0_66; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2253 = ~quene ? _GEN_717 : tag_0_67; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2254 = ~quene ? _GEN_718 : tag_0_68; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2255 = ~quene ? _GEN_719 : tag_0_69; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2256 = ~quene ? _GEN_720 : tag_0_70; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2257 = ~quene ? _GEN_721 : tag_0_71; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2258 = ~quene ? _GEN_722 : tag_0_72; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2259 = ~quene ? _GEN_723 : tag_0_73; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2260 = ~quene ? _GEN_724 : tag_0_74; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2261 = ~quene ? _GEN_725 : tag_0_75; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2262 = ~quene ? _GEN_726 : tag_0_76; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2263 = ~quene ? _GEN_727 : tag_0_77; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2264 = ~quene ? _GEN_728 : tag_0_78; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2265 = ~quene ? _GEN_729 : tag_0_79; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2266 = ~quene ? _GEN_730 : tag_0_80; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2267 = ~quene ? _GEN_731 : tag_0_81; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2268 = ~quene ? _GEN_732 : tag_0_82; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2269 = ~quene ? _GEN_733 : tag_0_83; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2270 = ~quene ? _GEN_734 : tag_0_84; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2271 = ~quene ? _GEN_735 : tag_0_85; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2272 = ~quene ? _GEN_736 : tag_0_86; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2273 = ~quene ? _GEN_737 : tag_0_87; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2274 = ~quene ? _GEN_738 : tag_0_88; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2275 = ~quene ? _GEN_739 : tag_0_89; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2276 = ~quene ? _GEN_740 : tag_0_90; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2277 = ~quene ? _GEN_741 : tag_0_91; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2278 = ~quene ? _GEN_742 : tag_0_92; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2279 = ~quene ? _GEN_743 : tag_0_93; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2280 = ~quene ? _GEN_744 : tag_0_94; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2281 = ~quene ? _GEN_745 : tag_0_95; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2282 = ~quene ? _GEN_746 : tag_0_96; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2283 = ~quene ? _GEN_747 : tag_0_97; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2284 = ~quene ? _GEN_748 : tag_0_98; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2285 = ~quene ? _GEN_749 : tag_0_99; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2286 = ~quene ? _GEN_750 : tag_0_100; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2287 = ~quene ? _GEN_751 : tag_0_101; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2288 = ~quene ? _GEN_752 : tag_0_102; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2289 = ~quene ? _GEN_753 : tag_0_103; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2290 = ~quene ? _GEN_754 : tag_0_104; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2291 = ~quene ? _GEN_755 : tag_0_105; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2292 = ~quene ? _GEN_756 : tag_0_106; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2293 = ~quene ? _GEN_757 : tag_0_107; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2294 = ~quene ? _GEN_758 : tag_0_108; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2295 = ~quene ? _GEN_759 : tag_0_109; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2296 = ~quene ? _GEN_760 : tag_0_110; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2297 = ~quene ? _GEN_761 : tag_0_111; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2298 = ~quene ? _GEN_762 : tag_0_112; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2299 = ~quene ? _GEN_763 : tag_0_113; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2300 = ~quene ? _GEN_764 : tag_0_114; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2301 = ~quene ? _GEN_765 : tag_0_115; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2302 = ~quene ? _GEN_766 : tag_0_116; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2303 = ~quene ? _GEN_767 : tag_0_117; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2304 = ~quene ? _GEN_768 : tag_0_118; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2305 = ~quene ? _GEN_769 : tag_0_119; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2306 = ~quene ? _GEN_770 : tag_0_120; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2307 = ~quene ? _GEN_771 : tag_0_121; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2308 = ~quene ? _GEN_772 : tag_0_122; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2309 = ~quene ? _GEN_773 : tag_0_123; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2310 = ~quene ? _GEN_774 : tag_0_124; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2311 = ~quene ? _GEN_775 : tag_0_125; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2312 = ~quene ? _GEN_776 : tag_0_126; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2313 = ~quene ? _GEN_777 : tag_0_127; // @[i_cache.scala 19:24 97:34]
  wire  _GEN_2314 = ~quene ? _GEN_778 : valid_0_0; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2315 = ~quene ? _GEN_779 : valid_0_1; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2316 = ~quene ? _GEN_780 : valid_0_2; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2317 = ~quene ? _GEN_781 : valid_0_3; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2318 = ~quene ? _GEN_782 : valid_0_4; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2319 = ~quene ? _GEN_783 : valid_0_5; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2320 = ~quene ? _GEN_784 : valid_0_6; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2321 = ~quene ? _GEN_785 : valid_0_7; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2322 = ~quene ? _GEN_786 : valid_0_8; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2323 = ~quene ? _GEN_787 : valid_0_9; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2324 = ~quene ? _GEN_788 : valid_0_10; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2325 = ~quene ? _GEN_789 : valid_0_11; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2326 = ~quene ? _GEN_790 : valid_0_12; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2327 = ~quene ? _GEN_791 : valid_0_13; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2328 = ~quene ? _GEN_792 : valid_0_14; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2329 = ~quene ? _GEN_793 : valid_0_15; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2330 = ~quene ? _GEN_794 : valid_0_16; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2331 = ~quene ? _GEN_795 : valid_0_17; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2332 = ~quene ? _GEN_796 : valid_0_18; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2333 = ~quene ? _GEN_797 : valid_0_19; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2334 = ~quene ? _GEN_798 : valid_0_20; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2335 = ~quene ? _GEN_799 : valid_0_21; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2336 = ~quene ? _GEN_800 : valid_0_22; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2337 = ~quene ? _GEN_801 : valid_0_23; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2338 = ~quene ? _GEN_802 : valid_0_24; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2339 = ~quene ? _GEN_803 : valid_0_25; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2340 = ~quene ? _GEN_804 : valid_0_26; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2341 = ~quene ? _GEN_805 : valid_0_27; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2342 = ~quene ? _GEN_806 : valid_0_28; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2343 = ~quene ? _GEN_807 : valid_0_29; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2344 = ~quene ? _GEN_808 : valid_0_30; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2345 = ~quene ? _GEN_809 : valid_0_31; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2346 = ~quene ? _GEN_810 : valid_0_32; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2347 = ~quene ? _GEN_811 : valid_0_33; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2348 = ~quene ? _GEN_812 : valid_0_34; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2349 = ~quene ? _GEN_813 : valid_0_35; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2350 = ~quene ? _GEN_814 : valid_0_36; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2351 = ~quene ? _GEN_815 : valid_0_37; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2352 = ~quene ? _GEN_816 : valid_0_38; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2353 = ~quene ? _GEN_817 : valid_0_39; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2354 = ~quene ? _GEN_818 : valid_0_40; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2355 = ~quene ? _GEN_819 : valid_0_41; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2356 = ~quene ? _GEN_820 : valid_0_42; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2357 = ~quene ? _GEN_821 : valid_0_43; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2358 = ~quene ? _GEN_822 : valid_0_44; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2359 = ~quene ? _GEN_823 : valid_0_45; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2360 = ~quene ? _GEN_824 : valid_0_46; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2361 = ~quene ? _GEN_825 : valid_0_47; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2362 = ~quene ? _GEN_826 : valid_0_48; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2363 = ~quene ? _GEN_827 : valid_0_49; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2364 = ~quene ? _GEN_828 : valid_0_50; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2365 = ~quene ? _GEN_829 : valid_0_51; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2366 = ~quene ? _GEN_830 : valid_0_52; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2367 = ~quene ? _GEN_831 : valid_0_53; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2368 = ~quene ? _GEN_832 : valid_0_54; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2369 = ~quene ? _GEN_833 : valid_0_55; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2370 = ~quene ? _GEN_834 : valid_0_56; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2371 = ~quene ? _GEN_835 : valid_0_57; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2372 = ~quene ? _GEN_836 : valid_0_58; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2373 = ~quene ? _GEN_837 : valid_0_59; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2374 = ~quene ? _GEN_838 : valid_0_60; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2375 = ~quene ? _GEN_839 : valid_0_61; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2376 = ~quene ? _GEN_840 : valid_0_62; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2377 = ~quene ? _GEN_841 : valid_0_63; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2378 = ~quene ? _GEN_842 : valid_0_64; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2379 = ~quene ? _GEN_843 : valid_0_65; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2380 = ~quene ? _GEN_844 : valid_0_66; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2381 = ~quene ? _GEN_845 : valid_0_67; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2382 = ~quene ? _GEN_846 : valid_0_68; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2383 = ~quene ? _GEN_847 : valid_0_69; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2384 = ~quene ? _GEN_848 : valid_0_70; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2385 = ~quene ? _GEN_849 : valid_0_71; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2386 = ~quene ? _GEN_850 : valid_0_72; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2387 = ~quene ? _GEN_851 : valid_0_73; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2388 = ~quene ? _GEN_852 : valid_0_74; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2389 = ~quene ? _GEN_853 : valid_0_75; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2390 = ~quene ? _GEN_854 : valid_0_76; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2391 = ~quene ? _GEN_855 : valid_0_77; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2392 = ~quene ? _GEN_856 : valid_0_78; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2393 = ~quene ? _GEN_857 : valid_0_79; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2394 = ~quene ? _GEN_858 : valid_0_80; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2395 = ~quene ? _GEN_859 : valid_0_81; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2396 = ~quene ? _GEN_860 : valid_0_82; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2397 = ~quene ? _GEN_861 : valid_0_83; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2398 = ~quene ? _GEN_862 : valid_0_84; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2399 = ~quene ? _GEN_863 : valid_0_85; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2400 = ~quene ? _GEN_864 : valid_0_86; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2401 = ~quene ? _GEN_865 : valid_0_87; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2402 = ~quene ? _GEN_866 : valid_0_88; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2403 = ~quene ? _GEN_867 : valid_0_89; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2404 = ~quene ? _GEN_868 : valid_0_90; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2405 = ~quene ? _GEN_869 : valid_0_91; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2406 = ~quene ? _GEN_870 : valid_0_92; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2407 = ~quene ? _GEN_871 : valid_0_93; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2408 = ~quene ? _GEN_872 : valid_0_94; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2409 = ~quene ? _GEN_873 : valid_0_95; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2410 = ~quene ? _GEN_874 : valid_0_96; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2411 = ~quene ? _GEN_875 : valid_0_97; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2412 = ~quene ? _GEN_876 : valid_0_98; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2413 = ~quene ? _GEN_877 : valid_0_99; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2414 = ~quene ? _GEN_878 : valid_0_100; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2415 = ~quene ? _GEN_879 : valid_0_101; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2416 = ~quene ? _GEN_880 : valid_0_102; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2417 = ~quene ? _GEN_881 : valid_0_103; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2418 = ~quene ? _GEN_882 : valid_0_104; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2419 = ~quene ? _GEN_883 : valid_0_105; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2420 = ~quene ? _GEN_884 : valid_0_106; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2421 = ~quene ? _GEN_885 : valid_0_107; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2422 = ~quene ? _GEN_886 : valid_0_108; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2423 = ~quene ? _GEN_887 : valid_0_109; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2424 = ~quene ? _GEN_888 : valid_0_110; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2425 = ~quene ? _GEN_889 : valid_0_111; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2426 = ~quene ? _GEN_890 : valid_0_112; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2427 = ~quene ? _GEN_891 : valid_0_113; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2428 = ~quene ? _GEN_892 : valid_0_114; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2429 = ~quene ? _GEN_893 : valid_0_115; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2430 = ~quene ? _GEN_894 : valid_0_116; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2431 = ~quene ? _GEN_895 : valid_0_117; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2432 = ~quene ? _GEN_896 : valid_0_118; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2433 = ~quene ? _GEN_897 : valid_0_119; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2434 = ~quene ? _GEN_898 : valid_0_120; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2435 = ~quene ? _GEN_899 : valid_0_121; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2436 = ~quene ? _GEN_900 : valid_0_122; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2437 = ~quene ? _GEN_901 : valid_0_123; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2438 = ~quene ? _GEN_902 : valid_0_124; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2439 = ~quene ? _GEN_903 : valid_0_125; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2440 = ~quene ? _GEN_904 : valid_0_126; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2441 = ~quene ? _GEN_905 : valid_0_127; // @[i_cache.scala 21:26 97:34]
  wire [63:0] _GEN_2443 = ~quene ? ram_1_0 : _GEN_906; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2444 = ~quene ? ram_1_1 : _GEN_907; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2445 = ~quene ? ram_1_2 : _GEN_908; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2446 = ~quene ? ram_1_3 : _GEN_909; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2447 = ~quene ? ram_1_4 : _GEN_910; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2448 = ~quene ? ram_1_5 : _GEN_911; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2449 = ~quene ? ram_1_6 : _GEN_912; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2450 = ~quene ? ram_1_7 : _GEN_913; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2451 = ~quene ? ram_1_8 : _GEN_914; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2452 = ~quene ? ram_1_9 : _GEN_915; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2453 = ~quene ? ram_1_10 : _GEN_916; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2454 = ~quene ? ram_1_11 : _GEN_917; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2455 = ~quene ? ram_1_12 : _GEN_918; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2456 = ~quene ? ram_1_13 : _GEN_919; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2457 = ~quene ? ram_1_14 : _GEN_920; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2458 = ~quene ? ram_1_15 : _GEN_921; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2459 = ~quene ? ram_1_16 : _GEN_922; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2460 = ~quene ? ram_1_17 : _GEN_923; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2461 = ~quene ? ram_1_18 : _GEN_924; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2462 = ~quene ? ram_1_19 : _GEN_925; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2463 = ~quene ? ram_1_20 : _GEN_926; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2464 = ~quene ? ram_1_21 : _GEN_927; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2465 = ~quene ? ram_1_22 : _GEN_928; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2466 = ~quene ? ram_1_23 : _GEN_929; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2467 = ~quene ? ram_1_24 : _GEN_930; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2468 = ~quene ? ram_1_25 : _GEN_931; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2469 = ~quene ? ram_1_26 : _GEN_932; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2470 = ~quene ? ram_1_27 : _GEN_933; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2471 = ~quene ? ram_1_28 : _GEN_934; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2472 = ~quene ? ram_1_29 : _GEN_935; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2473 = ~quene ? ram_1_30 : _GEN_936; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2474 = ~quene ? ram_1_31 : _GEN_937; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2475 = ~quene ? ram_1_32 : _GEN_938; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2476 = ~quene ? ram_1_33 : _GEN_939; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2477 = ~quene ? ram_1_34 : _GEN_940; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2478 = ~quene ? ram_1_35 : _GEN_941; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2479 = ~quene ? ram_1_36 : _GEN_942; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2480 = ~quene ? ram_1_37 : _GEN_943; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2481 = ~quene ? ram_1_38 : _GEN_944; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2482 = ~quene ? ram_1_39 : _GEN_945; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2483 = ~quene ? ram_1_40 : _GEN_946; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2484 = ~quene ? ram_1_41 : _GEN_947; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2485 = ~quene ? ram_1_42 : _GEN_948; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2486 = ~quene ? ram_1_43 : _GEN_949; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2487 = ~quene ? ram_1_44 : _GEN_950; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2488 = ~quene ? ram_1_45 : _GEN_951; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2489 = ~quene ? ram_1_46 : _GEN_952; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2490 = ~quene ? ram_1_47 : _GEN_953; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2491 = ~quene ? ram_1_48 : _GEN_954; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2492 = ~quene ? ram_1_49 : _GEN_955; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2493 = ~quene ? ram_1_50 : _GEN_956; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2494 = ~quene ? ram_1_51 : _GEN_957; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2495 = ~quene ? ram_1_52 : _GEN_958; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2496 = ~quene ? ram_1_53 : _GEN_959; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2497 = ~quene ? ram_1_54 : _GEN_960; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2498 = ~quene ? ram_1_55 : _GEN_961; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2499 = ~quene ? ram_1_56 : _GEN_962; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2500 = ~quene ? ram_1_57 : _GEN_963; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2501 = ~quene ? ram_1_58 : _GEN_964; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2502 = ~quene ? ram_1_59 : _GEN_965; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2503 = ~quene ? ram_1_60 : _GEN_966; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2504 = ~quene ? ram_1_61 : _GEN_967; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2505 = ~quene ? ram_1_62 : _GEN_968; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2506 = ~quene ? ram_1_63 : _GEN_969; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2507 = ~quene ? ram_1_64 : _GEN_970; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2508 = ~quene ? ram_1_65 : _GEN_971; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2509 = ~quene ? ram_1_66 : _GEN_972; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2510 = ~quene ? ram_1_67 : _GEN_973; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2511 = ~quene ? ram_1_68 : _GEN_974; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2512 = ~quene ? ram_1_69 : _GEN_975; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2513 = ~quene ? ram_1_70 : _GEN_976; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2514 = ~quene ? ram_1_71 : _GEN_977; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2515 = ~quene ? ram_1_72 : _GEN_978; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2516 = ~quene ? ram_1_73 : _GEN_979; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2517 = ~quene ? ram_1_74 : _GEN_980; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2518 = ~quene ? ram_1_75 : _GEN_981; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2519 = ~quene ? ram_1_76 : _GEN_982; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2520 = ~quene ? ram_1_77 : _GEN_983; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2521 = ~quene ? ram_1_78 : _GEN_984; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2522 = ~quene ? ram_1_79 : _GEN_985; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2523 = ~quene ? ram_1_80 : _GEN_986; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2524 = ~quene ? ram_1_81 : _GEN_987; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2525 = ~quene ? ram_1_82 : _GEN_988; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2526 = ~quene ? ram_1_83 : _GEN_989; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2527 = ~quene ? ram_1_84 : _GEN_990; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2528 = ~quene ? ram_1_85 : _GEN_991; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2529 = ~quene ? ram_1_86 : _GEN_992; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2530 = ~quene ? ram_1_87 : _GEN_993; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2531 = ~quene ? ram_1_88 : _GEN_994; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2532 = ~quene ? ram_1_89 : _GEN_995; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2533 = ~quene ? ram_1_90 : _GEN_996; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2534 = ~quene ? ram_1_91 : _GEN_997; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2535 = ~quene ? ram_1_92 : _GEN_998; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2536 = ~quene ? ram_1_93 : _GEN_999; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2537 = ~quene ? ram_1_94 : _GEN_1000; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2538 = ~quene ? ram_1_95 : _GEN_1001; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2539 = ~quene ? ram_1_96 : _GEN_1002; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2540 = ~quene ? ram_1_97 : _GEN_1003; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2541 = ~quene ? ram_1_98 : _GEN_1004; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2542 = ~quene ? ram_1_99 : _GEN_1005; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2543 = ~quene ? ram_1_100 : _GEN_1006; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2544 = ~quene ? ram_1_101 : _GEN_1007; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2545 = ~quene ? ram_1_102 : _GEN_1008; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2546 = ~quene ? ram_1_103 : _GEN_1009; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2547 = ~quene ? ram_1_104 : _GEN_1010; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2548 = ~quene ? ram_1_105 : _GEN_1011; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2549 = ~quene ? ram_1_106 : _GEN_1012; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2550 = ~quene ? ram_1_107 : _GEN_1013; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2551 = ~quene ? ram_1_108 : _GEN_1014; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2552 = ~quene ? ram_1_109 : _GEN_1015; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2553 = ~quene ? ram_1_110 : _GEN_1016; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2554 = ~quene ? ram_1_111 : _GEN_1017; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2555 = ~quene ? ram_1_112 : _GEN_1018; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2556 = ~quene ? ram_1_113 : _GEN_1019; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2557 = ~quene ? ram_1_114 : _GEN_1020; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2558 = ~quene ? ram_1_115 : _GEN_1021; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2559 = ~quene ? ram_1_116 : _GEN_1022; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2560 = ~quene ? ram_1_117 : _GEN_1023; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2561 = ~quene ? ram_1_118 : _GEN_1024; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2562 = ~quene ? ram_1_119 : _GEN_1025; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2563 = ~quene ? ram_1_120 : _GEN_1026; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2564 = ~quene ? ram_1_121 : _GEN_1027; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2565 = ~quene ? ram_1_122 : _GEN_1028; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2566 = ~quene ? ram_1_123 : _GEN_1029; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2567 = ~quene ? ram_1_124 : _GEN_1030; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2568 = ~quene ? ram_1_125 : _GEN_1031; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2569 = ~quene ? ram_1_126 : _GEN_1032; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2570 = ~quene ? ram_1_127 : _GEN_1033; // @[i_cache.scala 18:24 97:34]
  wire [31:0] _GEN_2571 = ~quene ? tag_1_0 : _GEN_1034; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2572 = ~quene ? tag_1_1 : _GEN_1035; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2573 = ~quene ? tag_1_2 : _GEN_1036; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2574 = ~quene ? tag_1_3 : _GEN_1037; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2575 = ~quene ? tag_1_4 : _GEN_1038; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2576 = ~quene ? tag_1_5 : _GEN_1039; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2577 = ~quene ? tag_1_6 : _GEN_1040; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2578 = ~quene ? tag_1_7 : _GEN_1041; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2579 = ~quene ? tag_1_8 : _GEN_1042; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2580 = ~quene ? tag_1_9 : _GEN_1043; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2581 = ~quene ? tag_1_10 : _GEN_1044; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2582 = ~quene ? tag_1_11 : _GEN_1045; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2583 = ~quene ? tag_1_12 : _GEN_1046; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2584 = ~quene ? tag_1_13 : _GEN_1047; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2585 = ~quene ? tag_1_14 : _GEN_1048; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2586 = ~quene ? tag_1_15 : _GEN_1049; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2587 = ~quene ? tag_1_16 : _GEN_1050; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2588 = ~quene ? tag_1_17 : _GEN_1051; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2589 = ~quene ? tag_1_18 : _GEN_1052; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2590 = ~quene ? tag_1_19 : _GEN_1053; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2591 = ~quene ? tag_1_20 : _GEN_1054; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2592 = ~quene ? tag_1_21 : _GEN_1055; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2593 = ~quene ? tag_1_22 : _GEN_1056; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2594 = ~quene ? tag_1_23 : _GEN_1057; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2595 = ~quene ? tag_1_24 : _GEN_1058; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2596 = ~quene ? tag_1_25 : _GEN_1059; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2597 = ~quene ? tag_1_26 : _GEN_1060; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2598 = ~quene ? tag_1_27 : _GEN_1061; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2599 = ~quene ? tag_1_28 : _GEN_1062; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2600 = ~quene ? tag_1_29 : _GEN_1063; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2601 = ~quene ? tag_1_30 : _GEN_1064; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2602 = ~quene ? tag_1_31 : _GEN_1065; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2603 = ~quene ? tag_1_32 : _GEN_1066; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2604 = ~quene ? tag_1_33 : _GEN_1067; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2605 = ~quene ? tag_1_34 : _GEN_1068; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2606 = ~quene ? tag_1_35 : _GEN_1069; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2607 = ~quene ? tag_1_36 : _GEN_1070; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2608 = ~quene ? tag_1_37 : _GEN_1071; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2609 = ~quene ? tag_1_38 : _GEN_1072; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2610 = ~quene ? tag_1_39 : _GEN_1073; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2611 = ~quene ? tag_1_40 : _GEN_1074; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2612 = ~quene ? tag_1_41 : _GEN_1075; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2613 = ~quene ? tag_1_42 : _GEN_1076; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2614 = ~quene ? tag_1_43 : _GEN_1077; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2615 = ~quene ? tag_1_44 : _GEN_1078; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2616 = ~quene ? tag_1_45 : _GEN_1079; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2617 = ~quene ? tag_1_46 : _GEN_1080; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2618 = ~quene ? tag_1_47 : _GEN_1081; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2619 = ~quene ? tag_1_48 : _GEN_1082; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2620 = ~quene ? tag_1_49 : _GEN_1083; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2621 = ~quene ? tag_1_50 : _GEN_1084; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2622 = ~quene ? tag_1_51 : _GEN_1085; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2623 = ~quene ? tag_1_52 : _GEN_1086; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2624 = ~quene ? tag_1_53 : _GEN_1087; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2625 = ~quene ? tag_1_54 : _GEN_1088; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2626 = ~quene ? tag_1_55 : _GEN_1089; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2627 = ~quene ? tag_1_56 : _GEN_1090; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2628 = ~quene ? tag_1_57 : _GEN_1091; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2629 = ~quene ? tag_1_58 : _GEN_1092; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2630 = ~quene ? tag_1_59 : _GEN_1093; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2631 = ~quene ? tag_1_60 : _GEN_1094; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2632 = ~quene ? tag_1_61 : _GEN_1095; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2633 = ~quene ? tag_1_62 : _GEN_1096; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2634 = ~quene ? tag_1_63 : _GEN_1097; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2635 = ~quene ? tag_1_64 : _GEN_1098; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2636 = ~quene ? tag_1_65 : _GEN_1099; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2637 = ~quene ? tag_1_66 : _GEN_1100; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2638 = ~quene ? tag_1_67 : _GEN_1101; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2639 = ~quene ? tag_1_68 : _GEN_1102; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2640 = ~quene ? tag_1_69 : _GEN_1103; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2641 = ~quene ? tag_1_70 : _GEN_1104; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2642 = ~quene ? tag_1_71 : _GEN_1105; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2643 = ~quene ? tag_1_72 : _GEN_1106; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2644 = ~quene ? tag_1_73 : _GEN_1107; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2645 = ~quene ? tag_1_74 : _GEN_1108; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2646 = ~quene ? tag_1_75 : _GEN_1109; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2647 = ~quene ? tag_1_76 : _GEN_1110; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2648 = ~quene ? tag_1_77 : _GEN_1111; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2649 = ~quene ? tag_1_78 : _GEN_1112; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2650 = ~quene ? tag_1_79 : _GEN_1113; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2651 = ~quene ? tag_1_80 : _GEN_1114; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2652 = ~quene ? tag_1_81 : _GEN_1115; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2653 = ~quene ? tag_1_82 : _GEN_1116; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2654 = ~quene ? tag_1_83 : _GEN_1117; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2655 = ~quene ? tag_1_84 : _GEN_1118; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2656 = ~quene ? tag_1_85 : _GEN_1119; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2657 = ~quene ? tag_1_86 : _GEN_1120; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2658 = ~quene ? tag_1_87 : _GEN_1121; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2659 = ~quene ? tag_1_88 : _GEN_1122; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2660 = ~quene ? tag_1_89 : _GEN_1123; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2661 = ~quene ? tag_1_90 : _GEN_1124; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2662 = ~quene ? tag_1_91 : _GEN_1125; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2663 = ~quene ? tag_1_92 : _GEN_1126; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2664 = ~quene ? tag_1_93 : _GEN_1127; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2665 = ~quene ? tag_1_94 : _GEN_1128; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2666 = ~quene ? tag_1_95 : _GEN_1129; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2667 = ~quene ? tag_1_96 : _GEN_1130; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2668 = ~quene ? tag_1_97 : _GEN_1131; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2669 = ~quene ? tag_1_98 : _GEN_1132; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2670 = ~quene ? tag_1_99 : _GEN_1133; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2671 = ~quene ? tag_1_100 : _GEN_1134; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2672 = ~quene ? tag_1_101 : _GEN_1135; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2673 = ~quene ? tag_1_102 : _GEN_1136; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2674 = ~quene ? tag_1_103 : _GEN_1137; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2675 = ~quene ? tag_1_104 : _GEN_1138; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2676 = ~quene ? tag_1_105 : _GEN_1139; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2677 = ~quene ? tag_1_106 : _GEN_1140; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2678 = ~quene ? tag_1_107 : _GEN_1141; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2679 = ~quene ? tag_1_108 : _GEN_1142; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2680 = ~quene ? tag_1_109 : _GEN_1143; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2681 = ~quene ? tag_1_110 : _GEN_1144; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2682 = ~quene ? tag_1_111 : _GEN_1145; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2683 = ~quene ? tag_1_112 : _GEN_1146; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2684 = ~quene ? tag_1_113 : _GEN_1147; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2685 = ~quene ? tag_1_114 : _GEN_1148; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2686 = ~quene ? tag_1_115 : _GEN_1149; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2687 = ~quene ? tag_1_116 : _GEN_1150; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2688 = ~quene ? tag_1_117 : _GEN_1151; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2689 = ~quene ? tag_1_118 : _GEN_1152; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2690 = ~quene ? tag_1_119 : _GEN_1153; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2691 = ~quene ? tag_1_120 : _GEN_1154; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2692 = ~quene ? tag_1_121 : _GEN_1155; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2693 = ~quene ? tag_1_122 : _GEN_1156; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2694 = ~quene ? tag_1_123 : _GEN_1157; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2695 = ~quene ? tag_1_124 : _GEN_1158; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2696 = ~quene ? tag_1_125 : _GEN_1159; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2697 = ~quene ? tag_1_126 : _GEN_1160; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2698 = ~quene ? tag_1_127 : _GEN_1161; // @[i_cache.scala 20:24 97:34]
  wire  _GEN_2699 = ~quene ? valid_1_0 : _GEN_1162; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2700 = ~quene ? valid_1_1 : _GEN_1163; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2701 = ~quene ? valid_1_2 : _GEN_1164; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2702 = ~quene ? valid_1_3 : _GEN_1165; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2703 = ~quene ? valid_1_4 : _GEN_1166; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2704 = ~quene ? valid_1_5 : _GEN_1167; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2705 = ~quene ? valid_1_6 : _GEN_1168; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2706 = ~quene ? valid_1_7 : _GEN_1169; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2707 = ~quene ? valid_1_8 : _GEN_1170; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2708 = ~quene ? valid_1_9 : _GEN_1171; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2709 = ~quene ? valid_1_10 : _GEN_1172; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2710 = ~quene ? valid_1_11 : _GEN_1173; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2711 = ~quene ? valid_1_12 : _GEN_1174; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2712 = ~quene ? valid_1_13 : _GEN_1175; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2713 = ~quene ? valid_1_14 : _GEN_1176; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2714 = ~quene ? valid_1_15 : _GEN_1177; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2715 = ~quene ? valid_1_16 : _GEN_1178; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2716 = ~quene ? valid_1_17 : _GEN_1179; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2717 = ~quene ? valid_1_18 : _GEN_1180; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2718 = ~quene ? valid_1_19 : _GEN_1181; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2719 = ~quene ? valid_1_20 : _GEN_1182; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2720 = ~quene ? valid_1_21 : _GEN_1183; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2721 = ~quene ? valid_1_22 : _GEN_1184; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2722 = ~quene ? valid_1_23 : _GEN_1185; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2723 = ~quene ? valid_1_24 : _GEN_1186; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2724 = ~quene ? valid_1_25 : _GEN_1187; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2725 = ~quene ? valid_1_26 : _GEN_1188; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2726 = ~quene ? valid_1_27 : _GEN_1189; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2727 = ~quene ? valid_1_28 : _GEN_1190; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2728 = ~quene ? valid_1_29 : _GEN_1191; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2729 = ~quene ? valid_1_30 : _GEN_1192; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2730 = ~quene ? valid_1_31 : _GEN_1193; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2731 = ~quene ? valid_1_32 : _GEN_1194; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2732 = ~quene ? valid_1_33 : _GEN_1195; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2733 = ~quene ? valid_1_34 : _GEN_1196; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2734 = ~quene ? valid_1_35 : _GEN_1197; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2735 = ~quene ? valid_1_36 : _GEN_1198; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2736 = ~quene ? valid_1_37 : _GEN_1199; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2737 = ~quene ? valid_1_38 : _GEN_1200; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2738 = ~quene ? valid_1_39 : _GEN_1201; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2739 = ~quene ? valid_1_40 : _GEN_1202; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2740 = ~quene ? valid_1_41 : _GEN_1203; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2741 = ~quene ? valid_1_42 : _GEN_1204; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2742 = ~quene ? valid_1_43 : _GEN_1205; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2743 = ~quene ? valid_1_44 : _GEN_1206; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2744 = ~quene ? valid_1_45 : _GEN_1207; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2745 = ~quene ? valid_1_46 : _GEN_1208; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2746 = ~quene ? valid_1_47 : _GEN_1209; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2747 = ~quene ? valid_1_48 : _GEN_1210; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2748 = ~quene ? valid_1_49 : _GEN_1211; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2749 = ~quene ? valid_1_50 : _GEN_1212; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2750 = ~quene ? valid_1_51 : _GEN_1213; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2751 = ~quene ? valid_1_52 : _GEN_1214; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2752 = ~quene ? valid_1_53 : _GEN_1215; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2753 = ~quene ? valid_1_54 : _GEN_1216; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2754 = ~quene ? valid_1_55 : _GEN_1217; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2755 = ~quene ? valid_1_56 : _GEN_1218; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2756 = ~quene ? valid_1_57 : _GEN_1219; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2757 = ~quene ? valid_1_58 : _GEN_1220; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2758 = ~quene ? valid_1_59 : _GEN_1221; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2759 = ~quene ? valid_1_60 : _GEN_1222; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2760 = ~quene ? valid_1_61 : _GEN_1223; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2761 = ~quene ? valid_1_62 : _GEN_1224; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2762 = ~quene ? valid_1_63 : _GEN_1225; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2763 = ~quene ? valid_1_64 : _GEN_1226; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2764 = ~quene ? valid_1_65 : _GEN_1227; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2765 = ~quene ? valid_1_66 : _GEN_1228; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2766 = ~quene ? valid_1_67 : _GEN_1229; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2767 = ~quene ? valid_1_68 : _GEN_1230; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2768 = ~quene ? valid_1_69 : _GEN_1231; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2769 = ~quene ? valid_1_70 : _GEN_1232; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2770 = ~quene ? valid_1_71 : _GEN_1233; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2771 = ~quene ? valid_1_72 : _GEN_1234; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2772 = ~quene ? valid_1_73 : _GEN_1235; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2773 = ~quene ? valid_1_74 : _GEN_1236; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2774 = ~quene ? valid_1_75 : _GEN_1237; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2775 = ~quene ? valid_1_76 : _GEN_1238; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2776 = ~quene ? valid_1_77 : _GEN_1239; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2777 = ~quene ? valid_1_78 : _GEN_1240; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2778 = ~quene ? valid_1_79 : _GEN_1241; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2779 = ~quene ? valid_1_80 : _GEN_1242; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2780 = ~quene ? valid_1_81 : _GEN_1243; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2781 = ~quene ? valid_1_82 : _GEN_1244; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2782 = ~quene ? valid_1_83 : _GEN_1245; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2783 = ~quene ? valid_1_84 : _GEN_1246; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2784 = ~quene ? valid_1_85 : _GEN_1247; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2785 = ~quene ? valid_1_86 : _GEN_1248; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2786 = ~quene ? valid_1_87 : _GEN_1249; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2787 = ~quene ? valid_1_88 : _GEN_1250; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2788 = ~quene ? valid_1_89 : _GEN_1251; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2789 = ~quene ? valid_1_90 : _GEN_1252; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2790 = ~quene ? valid_1_91 : _GEN_1253; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2791 = ~quene ? valid_1_92 : _GEN_1254; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2792 = ~quene ? valid_1_93 : _GEN_1255; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2793 = ~quene ? valid_1_94 : _GEN_1256; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2794 = ~quene ? valid_1_95 : _GEN_1257; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2795 = ~quene ? valid_1_96 : _GEN_1258; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2796 = ~quene ? valid_1_97 : _GEN_1259; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2797 = ~quene ? valid_1_98 : _GEN_1260; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2798 = ~quene ? valid_1_99 : _GEN_1261; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2799 = ~quene ? valid_1_100 : _GEN_1262; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2800 = ~quene ? valid_1_101 : _GEN_1263; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2801 = ~quene ? valid_1_102 : _GEN_1264; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2802 = ~quene ? valid_1_103 : _GEN_1265; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2803 = ~quene ? valid_1_104 : _GEN_1266; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2804 = ~quene ? valid_1_105 : _GEN_1267; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2805 = ~quene ? valid_1_106 : _GEN_1268; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2806 = ~quene ? valid_1_107 : _GEN_1269; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2807 = ~quene ? valid_1_108 : _GEN_1270; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2808 = ~quene ? valid_1_109 : _GEN_1271; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2809 = ~quene ? valid_1_110 : _GEN_1272; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2810 = ~quene ? valid_1_111 : _GEN_1273; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2811 = ~quene ? valid_1_112 : _GEN_1274; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2812 = ~quene ? valid_1_113 : _GEN_1275; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2813 = ~quene ? valid_1_114 : _GEN_1276; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2814 = ~quene ? valid_1_115 : _GEN_1277; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2815 = ~quene ? valid_1_116 : _GEN_1278; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2816 = ~quene ? valid_1_117 : _GEN_1279; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2817 = ~quene ? valid_1_118 : _GEN_1280; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2818 = ~quene ? valid_1_119 : _GEN_1281; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2819 = ~quene ? valid_1_120 : _GEN_1282; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2820 = ~quene ? valid_1_121 : _GEN_1283; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2821 = ~quene ? valid_1_122 : _GEN_1284; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2822 = ~quene ? valid_1_123 : _GEN_1285; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2823 = ~quene ? valid_1_124 : _GEN_1286; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2824 = ~quene ? valid_1_125 : _GEN_1287; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2825 = ~quene ? valid_1_126 : _GEN_1288; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2826 = ~quene ? valid_1_127 : _GEN_1289; // @[i_cache.scala 22:26 97:34]
  wire [63:0] _GEN_2827 = unuse_way == 2'h2 ? _GEN_906 : _GEN_2443; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2828 = unuse_way == 2'h2 ? _GEN_907 : _GEN_2444; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2829 = unuse_way == 2'h2 ? _GEN_908 : _GEN_2445; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2830 = unuse_way == 2'h2 ? _GEN_909 : _GEN_2446; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2831 = unuse_way == 2'h2 ? _GEN_910 : _GEN_2447; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2832 = unuse_way == 2'h2 ? _GEN_911 : _GEN_2448; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2833 = unuse_way == 2'h2 ? _GEN_912 : _GEN_2449; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2834 = unuse_way == 2'h2 ? _GEN_913 : _GEN_2450; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2835 = unuse_way == 2'h2 ? _GEN_914 : _GEN_2451; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2836 = unuse_way == 2'h2 ? _GEN_915 : _GEN_2452; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2837 = unuse_way == 2'h2 ? _GEN_916 : _GEN_2453; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2838 = unuse_way == 2'h2 ? _GEN_917 : _GEN_2454; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2839 = unuse_way == 2'h2 ? _GEN_918 : _GEN_2455; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2840 = unuse_way == 2'h2 ? _GEN_919 : _GEN_2456; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2841 = unuse_way == 2'h2 ? _GEN_920 : _GEN_2457; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2842 = unuse_way == 2'h2 ? _GEN_921 : _GEN_2458; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2843 = unuse_way == 2'h2 ? _GEN_922 : _GEN_2459; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2844 = unuse_way == 2'h2 ? _GEN_923 : _GEN_2460; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2845 = unuse_way == 2'h2 ? _GEN_924 : _GEN_2461; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2846 = unuse_way == 2'h2 ? _GEN_925 : _GEN_2462; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2847 = unuse_way == 2'h2 ? _GEN_926 : _GEN_2463; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2848 = unuse_way == 2'h2 ? _GEN_927 : _GEN_2464; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2849 = unuse_way == 2'h2 ? _GEN_928 : _GEN_2465; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2850 = unuse_way == 2'h2 ? _GEN_929 : _GEN_2466; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2851 = unuse_way == 2'h2 ? _GEN_930 : _GEN_2467; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2852 = unuse_way == 2'h2 ? _GEN_931 : _GEN_2468; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2853 = unuse_way == 2'h2 ? _GEN_932 : _GEN_2469; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2854 = unuse_way == 2'h2 ? _GEN_933 : _GEN_2470; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2855 = unuse_way == 2'h2 ? _GEN_934 : _GEN_2471; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2856 = unuse_way == 2'h2 ? _GEN_935 : _GEN_2472; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2857 = unuse_way == 2'h2 ? _GEN_936 : _GEN_2473; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2858 = unuse_way == 2'h2 ? _GEN_937 : _GEN_2474; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2859 = unuse_way == 2'h2 ? _GEN_938 : _GEN_2475; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2860 = unuse_way == 2'h2 ? _GEN_939 : _GEN_2476; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2861 = unuse_way == 2'h2 ? _GEN_940 : _GEN_2477; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2862 = unuse_way == 2'h2 ? _GEN_941 : _GEN_2478; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2863 = unuse_way == 2'h2 ? _GEN_942 : _GEN_2479; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2864 = unuse_way == 2'h2 ? _GEN_943 : _GEN_2480; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2865 = unuse_way == 2'h2 ? _GEN_944 : _GEN_2481; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2866 = unuse_way == 2'h2 ? _GEN_945 : _GEN_2482; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2867 = unuse_way == 2'h2 ? _GEN_946 : _GEN_2483; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2868 = unuse_way == 2'h2 ? _GEN_947 : _GEN_2484; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2869 = unuse_way == 2'h2 ? _GEN_948 : _GEN_2485; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2870 = unuse_way == 2'h2 ? _GEN_949 : _GEN_2486; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2871 = unuse_way == 2'h2 ? _GEN_950 : _GEN_2487; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2872 = unuse_way == 2'h2 ? _GEN_951 : _GEN_2488; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2873 = unuse_way == 2'h2 ? _GEN_952 : _GEN_2489; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2874 = unuse_way == 2'h2 ? _GEN_953 : _GEN_2490; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2875 = unuse_way == 2'h2 ? _GEN_954 : _GEN_2491; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2876 = unuse_way == 2'h2 ? _GEN_955 : _GEN_2492; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2877 = unuse_way == 2'h2 ? _GEN_956 : _GEN_2493; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2878 = unuse_way == 2'h2 ? _GEN_957 : _GEN_2494; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2879 = unuse_way == 2'h2 ? _GEN_958 : _GEN_2495; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2880 = unuse_way == 2'h2 ? _GEN_959 : _GEN_2496; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2881 = unuse_way == 2'h2 ? _GEN_960 : _GEN_2497; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2882 = unuse_way == 2'h2 ? _GEN_961 : _GEN_2498; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2883 = unuse_way == 2'h2 ? _GEN_962 : _GEN_2499; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2884 = unuse_way == 2'h2 ? _GEN_963 : _GEN_2500; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2885 = unuse_way == 2'h2 ? _GEN_964 : _GEN_2501; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2886 = unuse_way == 2'h2 ? _GEN_965 : _GEN_2502; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2887 = unuse_way == 2'h2 ? _GEN_966 : _GEN_2503; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2888 = unuse_way == 2'h2 ? _GEN_967 : _GEN_2504; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2889 = unuse_way == 2'h2 ? _GEN_968 : _GEN_2505; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2890 = unuse_way == 2'h2 ? _GEN_969 : _GEN_2506; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2891 = unuse_way == 2'h2 ? _GEN_970 : _GEN_2507; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2892 = unuse_way == 2'h2 ? _GEN_971 : _GEN_2508; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2893 = unuse_way == 2'h2 ? _GEN_972 : _GEN_2509; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2894 = unuse_way == 2'h2 ? _GEN_973 : _GEN_2510; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2895 = unuse_way == 2'h2 ? _GEN_974 : _GEN_2511; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2896 = unuse_way == 2'h2 ? _GEN_975 : _GEN_2512; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2897 = unuse_way == 2'h2 ? _GEN_976 : _GEN_2513; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2898 = unuse_way == 2'h2 ? _GEN_977 : _GEN_2514; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2899 = unuse_way == 2'h2 ? _GEN_978 : _GEN_2515; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2900 = unuse_way == 2'h2 ? _GEN_979 : _GEN_2516; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2901 = unuse_way == 2'h2 ? _GEN_980 : _GEN_2517; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2902 = unuse_way == 2'h2 ? _GEN_981 : _GEN_2518; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2903 = unuse_way == 2'h2 ? _GEN_982 : _GEN_2519; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2904 = unuse_way == 2'h2 ? _GEN_983 : _GEN_2520; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2905 = unuse_way == 2'h2 ? _GEN_984 : _GEN_2521; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2906 = unuse_way == 2'h2 ? _GEN_985 : _GEN_2522; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2907 = unuse_way == 2'h2 ? _GEN_986 : _GEN_2523; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2908 = unuse_way == 2'h2 ? _GEN_987 : _GEN_2524; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2909 = unuse_way == 2'h2 ? _GEN_988 : _GEN_2525; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2910 = unuse_way == 2'h2 ? _GEN_989 : _GEN_2526; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2911 = unuse_way == 2'h2 ? _GEN_990 : _GEN_2527; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2912 = unuse_way == 2'h2 ? _GEN_991 : _GEN_2528; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2913 = unuse_way == 2'h2 ? _GEN_992 : _GEN_2529; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2914 = unuse_way == 2'h2 ? _GEN_993 : _GEN_2530; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2915 = unuse_way == 2'h2 ? _GEN_994 : _GEN_2531; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2916 = unuse_way == 2'h2 ? _GEN_995 : _GEN_2532; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2917 = unuse_way == 2'h2 ? _GEN_996 : _GEN_2533; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2918 = unuse_way == 2'h2 ? _GEN_997 : _GEN_2534; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2919 = unuse_way == 2'h2 ? _GEN_998 : _GEN_2535; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2920 = unuse_way == 2'h2 ? _GEN_999 : _GEN_2536; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2921 = unuse_way == 2'h2 ? _GEN_1000 : _GEN_2537; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2922 = unuse_way == 2'h2 ? _GEN_1001 : _GEN_2538; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2923 = unuse_way == 2'h2 ? _GEN_1002 : _GEN_2539; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2924 = unuse_way == 2'h2 ? _GEN_1003 : _GEN_2540; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2925 = unuse_way == 2'h2 ? _GEN_1004 : _GEN_2541; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2926 = unuse_way == 2'h2 ? _GEN_1005 : _GEN_2542; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2927 = unuse_way == 2'h2 ? _GEN_1006 : _GEN_2543; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2928 = unuse_way == 2'h2 ? _GEN_1007 : _GEN_2544; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2929 = unuse_way == 2'h2 ? _GEN_1008 : _GEN_2545; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2930 = unuse_way == 2'h2 ? _GEN_1009 : _GEN_2546; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2931 = unuse_way == 2'h2 ? _GEN_1010 : _GEN_2547; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2932 = unuse_way == 2'h2 ? _GEN_1011 : _GEN_2548; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2933 = unuse_way == 2'h2 ? _GEN_1012 : _GEN_2549; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2934 = unuse_way == 2'h2 ? _GEN_1013 : _GEN_2550; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2935 = unuse_way == 2'h2 ? _GEN_1014 : _GEN_2551; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2936 = unuse_way == 2'h2 ? _GEN_1015 : _GEN_2552; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2937 = unuse_way == 2'h2 ? _GEN_1016 : _GEN_2553; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2938 = unuse_way == 2'h2 ? _GEN_1017 : _GEN_2554; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2939 = unuse_way == 2'h2 ? _GEN_1018 : _GEN_2555; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2940 = unuse_way == 2'h2 ? _GEN_1019 : _GEN_2556; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2941 = unuse_way == 2'h2 ? _GEN_1020 : _GEN_2557; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2942 = unuse_way == 2'h2 ? _GEN_1021 : _GEN_2558; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2943 = unuse_way == 2'h2 ? _GEN_1022 : _GEN_2559; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2944 = unuse_way == 2'h2 ? _GEN_1023 : _GEN_2560; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2945 = unuse_way == 2'h2 ? _GEN_1024 : _GEN_2561; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2946 = unuse_way == 2'h2 ? _GEN_1025 : _GEN_2562; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2947 = unuse_way == 2'h2 ? _GEN_1026 : _GEN_2563; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2948 = unuse_way == 2'h2 ? _GEN_1027 : _GEN_2564; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2949 = unuse_way == 2'h2 ? _GEN_1028 : _GEN_2565; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2950 = unuse_way == 2'h2 ? _GEN_1029 : _GEN_2566; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2951 = unuse_way == 2'h2 ? _GEN_1030 : _GEN_2567; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2952 = unuse_way == 2'h2 ? _GEN_1031 : _GEN_2568; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2953 = unuse_way == 2'h2 ? _GEN_1032 : _GEN_2569; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2954 = unuse_way == 2'h2 ? _GEN_1033 : _GEN_2570; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2955 = unuse_way == 2'h2 ? _GEN_1034 : _GEN_2571; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2956 = unuse_way == 2'h2 ? _GEN_1035 : _GEN_2572; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2957 = unuse_way == 2'h2 ? _GEN_1036 : _GEN_2573; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2958 = unuse_way == 2'h2 ? _GEN_1037 : _GEN_2574; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2959 = unuse_way == 2'h2 ? _GEN_1038 : _GEN_2575; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2960 = unuse_way == 2'h2 ? _GEN_1039 : _GEN_2576; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2961 = unuse_way == 2'h2 ? _GEN_1040 : _GEN_2577; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2962 = unuse_way == 2'h2 ? _GEN_1041 : _GEN_2578; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2963 = unuse_way == 2'h2 ? _GEN_1042 : _GEN_2579; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2964 = unuse_way == 2'h2 ? _GEN_1043 : _GEN_2580; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2965 = unuse_way == 2'h2 ? _GEN_1044 : _GEN_2581; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2966 = unuse_way == 2'h2 ? _GEN_1045 : _GEN_2582; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2967 = unuse_way == 2'h2 ? _GEN_1046 : _GEN_2583; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2968 = unuse_way == 2'h2 ? _GEN_1047 : _GEN_2584; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2969 = unuse_way == 2'h2 ? _GEN_1048 : _GEN_2585; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2970 = unuse_way == 2'h2 ? _GEN_1049 : _GEN_2586; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2971 = unuse_way == 2'h2 ? _GEN_1050 : _GEN_2587; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2972 = unuse_way == 2'h2 ? _GEN_1051 : _GEN_2588; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2973 = unuse_way == 2'h2 ? _GEN_1052 : _GEN_2589; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2974 = unuse_way == 2'h2 ? _GEN_1053 : _GEN_2590; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2975 = unuse_way == 2'h2 ? _GEN_1054 : _GEN_2591; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2976 = unuse_way == 2'h2 ? _GEN_1055 : _GEN_2592; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2977 = unuse_way == 2'h2 ? _GEN_1056 : _GEN_2593; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2978 = unuse_way == 2'h2 ? _GEN_1057 : _GEN_2594; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2979 = unuse_way == 2'h2 ? _GEN_1058 : _GEN_2595; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2980 = unuse_way == 2'h2 ? _GEN_1059 : _GEN_2596; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2981 = unuse_way == 2'h2 ? _GEN_1060 : _GEN_2597; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2982 = unuse_way == 2'h2 ? _GEN_1061 : _GEN_2598; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2983 = unuse_way == 2'h2 ? _GEN_1062 : _GEN_2599; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2984 = unuse_way == 2'h2 ? _GEN_1063 : _GEN_2600; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2985 = unuse_way == 2'h2 ? _GEN_1064 : _GEN_2601; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2986 = unuse_way == 2'h2 ? _GEN_1065 : _GEN_2602; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2987 = unuse_way == 2'h2 ? _GEN_1066 : _GEN_2603; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2988 = unuse_way == 2'h2 ? _GEN_1067 : _GEN_2604; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2989 = unuse_way == 2'h2 ? _GEN_1068 : _GEN_2605; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2990 = unuse_way == 2'h2 ? _GEN_1069 : _GEN_2606; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2991 = unuse_way == 2'h2 ? _GEN_1070 : _GEN_2607; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2992 = unuse_way == 2'h2 ? _GEN_1071 : _GEN_2608; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2993 = unuse_way == 2'h2 ? _GEN_1072 : _GEN_2609; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2994 = unuse_way == 2'h2 ? _GEN_1073 : _GEN_2610; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2995 = unuse_way == 2'h2 ? _GEN_1074 : _GEN_2611; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2996 = unuse_way == 2'h2 ? _GEN_1075 : _GEN_2612; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2997 = unuse_way == 2'h2 ? _GEN_1076 : _GEN_2613; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2998 = unuse_way == 2'h2 ? _GEN_1077 : _GEN_2614; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2999 = unuse_way == 2'h2 ? _GEN_1078 : _GEN_2615; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3000 = unuse_way == 2'h2 ? _GEN_1079 : _GEN_2616; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3001 = unuse_way == 2'h2 ? _GEN_1080 : _GEN_2617; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3002 = unuse_way == 2'h2 ? _GEN_1081 : _GEN_2618; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3003 = unuse_way == 2'h2 ? _GEN_1082 : _GEN_2619; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3004 = unuse_way == 2'h2 ? _GEN_1083 : _GEN_2620; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3005 = unuse_way == 2'h2 ? _GEN_1084 : _GEN_2621; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3006 = unuse_way == 2'h2 ? _GEN_1085 : _GEN_2622; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3007 = unuse_way == 2'h2 ? _GEN_1086 : _GEN_2623; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3008 = unuse_way == 2'h2 ? _GEN_1087 : _GEN_2624; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3009 = unuse_way == 2'h2 ? _GEN_1088 : _GEN_2625; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3010 = unuse_way == 2'h2 ? _GEN_1089 : _GEN_2626; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3011 = unuse_way == 2'h2 ? _GEN_1090 : _GEN_2627; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3012 = unuse_way == 2'h2 ? _GEN_1091 : _GEN_2628; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3013 = unuse_way == 2'h2 ? _GEN_1092 : _GEN_2629; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3014 = unuse_way == 2'h2 ? _GEN_1093 : _GEN_2630; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3015 = unuse_way == 2'h2 ? _GEN_1094 : _GEN_2631; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3016 = unuse_way == 2'h2 ? _GEN_1095 : _GEN_2632; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3017 = unuse_way == 2'h2 ? _GEN_1096 : _GEN_2633; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3018 = unuse_way == 2'h2 ? _GEN_1097 : _GEN_2634; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3019 = unuse_way == 2'h2 ? _GEN_1098 : _GEN_2635; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3020 = unuse_way == 2'h2 ? _GEN_1099 : _GEN_2636; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3021 = unuse_way == 2'h2 ? _GEN_1100 : _GEN_2637; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3022 = unuse_way == 2'h2 ? _GEN_1101 : _GEN_2638; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3023 = unuse_way == 2'h2 ? _GEN_1102 : _GEN_2639; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3024 = unuse_way == 2'h2 ? _GEN_1103 : _GEN_2640; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3025 = unuse_way == 2'h2 ? _GEN_1104 : _GEN_2641; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3026 = unuse_way == 2'h2 ? _GEN_1105 : _GEN_2642; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3027 = unuse_way == 2'h2 ? _GEN_1106 : _GEN_2643; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3028 = unuse_way == 2'h2 ? _GEN_1107 : _GEN_2644; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3029 = unuse_way == 2'h2 ? _GEN_1108 : _GEN_2645; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3030 = unuse_way == 2'h2 ? _GEN_1109 : _GEN_2646; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3031 = unuse_way == 2'h2 ? _GEN_1110 : _GEN_2647; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3032 = unuse_way == 2'h2 ? _GEN_1111 : _GEN_2648; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3033 = unuse_way == 2'h2 ? _GEN_1112 : _GEN_2649; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3034 = unuse_way == 2'h2 ? _GEN_1113 : _GEN_2650; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3035 = unuse_way == 2'h2 ? _GEN_1114 : _GEN_2651; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3036 = unuse_way == 2'h2 ? _GEN_1115 : _GEN_2652; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3037 = unuse_way == 2'h2 ? _GEN_1116 : _GEN_2653; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3038 = unuse_way == 2'h2 ? _GEN_1117 : _GEN_2654; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3039 = unuse_way == 2'h2 ? _GEN_1118 : _GEN_2655; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3040 = unuse_way == 2'h2 ? _GEN_1119 : _GEN_2656; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3041 = unuse_way == 2'h2 ? _GEN_1120 : _GEN_2657; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3042 = unuse_way == 2'h2 ? _GEN_1121 : _GEN_2658; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3043 = unuse_way == 2'h2 ? _GEN_1122 : _GEN_2659; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3044 = unuse_way == 2'h2 ? _GEN_1123 : _GEN_2660; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3045 = unuse_way == 2'h2 ? _GEN_1124 : _GEN_2661; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3046 = unuse_way == 2'h2 ? _GEN_1125 : _GEN_2662; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3047 = unuse_way == 2'h2 ? _GEN_1126 : _GEN_2663; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3048 = unuse_way == 2'h2 ? _GEN_1127 : _GEN_2664; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3049 = unuse_way == 2'h2 ? _GEN_1128 : _GEN_2665; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3050 = unuse_way == 2'h2 ? _GEN_1129 : _GEN_2666; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3051 = unuse_way == 2'h2 ? _GEN_1130 : _GEN_2667; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3052 = unuse_way == 2'h2 ? _GEN_1131 : _GEN_2668; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3053 = unuse_way == 2'h2 ? _GEN_1132 : _GEN_2669; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3054 = unuse_way == 2'h2 ? _GEN_1133 : _GEN_2670; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3055 = unuse_way == 2'h2 ? _GEN_1134 : _GEN_2671; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3056 = unuse_way == 2'h2 ? _GEN_1135 : _GEN_2672; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3057 = unuse_way == 2'h2 ? _GEN_1136 : _GEN_2673; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3058 = unuse_way == 2'h2 ? _GEN_1137 : _GEN_2674; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3059 = unuse_way == 2'h2 ? _GEN_1138 : _GEN_2675; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3060 = unuse_way == 2'h2 ? _GEN_1139 : _GEN_2676; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3061 = unuse_way == 2'h2 ? _GEN_1140 : _GEN_2677; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3062 = unuse_way == 2'h2 ? _GEN_1141 : _GEN_2678; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3063 = unuse_way == 2'h2 ? _GEN_1142 : _GEN_2679; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3064 = unuse_way == 2'h2 ? _GEN_1143 : _GEN_2680; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3065 = unuse_way == 2'h2 ? _GEN_1144 : _GEN_2681; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3066 = unuse_way == 2'h2 ? _GEN_1145 : _GEN_2682; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3067 = unuse_way == 2'h2 ? _GEN_1146 : _GEN_2683; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3068 = unuse_way == 2'h2 ? _GEN_1147 : _GEN_2684; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3069 = unuse_way == 2'h2 ? _GEN_1148 : _GEN_2685; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3070 = unuse_way == 2'h2 ? _GEN_1149 : _GEN_2686; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3071 = unuse_way == 2'h2 ? _GEN_1150 : _GEN_2687; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3072 = unuse_way == 2'h2 ? _GEN_1151 : _GEN_2688; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3073 = unuse_way == 2'h2 ? _GEN_1152 : _GEN_2689; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3074 = unuse_way == 2'h2 ? _GEN_1153 : _GEN_2690; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3075 = unuse_way == 2'h2 ? _GEN_1154 : _GEN_2691; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3076 = unuse_way == 2'h2 ? _GEN_1155 : _GEN_2692; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3077 = unuse_way == 2'h2 ? _GEN_1156 : _GEN_2693; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3078 = unuse_way == 2'h2 ? _GEN_1157 : _GEN_2694; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3079 = unuse_way == 2'h2 ? _GEN_1158 : _GEN_2695; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3080 = unuse_way == 2'h2 ? _GEN_1159 : _GEN_2696; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3081 = unuse_way == 2'h2 ? _GEN_1160 : _GEN_2697; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3082 = unuse_way == 2'h2 ? _GEN_1161 : _GEN_2698; // @[i_cache.scala 91:40]
  wire  _GEN_3083 = unuse_way == 2'h2 ? _GEN_1162 : _GEN_2699; // @[i_cache.scala 91:40]
  wire  _GEN_3084 = unuse_way == 2'h2 ? _GEN_1163 : _GEN_2700; // @[i_cache.scala 91:40]
  wire  _GEN_3085 = unuse_way == 2'h2 ? _GEN_1164 : _GEN_2701; // @[i_cache.scala 91:40]
  wire  _GEN_3086 = unuse_way == 2'h2 ? _GEN_1165 : _GEN_2702; // @[i_cache.scala 91:40]
  wire  _GEN_3087 = unuse_way == 2'h2 ? _GEN_1166 : _GEN_2703; // @[i_cache.scala 91:40]
  wire  _GEN_3088 = unuse_way == 2'h2 ? _GEN_1167 : _GEN_2704; // @[i_cache.scala 91:40]
  wire  _GEN_3089 = unuse_way == 2'h2 ? _GEN_1168 : _GEN_2705; // @[i_cache.scala 91:40]
  wire  _GEN_3090 = unuse_way == 2'h2 ? _GEN_1169 : _GEN_2706; // @[i_cache.scala 91:40]
  wire  _GEN_3091 = unuse_way == 2'h2 ? _GEN_1170 : _GEN_2707; // @[i_cache.scala 91:40]
  wire  _GEN_3092 = unuse_way == 2'h2 ? _GEN_1171 : _GEN_2708; // @[i_cache.scala 91:40]
  wire  _GEN_3093 = unuse_way == 2'h2 ? _GEN_1172 : _GEN_2709; // @[i_cache.scala 91:40]
  wire  _GEN_3094 = unuse_way == 2'h2 ? _GEN_1173 : _GEN_2710; // @[i_cache.scala 91:40]
  wire  _GEN_3095 = unuse_way == 2'h2 ? _GEN_1174 : _GEN_2711; // @[i_cache.scala 91:40]
  wire  _GEN_3096 = unuse_way == 2'h2 ? _GEN_1175 : _GEN_2712; // @[i_cache.scala 91:40]
  wire  _GEN_3097 = unuse_way == 2'h2 ? _GEN_1176 : _GEN_2713; // @[i_cache.scala 91:40]
  wire  _GEN_3098 = unuse_way == 2'h2 ? _GEN_1177 : _GEN_2714; // @[i_cache.scala 91:40]
  wire  _GEN_3099 = unuse_way == 2'h2 ? _GEN_1178 : _GEN_2715; // @[i_cache.scala 91:40]
  wire  _GEN_3100 = unuse_way == 2'h2 ? _GEN_1179 : _GEN_2716; // @[i_cache.scala 91:40]
  wire  _GEN_3101 = unuse_way == 2'h2 ? _GEN_1180 : _GEN_2717; // @[i_cache.scala 91:40]
  wire  _GEN_3102 = unuse_way == 2'h2 ? _GEN_1181 : _GEN_2718; // @[i_cache.scala 91:40]
  wire  _GEN_3103 = unuse_way == 2'h2 ? _GEN_1182 : _GEN_2719; // @[i_cache.scala 91:40]
  wire  _GEN_3104 = unuse_way == 2'h2 ? _GEN_1183 : _GEN_2720; // @[i_cache.scala 91:40]
  wire  _GEN_3105 = unuse_way == 2'h2 ? _GEN_1184 : _GEN_2721; // @[i_cache.scala 91:40]
  wire  _GEN_3106 = unuse_way == 2'h2 ? _GEN_1185 : _GEN_2722; // @[i_cache.scala 91:40]
  wire  _GEN_3107 = unuse_way == 2'h2 ? _GEN_1186 : _GEN_2723; // @[i_cache.scala 91:40]
  wire  _GEN_3108 = unuse_way == 2'h2 ? _GEN_1187 : _GEN_2724; // @[i_cache.scala 91:40]
  wire  _GEN_3109 = unuse_way == 2'h2 ? _GEN_1188 : _GEN_2725; // @[i_cache.scala 91:40]
  wire  _GEN_3110 = unuse_way == 2'h2 ? _GEN_1189 : _GEN_2726; // @[i_cache.scala 91:40]
  wire  _GEN_3111 = unuse_way == 2'h2 ? _GEN_1190 : _GEN_2727; // @[i_cache.scala 91:40]
  wire  _GEN_3112 = unuse_way == 2'h2 ? _GEN_1191 : _GEN_2728; // @[i_cache.scala 91:40]
  wire  _GEN_3113 = unuse_way == 2'h2 ? _GEN_1192 : _GEN_2729; // @[i_cache.scala 91:40]
  wire  _GEN_3114 = unuse_way == 2'h2 ? _GEN_1193 : _GEN_2730; // @[i_cache.scala 91:40]
  wire  _GEN_3115 = unuse_way == 2'h2 ? _GEN_1194 : _GEN_2731; // @[i_cache.scala 91:40]
  wire  _GEN_3116 = unuse_way == 2'h2 ? _GEN_1195 : _GEN_2732; // @[i_cache.scala 91:40]
  wire  _GEN_3117 = unuse_way == 2'h2 ? _GEN_1196 : _GEN_2733; // @[i_cache.scala 91:40]
  wire  _GEN_3118 = unuse_way == 2'h2 ? _GEN_1197 : _GEN_2734; // @[i_cache.scala 91:40]
  wire  _GEN_3119 = unuse_way == 2'h2 ? _GEN_1198 : _GEN_2735; // @[i_cache.scala 91:40]
  wire  _GEN_3120 = unuse_way == 2'h2 ? _GEN_1199 : _GEN_2736; // @[i_cache.scala 91:40]
  wire  _GEN_3121 = unuse_way == 2'h2 ? _GEN_1200 : _GEN_2737; // @[i_cache.scala 91:40]
  wire  _GEN_3122 = unuse_way == 2'h2 ? _GEN_1201 : _GEN_2738; // @[i_cache.scala 91:40]
  wire  _GEN_3123 = unuse_way == 2'h2 ? _GEN_1202 : _GEN_2739; // @[i_cache.scala 91:40]
  wire  _GEN_3124 = unuse_way == 2'h2 ? _GEN_1203 : _GEN_2740; // @[i_cache.scala 91:40]
  wire  _GEN_3125 = unuse_way == 2'h2 ? _GEN_1204 : _GEN_2741; // @[i_cache.scala 91:40]
  wire  _GEN_3126 = unuse_way == 2'h2 ? _GEN_1205 : _GEN_2742; // @[i_cache.scala 91:40]
  wire  _GEN_3127 = unuse_way == 2'h2 ? _GEN_1206 : _GEN_2743; // @[i_cache.scala 91:40]
  wire  _GEN_3128 = unuse_way == 2'h2 ? _GEN_1207 : _GEN_2744; // @[i_cache.scala 91:40]
  wire  _GEN_3129 = unuse_way == 2'h2 ? _GEN_1208 : _GEN_2745; // @[i_cache.scala 91:40]
  wire  _GEN_3130 = unuse_way == 2'h2 ? _GEN_1209 : _GEN_2746; // @[i_cache.scala 91:40]
  wire  _GEN_3131 = unuse_way == 2'h2 ? _GEN_1210 : _GEN_2747; // @[i_cache.scala 91:40]
  wire  _GEN_3132 = unuse_way == 2'h2 ? _GEN_1211 : _GEN_2748; // @[i_cache.scala 91:40]
  wire  _GEN_3133 = unuse_way == 2'h2 ? _GEN_1212 : _GEN_2749; // @[i_cache.scala 91:40]
  wire  _GEN_3134 = unuse_way == 2'h2 ? _GEN_1213 : _GEN_2750; // @[i_cache.scala 91:40]
  wire  _GEN_3135 = unuse_way == 2'h2 ? _GEN_1214 : _GEN_2751; // @[i_cache.scala 91:40]
  wire  _GEN_3136 = unuse_way == 2'h2 ? _GEN_1215 : _GEN_2752; // @[i_cache.scala 91:40]
  wire  _GEN_3137 = unuse_way == 2'h2 ? _GEN_1216 : _GEN_2753; // @[i_cache.scala 91:40]
  wire  _GEN_3138 = unuse_way == 2'h2 ? _GEN_1217 : _GEN_2754; // @[i_cache.scala 91:40]
  wire  _GEN_3139 = unuse_way == 2'h2 ? _GEN_1218 : _GEN_2755; // @[i_cache.scala 91:40]
  wire  _GEN_3140 = unuse_way == 2'h2 ? _GEN_1219 : _GEN_2756; // @[i_cache.scala 91:40]
  wire  _GEN_3141 = unuse_way == 2'h2 ? _GEN_1220 : _GEN_2757; // @[i_cache.scala 91:40]
  wire  _GEN_3142 = unuse_way == 2'h2 ? _GEN_1221 : _GEN_2758; // @[i_cache.scala 91:40]
  wire  _GEN_3143 = unuse_way == 2'h2 ? _GEN_1222 : _GEN_2759; // @[i_cache.scala 91:40]
  wire  _GEN_3144 = unuse_way == 2'h2 ? _GEN_1223 : _GEN_2760; // @[i_cache.scala 91:40]
  wire  _GEN_3145 = unuse_way == 2'h2 ? _GEN_1224 : _GEN_2761; // @[i_cache.scala 91:40]
  wire  _GEN_3146 = unuse_way == 2'h2 ? _GEN_1225 : _GEN_2762; // @[i_cache.scala 91:40]
  wire  _GEN_3147 = unuse_way == 2'h2 ? _GEN_1226 : _GEN_2763; // @[i_cache.scala 91:40]
  wire  _GEN_3148 = unuse_way == 2'h2 ? _GEN_1227 : _GEN_2764; // @[i_cache.scala 91:40]
  wire  _GEN_3149 = unuse_way == 2'h2 ? _GEN_1228 : _GEN_2765; // @[i_cache.scala 91:40]
  wire  _GEN_3150 = unuse_way == 2'h2 ? _GEN_1229 : _GEN_2766; // @[i_cache.scala 91:40]
  wire  _GEN_3151 = unuse_way == 2'h2 ? _GEN_1230 : _GEN_2767; // @[i_cache.scala 91:40]
  wire  _GEN_3152 = unuse_way == 2'h2 ? _GEN_1231 : _GEN_2768; // @[i_cache.scala 91:40]
  wire  _GEN_3153 = unuse_way == 2'h2 ? _GEN_1232 : _GEN_2769; // @[i_cache.scala 91:40]
  wire  _GEN_3154 = unuse_way == 2'h2 ? _GEN_1233 : _GEN_2770; // @[i_cache.scala 91:40]
  wire  _GEN_3155 = unuse_way == 2'h2 ? _GEN_1234 : _GEN_2771; // @[i_cache.scala 91:40]
  wire  _GEN_3156 = unuse_way == 2'h2 ? _GEN_1235 : _GEN_2772; // @[i_cache.scala 91:40]
  wire  _GEN_3157 = unuse_way == 2'h2 ? _GEN_1236 : _GEN_2773; // @[i_cache.scala 91:40]
  wire  _GEN_3158 = unuse_way == 2'h2 ? _GEN_1237 : _GEN_2774; // @[i_cache.scala 91:40]
  wire  _GEN_3159 = unuse_way == 2'h2 ? _GEN_1238 : _GEN_2775; // @[i_cache.scala 91:40]
  wire  _GEN_3160 = unuse_way == 2'h2 ? _GEN_1239 : _GEN_2776; // @[i_cache.scala 91:40]
  wire  _GEN_3161 = unuse_way == 2'h2 ? _GEN_1240 : _GEN_2777; // @[i_cache.scala 91:40]
  wire  _GEN_3162 = unuse_way == 2'h2 ? _GEN_1241 : _GEN_2778; // @[i_cache.scala 91:40]
  wire  _GEN_3163 = unuse_way == 2'h2 ? _GEN_1242 : _GEN_2779; // @[i_cache.scala 91:40]
  wire  _GEN_3164 = unuse_way == 2'h2 ? _GEN_1243 : _GEN_2780; // @[i_cache.scala 91:40]
  wire  _GEN_3165 = unuse_way == 2'h2 ? _GEN_1244 : _GEN_2781; // @[i_cache.scala 91:40]
  wire  _GEN_3166 = unuse_way == 2'h2 ? _GEN_1245 : _GEN_2782; // @[i_cache.scala 91:40]
  wire  _GEN_3167 = unuse_way == 2'h2 ? _GEN_1246 : _GEN_2783; // @[i_cache.scala 91:40]
  wire  _GEN_3168 = unuse_way == 2'h2 ? _GEN_1247 : _GEN_2784; // @[i_cache.scala 91:40]
  wire  _GEN_3169 = unuse_way == 2'h2 ? _GEN_1248 : _GEN_2785; // @[i_cache.scala 91:40]
  wire  _GEN_3170 = unuse_way == 2'h2 ? _GEN_1249 : _GEN_2786; // @[i_cache.scala 91:40]
  wire  _GEN_3171 = unuse_way == 2'h2 ? _GEN_1250 : _GEN_2787; // @[i_cache.scala 91:40]
  wire  _GEN_3172 = unuse_way == 2'h2 ? _GEN_1251 : _GEN_2788; // @[i_cache.scala 91:40]
  wire  _GEN_3173 = unuse_way == 2'h2 ? _GEN_1252 : _GEN_2789; // @[i_cache.scala 91:40]
  wire  _GEN_3174 = unuse_way == 2'h2 ? _GEN_1253 : _GEN_2790; // @[i_cache.scala 91:40]
  wire  _GEN_3175 = unuse_way == 2'h2 ? _GEN_1254 : _GEN_2791; // @[i_cache.scala 91:40]
  wire  _GEN_3176 = unuse_way == 2'h2 ? _GEN_1255 : _GEN_2792; // @[i_cache.scala 91:40]
  wire  _GEN_3177 = unuse_way == 2'h2 ? _GEN_1256 : _GEN_2793; // @[i_cache.scala 91:40]
  wire  _GEN_3178 = unuse_way == 2'h2 ? _GEN_1257 : _GEN_2794; // @[i_cache.scala 91:40]
  wire  _GEN_3179 = unuse_way == 2'h2 ? _GEN_1258 : _GEN_2795; // @[i_cache.scala 91:40]
  wire  _GEN_3180 = unuse_way == 2'h2 ? _GEN_1259 : _GEN_2796; // @[i_cache.scala 91:40]
  wire  _GEN_3181 = unuse_way == 2'h2 ? _GEN_1260 : _GEN_2797; // @[i_cache.scala 91:40]
  wire  _GEN_3182 = unuse_way == 2'h2 ? _GEN_1261 : _GEN_2798; // @[i_cache.scala 91:40]
  wire  _GEN_3183 = unuse_way == 2'h2 ? _GEN_1262 : _GEN_2799; // @[i_cache.scala 91:40]
  wire  _GEN_3184 = unuse_way == 2'h2 ? _GEN_1263 : _GEN_2800; // @[i_cache.scala 91:40]
  wire  _GEN_3185 = unuse_way == 2'h2 ? _GEN_1264 : _GEN_2801; // @[i_cache.scala 91:40]
  wire  _GEN_3186 = unuse_way == 2'h2 ? _GEN_1265 : _GEN_2802; // @[i_cache.scala 91:40]
  wire  _GEN_3187 = unuse_way == 2'h2 ? _GEN_1266 : _GEN_2803; // @[i_cache.scala 91:40]
  wire  _GEN_3188 = unuse_way == 2'h2 ? _GEN_1267 : _GEN_2804; // @[i_cache.scala 91:40]
  wire  _GEN_3189 = unuse_way == 2'h2 ? _GEN_1268 : _GEN_2805; // @[i_cache.scala 91:40]
  wire  _GEN_3190 = unuse_way == 2'h2 ? _GEN_1269 : _GEN_2806; // @[i_cache.scala 91:40]
  wire  _GEN_3191 = unuse_way == 2'h2 ? _GEN_1270 : _GEN_2807; // @[i_cache.scala 91:40]
  wire  _GEN_3192 = unuse_way == 2'h2 ? _GEN_1271 : _GEN_2808; // @[i_cache.scala 91:40]
  wire  _GEN_3193 = unuse_way == 2'h2 ? _GEN_1272 : _GEN_2809; // @[i_cache.scala 91:40]
  wire  _GEN_3194 = unuse_way == 2'h2 ? _GEN_1273 : _GEN_2810; // @[i_cache.scala 91:40]
  wire  _GEN_3195 = unuse_way == 2'h2 ? _GEN_1274 : _GEN_2811; // @[i_cache.scala 91:40]
  wire  _GEN_3196 = unuse_way == 2'h2 ? _GEN_1275 : _GEN_2812; // @[i_cache.scala 91:40]
  wire  _GEN_3197 = unuse_way == 2'h2 ? _GEN_1276 : _GEN_2813; // @[i_cache.scala 91:40]
  wire  _GEN_3198 = unuse_way == 2'h2 ? _GEN_1277 : _GEN_2814; // @[i_cache.scala 91:40]
  wire  _GEN_3199 = unuse_way == 2'h2 ? _GEN_1278 : _GEN_2815; // @[i_cache.scala 91:40]
  wire  _GEN_3200 = unuse_way == 2'h2 ? _GEN_1279 : _GEN_2816; // @[i_cache.scala 91:40]
  wire  _GEN_3201 = unuse_way == 2'h2 ? _GEN_1280 : _GEN_2817; // @[i_cache.scala 91:40]
  wire  _GEN_3202 = unuse_way == 2'h2 ? _GEN_1281 : _GEN_2818; // @[i_cache.scala 91:40]
  wire  _GEN_3203 = unuse_way == 2'h2 ? _GEN_1282 : _GEN_2819; // @[i_cache.scala 91:40]
  wire  _GEN_3204 = unuse_way == 2'h2 ? _GEN_1283 : _GEN_2820; // @[i_cache.scala 91:40]
  wire  _GEN_3205 = unuse_way == 2'h2 ? _GEN_1284 : _GEN_2821; // @[i_cache.scala 91:40]
  wire  _GEN_3206 = unuse_way == 2'h2 ? _GEN_1285 : _GEN_2822; // @[i_cache.scala 91:40]
  wire  _GEN_3207 = unuse_way == 2'h2 ? _GEN_1286 : _GEN_2823; // @[i_cache.scala 91:40]
  wire  _GEN_3208 = unuse_way == 2'h2 ? _GEN_1287 : _GEN_2824; // @[i_cache.scala 91:40]
  wire  _GEN_3209 = unuse_way == 2'h2 ? _GEN_1288 : _GEN_2825; // @[i_cache.scala 91:40]
  wire  _GEN_3210 = unuse_way == 2'h2 ? _GEN_1289 : _GEN_2826; // @[i_cache.scala 91:40]
  wire  _GEN_3211 = unuse_way == 2'h2 ? 1'h0 : _T_14; // @[i_cache.scala 91:40 95:23]
  wire [63:0] _GEN_3212 = unuse_way == 2'h2 ? ram_0_0 : _GEN_2058; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3213 = unuse_way == 2'h2 ? ram_0_1 : _GEN_2059; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3214 = unuse_way == 2'h2 ? ram_0_2 : _GEN_2060; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3215 = unuse_way == 2'h2 ? ram_0_3 : _GEN_2061; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3216 = unuse_way == 2'h2 ? ram_0_4 : _GEN_2062; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3217 = unuse_way == 2'h2 ? ram_0_5 : _GEN_2063; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3218 = unuse_way == 2'h2 ? ram_0_6 : _GEN_2064; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3219 = unuse_way == 2'h2 ? ram_0_7 : _GEN_2065; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3220 = unuse_way == 2'h2 ? ram_0_8 : _GEN_2066; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3221 = unuse_way == 2'h2 ? ram_0_9 : _GEN_2067; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3222 = unuse_way == 2'h2 ? ram_0_10 : _GEN_2068; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3223 = unuse_way == 2'h2 ? ram_0_11 : _GEN_2069; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3224 = unuse_way == 2'h2 ? ram_0_12 : _GEN_2070; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3225 = unuse_way == 2'h2 ? ram_0_13 : _GEN_2071; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3226 = unuse_way == 2'h2 ? ram_0_14 : _GEN_2072; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3227 = unuse_way == 2'h2 ? ram_0_15 : _GEN_2073; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3228 = unuse_way == 2'h2 ? ram_0_16 : _GEN_2074; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3229 = unuse_way == 2'h2 ? ram_0_17 : _GEN_2075; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3230 = unuse_way == 2'h2 ? ram_0_18 : _GEN_2076; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3231 = unuse_way == 2'h2 ? ram_0_19 : _GEN_2077; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3232 = unuse_way == 2'h2 ? ram_0_20 : _GEN_2078; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3233 = unuse_way == 2'h2 ? ram_0_21 : _GEN_2079; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3234 = unuse_way == 2'h2 ? ram_0_22 : _GEN_2080; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3235 = unuse_way == 2'h2 ? ram_0_23 : _GEN_2081; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3236 = unuse_way == 2'h2 ? ram_0_24 : _GEN_2082; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3237 = unuse_way == 2'h2 ? ram_0_25 : _GEN_2083; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3238 = unuse_way == 2'h2 ? ram_0_26 : _GEN_2084; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3239 = unuse_way == 2'h2 ? ram_0_27 : _GEN_2085; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3240 = unuse_way == 2'h2 ? ram_0_28 : _GEN_2086; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3241 = unuse_way == 2'h2 ? ram_0_29 : _GEN_2087; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3242 = unuse_way == 2'h2 ? ram_0_30 : _GEN_2088; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3243 = unuse_way == 2'h2 ? ram_0_31 : _GEN_2089; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3244 = unuse_way == 2'h2 ? ram_0_32 : _GEN_2090; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3245 = unuse_way == 2'h2 ? ram_0_33 : _GEN_2091; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3246 = unuse_way == 2'h2 ? ram_0_34 : _GEN_2092; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3247 = unuse_way == 2'h2 ? ram_0_35 : _GEN_2093; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3248 = unuse_way == 2'h2 ? ram_0_36 : _GEN_2094; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3249 = unuse_way == 2'h2 ? ram_0_37 : _GEN_2095; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3250 = unuse_way == 2'h2 ? ram_0_38 : _GEN_2096; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3251 = unuse_way == 2'h2 ? ram_0_39 : _GEN_2097; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3252 = unuse_way == 2'h2 ? ram_0_40 : _GEN_2098; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3253 = unuse_way == 2'h2 ? ram_0_41 : _GEN_2099; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3254 = unuse_way == 2'h2 ? ram_0_42 : _GEN_2100; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3255 = unuse_way == 2'h2 ? ram_0_43 : _GEN_2101; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3256 = unuse_way == 2'h2 ? ram_0_44 : _GEN_2102; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3257 = unuse_way == 2'h2 ? ram_0_45 : _GEN_2103; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3258 = unuse_way == 2'h2 ? ram_0_46 : _GEN_2104; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3259 = unuse_way == 2'h2 ? ram_0_47 : _GEN_2105; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3260 = unuse_way == 2'h2 ? ram_0_48 : _GEN_2106; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3261 = unuse_way == 2'h2 ? ram_0_49 : _GEN_2107; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3262 = unuse_way == 2'h2 ? ram_0_50 : _GEN_2108; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3263 = unuse_way == 2'h2 ? ram_0_51 : _GEN_2109; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3264 = unuse_way == 2'h2 ? ram_0_52 : _GEN_2110; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3265 = unuse_way == 2'h2 ? ram_0_53 : _GEN_2111; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3266 = unuse_way == 2'h2 ? ram_0_54 : _GEN_2112; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3267 = unuse_way == 2'h2 ? ram_0_55 : _GEN_2113; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3268 = unuse_way == 2'h2 ? ram_0_56 : _GEN_2114; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3269 = unuse_way == 2'h2 ? ram_0_57 : _GEN_2115; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3270 = unuse_way == 2'h2 ? ram_0_58 : _GEN_2116; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3271 = unuse_way == 2'h2 ? ram_0_59 : _GEN_2117; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3272 = unuse_way == 2'h2 ? ram_0_60 : _GEN_2118; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3273 = unuse_way == 2'h2 ? ram_0_61 : _GEN_2119; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3274 = unuse_way == 2'h2 ? ram_0_62 : _GEN_2120; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3275 = unuse_way == 2'h2 ? ram_0_63 : _GEN_2121; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3276 = unuse_way == 2'h2 ? ram_0_64 : _GEN_2122; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3277 = unuse_way == 2'h2 ? ram_0_65 : _GEN_2123; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3278 = unuse_way == 2'h2 ? ram_0_66 : _GEN_2124; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3279 = unuse_way == 2'h2 ? ram_0_67 : _GEN_2125; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3280 = unuse_way == 2'h2 ? ram_0_68 : _GEN_2126; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3281 = unuse_way == 2'h2 ? ram_0_69 : _GEN_2127; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3282 = unuse_way == 2'h2 ? ram_0_70 : _GEN_2128; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3283 = unuse_way == 2'h2 ? ram_0_71 : _GEN_2129; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3284 = unuse_way == 2'h2 ? ram_0_72 : _GEN_2130; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3285 = unuse_way == 2'h2 ? ram_0_73 : _GEN_2131; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3286 = unuse_way == 2'h2 ? ram_0_74 : _GEN_2132; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3287 = unuse_way == 2'h2 ? ram_0_75 : _GEN_2133; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3288 = unuse_way == 2'h2 ? ram_0_76 : _GEN_2134; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3289 = unuse_way == 2'h2 ? ram_0_77 : _GEN_2135; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3290 = unuse_way == 2'h2 ? ram_0_78 : _GEN_2136; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3291 = unuse_way == 2'h2 ? ram_0_79 : _GEN_2137; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3292 = unuse_way == 2'h2 ? ram_0_80 : _GEN_2138; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3293 = unuse_way == 2'h2 ? ram_0_81 : _GEN_2139; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3294 = unuse_way == 2'h2 ? ram_0_82 : _GEN_2140; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3295 = unuse_way == 2'h2 ? ram_0_83 : _GEN_2141; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3296 = unuse_way == 2'h2 ? ram_0_84 : _GEN_2142; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3297 = unuse_way == 2'h2 ? ram_0_85 : _GEN_2143; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3298 = unuse_way == 2'h2 ? ram_0_86 : _GEN_2144; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3299 = unuse_way == 2'h2 ? ram_0_87 : _GEN_2145; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3300 = unuse_way == 2'h2 ? ram_0_88 : _GEN_2146; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3301 = unuse_way == 2'h2 ? ram_0_89 : _GEN_2147; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3302 = unuse_way == 2'h2 ? ram_0_90 : _GEN_2148; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3303 = unuse_way == 2'h2 ? ram_0_91 : _GEN_2149; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3304 = unuse_way == 2'h2 ? ram_0_92 : _GEN_2150; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3305 = unuse_way == 2'h2 ? ram_0_93 : _GEN_2151; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3306 = unuse_way == 2'h2 ? ram_0_94 : _GEN_2152; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3307 = unuse_way == 2'h2 ? ram_0_95 : _GEN_2153; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3308 = unuse_way == 2'h2 ? ram_0_96 : _GEN_2154; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3309 = unuse_way == 2'h2 ? ram_0_97 : _GEN_2155; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3310 = unuse_way == 2'h2 ? ram_0_98 : _GEN_2156; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3311 = unuse_way == 2'h2 ? ram_0_99 : _GEN_2157; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3312 = unuse_way == 2'h2 ? ram_0_100 : _GEN_2158; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3313 = unuse_way == 2'h2 ? ram_0_101 : _GEN_2159; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3314 = unuse_way == 2'h2 ? ram_0_102 : _GEN_2160; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3315 = unuse_way == 2'h2 ? ram_0_103 : _GEN_2161; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3316 = unuse_way == 2'h2 ? ram_0_104 : _GEN_2162; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3317 = unuse_way == 2'h2 ? ram_0_105 : _GEN_2163; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3318 = unuse_way == 2'h2 ? ram_0_106 : _GEN_2164; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3319 = unuse_way == 2'h2 ? ram_0_107 : _GEN_2165; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3320 = unuse_way == 2'h2 ? ram_0_108 : _GEN_2166; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3321 = unuse_way == 2'h2 ? ram_0_109 : _GEN_2167; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3322 = unuse_way == 2'h2 ? ram_0_110 : _GEN_2168; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3323 = unuse_way == 2'h2 ? ram_0_111 : _GEN_2169; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3324 = unuse_way == 2'h2 ? ram_0_112 : _GEN_2170; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3325 = unuse_way == 2'h2 ? ram_0_113 : _GEN_2171; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3326 = unuse_way == 2'h2 ? ram_0_114 : _GEN_2172; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3327 = unuse_way == 2'h2 ? ram_0_115 : _GEN_2173; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3328 = unuse_way == 2'h2 ? ram_0_116 : _GEN_2174; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3329 = unuse_way == 2'h2 ? ram_0_117 : _GEN_2175; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3330 = unuse_way == 2'h2 ? ram_0_118 : _GEN_2176; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3331 = unuse_way == 2'h2 ? ram_0_119 : _GEN_2177; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3332 = unuse_way == 2'h2 ? ram_0_120 : _GEN_2178; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3333 = unuse_way == 2'h2 ? ram_0_121 : _GEN_2179; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3334 = unuse_way == 2'h2 ? ram_0_122 : _GEN_2180; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3335 = unuse_way == 2'h2 ? ram_0_123 : _GEN_2181; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3336 = unuse_way == 2'h2 ? ram_0_124 : _GEN_2182; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3337 = unuse_way == 2'h2 ? ram_0_125 : _GEN_2183; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3338 = unuse_way == 2'h2 ? ram_0_126 : _GEN_2184; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3339 = unuse_way == 2'h2 ? ram_0_127 : _GEN_2185; // @[i_cache.scala 17:24 91:40]
  wire [31:0] _GEN_3340 = unuse_way == 2'h2 ? tag_0_0 : _GEN_2186; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3341 = unuse_way == 2'h2 ? tag_0_1 : _GEN_2187; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3342 = unuse_way == 2'h2 ? tag_0_2 : _GEN_2188; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3343 = unuse_way == 2'h2 ? tag_0_3 : _GEN_2189; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3344 = unuse_way == 2'h2 ? tag_0_4 : _GEN_2190; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3345 = unuse_way == 2'h2 ? tag_0_5 : _GEN_2191; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3346 = unuse_way == 2'h2 ? tag_0_6 : _GEN_2192; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3347 = unuse_way == 2'h2 ? tag_0_7 : _GEN_2193; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3348 = unuse_way == 2'h2 ? tag_0_8 : _GEN_2194; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3349 = unuse_way == 2'h2 ? tag_0_9 : _GEN_2195; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3350 = unuse_way == 2'h2 ? tag_0_10 : _GEN_2196; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3351 = unuse_way == 2'h2 ? tag_0_11 : _GEN_2197; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3352 = unuse_way == 2'h2 ? tag_0_12 : _GEN_2198; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3353 = unuse_way == 2'h2 ? tag_0_13 : _GEN_2199; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3354 = unuse_way == 2'h2 ? tag_0_14 : _GEN_2200; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3355 = unuse_way == 2'h2 ? tag_0_15 : _GEN_2201; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3356 = unuse_way == 2'h2 ? tag_0_16 : _GEN_2202; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3357 = unuse_way == 2'h2 ? tag_0_17 : _GEN_2203; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3358 = unuse_way == 2'h2 ? tag_0_18 : _GEN_2204; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3359 = unuse_way == 2'h2 ? tag_0_19 : _GEN_2205; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3360 = unuse_way == 2'h2 ? tag_0_20 : _GEN_2206; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3361 = unuse_way == 2'h2 ? tag_0_21 : _GEN_2207; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3362 = unuse_way == 2'h2 ? tag_0_22 : _GEN_2208; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3363 = unuse_way == 2'h2 ? tag_0_23 : _GEN_2209; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3364 = unuse_way == 2'h2 ? tag_0_24 : _GEN_2210; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3365 = unuse_way == 2'h2 ? tag_0_25 : _GEN_2211; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3366 = unuse_way == 2'h2 ? tag_0_26 : _GEN_2212; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3367 = unuse_way == 2'h2 ? tag_0_27 : _GEN_2213; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3368 = unuse_way == 2'h2 ? tag_0_28 : _GEN_2214; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3369 = unuse_way == 2'h2 ? tag_0_29 : _GEN_2215; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3370 = unuse_way == 2'h2 ? tag_0_30 : _GEN_2216; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3371 = unuse_way == 2'h2 ? tag_0_31 : _GEN_2217; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3372 = unuse_way == 2'h2 ? tag_0_32 : _GEN_2218; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3373 = unuse_way == 2'h2 ? tag_0_33 : _GEN_2219; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3374 = unuse_way == 2'h2 ? tag_0_34 : _GEN_2220; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3375 = unuse_way == 2'h2 ? tag_0_35 : _GEN_2221; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3376 = unuse_way == 2'h2 ? tag_0_36 : _GEN_2222; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3377 = unuse_way == 2'h2 ? tag_0_37 : _GEN_2223; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3378 = unuse_way == 2'h2 ? tag_0_38 : _GEN_2224; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3379 = unuse_way == 2'h2 ? tag_0_39 : _GEN_2225; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3380 = unuse_way == 2'h2 ? tag_0_40 : _GEN_2226; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3381 = unuse_way == 2'h2 ? tag_0_41 : _GEN_2227; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3382 = unuse_way == 2'h2 ? tag_0_42 : _GEN_2228; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3383 = unuse_way == 2'h2 ? tag_0_43 : _GEN_2229; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3384 = unuse_way == 2'h2 ? tag_0_44 : _GEN_2230; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3385 = unuse_way == 2'h2 ? tag_0_45 : _GEN_2231; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3386 = unuse_way == 2'h2 ? tag_0_46 : _GEN_2232; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3387 = unuse_way == 2'h2 ? tag_0_47 : _GEN_2233; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3388 = unuse_way == 2'h2 ? tag_0_48 : _GEN_2234; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3389 = unuse_way == 2'h2 ? tag_0_49 : _GEN_2235; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3390 = unuse_way == 2'h2 ? tag_0_50 : _GEN_2236; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3391 = unuse_way == 2'h2 ? tag_0_51 : _GEN_2237; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3392 = unuse_way == 2'h2 ? tag_0_52 : _GEN_2238; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3393 = unuse_way == 2'h2 ? tag_0_53 : _GEN_2239; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3394 = unuse_way == 2'h2 ? tag_0_54 : _GEN_2240; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3395 = unuse_way == 2'h2 ? tag_0_55 : _GEN_2241; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3396 = unuse_way == 2'h2 ? tag_0_56 : _GEN_2242; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3397 = unuse_way == 2'h2 ? tag_0_57 : _GEN_2243; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3398 = unuse_way == 2'h2 ? tag_0_58 : _GEN_2244; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3399 = unuse_way == 2'h2 ? tag_0_59 : _GEN_2245; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3400 = unuse_way == 2'h2 ? tag_0_60 : _GEN_2246; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3401 = unuse_way == 2'h2 ? tag_0_61 : _GEN_2247; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3402 = unuse_way == 2'h2 ? tag_0_62 : _GEN_2248; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3403 = unuse_way == 2'h2 ? tag_0_63 : _GEN_2249; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3404 = unuse_way == 2'h2 ? tag_0_64 : _GEN_2250; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3405 = unuse_way == 2'h2 ? tag_0_65 : _GEN_2251; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3406 = unuse_way == 2'h2 ? tag_0_66 : _GEN_2252; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3407 = unuse_way == 2'h2 ? tag_0_67 : _GEN_2253; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3408 = unuse_way == 2'h2 ? tag_0_68 : _GEN_2254; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3409 = unuse_way == 2'h2 ? tag_0_69 : _GEN_2255; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3410 = unuse_way == 2'h2 ? tag_0_70 : _GEN_2256; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3411 = unuse_way == 2'h2 ? tag_0_71 : _GEN_2257; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3412 = unuse_way == 2'h2 ? tag_0_72 : _GEN_2258; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3413 = unuse_way == 2'h2 ? tag_0_73 : _GEN_2259; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3414 = unuse_way == 2'h2 ? tag_0_74 : _GEN_2260; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3415 = unuse_way == 2'h2 ? tag_0_75 : _GEN_2261; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3416 = unuse_way == 2'h2 ? tag_0_76 : _GEN_2262; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3417 = unuse_way == 2'h2 ? tag_0_77 : _GEN_2263; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3418 = unuse_way == 2'h2 ? tag_0_78 : _GEN_2264; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3419 = unuse_way == 2'h2 ? tag_0_79 : _GEN_2265; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3420 = unuse_way == 2'h2 ? tag_0_80 : _GEN_2266; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3421 = unuse_way == 2'h2 ? tag_0_81 : _GEN_2267; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3422 = unuse_way == 2'h2 ? tag_0_82 : _GEN_2268; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3423 = unuse_way == 2'h2 ? tag_0_83 : _GEN_2269; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3424 = unuse_way == 2'h2 ? tag_0_84 : _GEN_2270; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3425 = unuse_way == 2'h2 ? tag_0_85 : _GEN_2271; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3426 = unuse_way == 2'h2 ? tag_0_86 : _GEN_2272; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3427 = unuse_way == 2'h2 ? tag_0_87 : _GEN_2273; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3428 = unuse_way == 2'h2 ? tag_0_88 : _GEN_2274; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3429 = unuse_way == 2'h2 ? tag_0_89 : _GEN_2275; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3430 = unuse_way == 2'h2 ? tag_0_90 : _GEN_2276; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3431 = unuse_way == 2'h2 ? tag_0_91 : _GEN_2277; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3432 = unuse_way == 2'h2 ? tag_0_92 : _GEN_2278; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3433 = unuse_way == 2'h2 ? tag_0_93 : _GEN_2279; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3434 = unuse_way == 2'h2 ? tag_0_94 : _GEN_2280; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3435 = unuse_way == 2'h2 ? tag_0_95 : _GEN_2281; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3436 = unuse_way == 2'h2 ? tag_0_96 : _GEN_2282; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3437 = unuse_way == 2'h2 ? tag_0_97 : _GEN_2283; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3438 = unuse_way == 2'h2 ? tag_0_98 : _GEN_2284; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3439 = unuse_way == 2'h2 ? tag_0_99 : _GEN_2285; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3440 = unuse_way == 2'h2 ? tag_0_100 : _GEN_2286; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3441 = unuse_way == 2'h2 ? tag_0_101 : _GEN_2287; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3442 = unuse_way == 2'h2 ? tag_0_102 : _GEN_2288; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3443 = unuse_way == 2'h2 ? tag_0_103 : _GEN_2289; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3444 = unuse_way == 2'h2 ? tag_0_104 : _GEN_2290; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3445 = unuse_way == 2'h2 ? tag_0_105 : _GEN_2291; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3446 = unuse_way == 2'h2 ? tag_0_106 : _GEN_2292; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3447 = unuse_way == 2'h2 ? tag_0_107 : _GEN_2293; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3448 = unuse_way == 2'h2 ? tag_0_108 : _GEN_2294; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3449 = unuse_way == 2'h2 ? tag_0_109 : _GEN_2295; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3450 = unuse_way == 2'h2 ? tag_0_110 : _GEN_2296; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3451 = unuse_way == 2'h2 ? tag_0_111 : _GEN_2297; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3452 = unuse_way == 2'h2 ? tag_0_112 : _GEN_2298; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3453 = unuse_way == 2'h2 ? tag_0_113 : _GEN_2299; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3454 = unuse_way == 2'h2 ? tag_0_114 : _GEN_2300; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3455 = unuse_way == 2'h2 ? tag_0_115 : _GEN_2301; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3456 = unuse_way == 2'h2 ? tag_0_116 : _GEN_2302; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3457 = unuse_way == 2'h2 ? tag_0_117 : _GEN_2303; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3458 = unuse_way == 2'h2 ? tag_0_118 : _GEN_2304; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3459 = unuse_way == 2'h2 ? tag_0_119 : _GEN_2305; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3460 = unuse_way == 2'h2 ? tag_0_120 : _GEN_2306; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3461 = unuse_way == 2'h2 ? tag_0_121 : _GEN_2307; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3462 = unuse_way == 2'h2 ? tag_0_122 : _GEN_2308; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3463 = unuse_way == 2'h2 ? tag_0_123 : _GEN_2309; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3464 = unuse_way == 2'h2 ? tag_0_124 : _GEN_2310; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3465 = unuse_way == 2'h2 ? tag_0_125 : _GEN_2311; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3466 = unuse_way == 2'h2 ? tag_0_126 : _GEN_2312; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3467 = unuse_way == 2'h2 ? tag_0_127 : _GEN_2313; // @[i_cache.scala 19:24 91:40]
  wire  _GEN_3468 = unuse_way == 2'h2 ? valid_0_0 : _GEN_2314; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3469 = unuse_way == 2'h2 ? valid_0_1 : _GEN_2315; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3470 = unuse_way == 2'h2 ? valid_0_2 : _GEN_2316; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3471 = unuse_way == 2'h2 ? valid_0_3 : _GEN_2317; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3472 = unuse_way == 2'h2 ? valid_0_4 : _GEN_2318; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3473 = unuse_way == 2'h2 ? valid_0_5 : _GEN_2319; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3474 = unuse_way == 2'h2 ? valid_0_6 : _GEN_2320; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3475 = unuse_way == 2'h2 ? valid_0_7 : _GEN_2321; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3476 = unuse_way == 2'h2 ? valid_0_8 : _GEN_2322; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3477 = unuse_way == 2'h2 ? valid_0_9 : _GEN_2323; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3478 = unuse_way == 2'h2 ? valid_0_10 : _GEN_2324; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3479 = unuse_way == 2'h2 ? valid_0_11 : _GEN_2325; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3480 = unuse_way == 2'h2 ? valid_0_12 : _GEN_2326; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3481 = unuse_way == 2'h2 ? valid_0_13 : _GEN_2327; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3482 = unuse_way == 2'h2 ? valid_0_14 : _GEN_2328; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3483 = unuse_way == 2'h2 ? valid_0_15 : _GEN_2329; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3484 = unuse_way == 2'h2 ? valid_0_16 : _GEN_2330; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3485 = unuse_way == 2'h2 ? valid_0_17 : _GEN_2331; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3486 = unuse_way == 2'h2 ? valid_0_18 : _GEN_2332; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3487 = unuse_way == 2'h2 ? valid_0_19 : _GEN_2333; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3488 = unuse_way == 2'h2 ? valid_0_20 : _GEN_2334; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3489 = unuse_way == 2'h2 ? valid_0_21 : _GEN_2335; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3490 = unuse_way == 2'h2 ? valid_0_22 : _GEN_2336; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3491 = unuse_way == 2'h2 ? valid_0_23 : _GEN_2337; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3492 = unuse_way == 2'h2 ? valid_0_24 : _GEN_2338; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3493 = unuse_way == 2'h2 ? valid_0_25 : _GEN_2339; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3494 = unuse_way == 2'h2 ? valid_0_26 : _GEN_2340; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3495 = unuse_way == 2'h2 ? valid_0_27 : _GEN_2341; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3496 = unuse_way == 2'h2 ? valid_0_28 : _GEN_2342; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3497 = unuse_way == 2'h2 ? valid_0_29 : _GEN_2343; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3498 = unuse_way == 2'h2 ? valid_0_30 : _GEN_2344; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3499 = unuse_way == 2'h2 ? valid_0_31 : _GEN_2345; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3500 = unuse_way == 2'h2 ? valid_0_32 : _GEN_2346; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3501 = unuse_way == 2'h2 ? valid_0_33 : _GEN_2347; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3502 = unuse_way == 2'h2 ? valid_0_34 : _GEN_2348; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3503 = unuse_way == 2'h2 ? valid_0_35 : _GEN_2349; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3504 = unuse_way == 2'h2 ? valid_0_36 : _GEN_2350; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3505 = unuse_way == 2'h2 ? valid_0_37 : _GEN_2351; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3506 = unuse_way == 2'h2 ? valid_0_38 : _GEN_2352; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3507 = unuse_way == 2'h2 ? valid_0_39 : _GEN_2353; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3508 = unuse_way == 2'h2 ? valid_0_40 : _GEN_2354; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3509 = unuse_way == 2'h2 ? valid_0_41 : _GEN_2355; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3510 = unuse_way == 2'h2 ? valid_0_42 : _GEN_2356; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3511 = unuse_way == 2'h2 ? valid_0_43 : _GEN_2357; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3512 = unuse_way == 2'h2 ? valid_0_44 : _GEN_2358; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3513 = unuse_way == 2'h2 ? valid_0_45 : _GEN_2359; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3514 = unuse_way == 2'h2 ? valid_0_46 : _GEN_2360; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3515 = unuse_way == 2'h2 ? valid_0_47 : _GEN_2361; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3516 = unuse_way == 2'h2 ? valid_0_48 : _GEN_2362; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3517 = unuse_way == 2'h2 ? valid_0_49 : _GEN_2363; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3518 = unuse_way == 2'h2 ? valid_0_50 : _GEN_2364; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3519 = unuse_way == 2'h2 ? valid_0_51 : _GEN_2365; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3520 = unuse_way == 2'h2 ? valid_0_52 : _GEN_2366; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3521 = unuse_way == 2'h2 ? valid_0_53 : _GEN_2367; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3522 = unuse_way == 2'h2 ? valid_0_54 : _GEN_2368; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3523 = unuse_way == 2'h2 ? valid_0_55 : _GEN_2369; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3524 = unuse_way == 2'h2 ? valid_0_56 : _GEN_2370; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3525 = unuse_way == 2'h2 ? valid_0_57 : _GEN_2371; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3526 = unuse_way == 2'h2 ? valid_0_58 : _GEN_2372; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3527 = unuse_way == 2'h2 ? valid_0_59 : _GEN_2373; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3528 = unuse_way == 2'h2 ? valid_0_60 : _GEN_2374; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3529 = unuse_way == 2'h2 ? valid_0_61 : _GEN_2375; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3530 = unuse_way == 2'h2 ? valid_0_62 : _GEN_2376; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3531 = unuse_way == 2'h2 ? valid_0_63 : _GEN_2377; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3532 = unuse_way == 2'h2 ? valid_0_64 : _GEN_2378; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3533 = unuse_way == 2'h2 ? valid_0_65 : _GEN_2379; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3534 = unuse_way == 2'h2 ? valid_0_66 : _GEN_2380; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3535 = unuse_way == 2'h2 ? valid_0_67 : _GEN_2381; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3536 = unuse_way == 2'h2 ? valid_0_68 : _GEN_2382; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3537 = unuse_way == 2'h2 ? valid_0_69 : _GEN_2383; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3538 = unuse_way == 2'h2 ? valid_0_70 : _GEN_2384; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3539 = unuse_way == 2'h2 ? valid_0_71 : _GEN_2385; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3540 = unuse_way == 2'h2 ? valid_0_72 : _GEN_2386; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3541 = unuse_way == 2'h2 ? valid_0_73 : _GEN_2387; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3542 = unuse_way == 2'h2 ? valid_0_74 : _GEN_2388; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3543 = unuse_way == 2'h2 ? valid_0_75 : _GEN_2389; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3544 = unuse_way == 2'h2 ? valid_0_76 : _GEN_2390; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3545 = unuse_way == 2'h2 ? valid_0_77 : _GEN_2391; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3546 = unuse_way == 2'h2 ? valid_0_78 : _GEN_2392; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3547 = unuse_way == 2'h2 ? valid_0_79 : _GEN_2393; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3548 = unuse_way == 2'h2 ? valid_0_80 : _GEN_2394; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3549 = unuse_way == 2'h2 ? valid_0_81 : _GEN_2395; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3550 = unuse_way == 2'h2 ? valid_0_82 : _GEN_2396; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3551 = unuse_way == 2'h2 ? valid_0_83 : _GEN_2397; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3552 = unuse_way == 2'h2 ? valid_0_84 : _GEN_2398; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3553 = unuse_way == 2'h2 ? valid_0_85 : _GEN_2399; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3554 = unuse_way == 2'h2 ? valid_0_86 : _GEN_2400; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3555 = unuse_way == 2'h2 ? valid_0_87 : _GEN_2401; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3556 = unuse_way == 2'h2 ? valid_0_88 : _GEN_2402; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3557 = unuse_way == 2'h2 ? valid_0_89 : _GEN_2403; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3558 = unuse_way == 2'h2 ? valid_0_90 : _GEN_2404; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3559 = unuse_way == 2'h2 ? valid_0_91 : _GEN_2405; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3560 = unuse_way == 2'h2 ? valid_0_92 : _GEN_2406; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3561 = unuse_way == 2'h2 ? valid_0_93 : _GEN_2407; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3562 = unuse_way == 2'h2 ? valid_0_94 : _GEN_2408; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3563 = unuse_way == 2'h2 ? valid_0_95 : _GEN_2409; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3564 = unuse_way == 2'h2 ? valid_0_96 : _GEN_2410; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3565 = unuse_way == 2'h2 ? valid_0_97 : _GEN_2411; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3566 = unuse_way == 2'h2 ? valid_0_98 : _GEN_2412; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3567 = unuse_way == 2'h2 ? valid_0_99 : _GEN_2413; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3568 = unuse_way == 2'h2 ? valid_0_100 : _GEN_2414; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3569 = unuse_way == 2'h2 ? valid_0_101 : _GEN_2415; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3570 = unuse_way == 2'h2 ? valid_0_102 : _GEN_2416; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3571 = unuse_way == 2'h2 ? valid_0_103 : _GEN_2417; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3572 = unuse_way == 2'h2 ? valid_0_104 : _GEN_2418; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3573 = unuse_way == 2'h2 ? valid_0_105 : _GEN_2419; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3574 = unuse_way == 2'h2 ? valid_0_106 : _GEN_2420; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3575 = unuse_way == 2'h2 ? valid_0_107 : _GEN_2421; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3576 = unuse_way == 2'h2 ? valid_0_108 : _GEN_2422; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3577 = unuse_way == 2'h2 ? valid_0_109 : _GEN_2423; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3578 = unuse_way == 2'h2 ? valid_0_110 : _GEN_2424; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3579 = unuse_way == 2'h2 ? valid_0_111 : _GEN_2425; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3580 = unuse_way == 2'h2 ? valid_0_112 : _GEN_2426; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3581 = unuse_way == 2'h2 ? valid_0_113 : _GEN_2427; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3582 = unuse_way == 2'h2 ? valid_0_114 : _GEN_2428; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3583 = unuse_way == 2'h2 ? valid_0_115 : _GEN_2429; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3584 = unuse_way == 2'h2 ? valid_0_116 : _GEN_2430; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3585 = unuse_way == 2'h2 ? valid_0_117 : _GEN_2431; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3586 = unuse_way == 2'h2 ? valid_0_118 : _GEN_2432; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3587 = unuse_way == 2'h2 ? valid_0_119 : _GEN_2433; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3588 = unuse_way == 2'h2 ? valid_0_120 : _GEN_2434; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3589 = unuse_way == 2'h2 ? valid_0_121 : _GEN_2435; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3590 = unuse_way == 2'h2 ? valid_0_122 : _GEN_2436; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3591 = unuse_way == 2'h2 ? valid_0_123 : _GEN_2437; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3592 = unuse_way == 2'h2 ? valid_0_124 : _GEN_2438; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3593 = unuse_way == 2'h2 ? valid_0_125 : _GEN_2439; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3594 = unuse_way == 2'h2 ? valid_0_126 : _GEN_2440; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3595 = unuse_way == 2'h2 ? valid_0_127 : _GEN_2441; // @[i_cache.scala 21:26 91:40]
  wire [63:0] _GEN_3596 = unuse_way == 2'h1 ? _GEN_522 : _GEN_3212; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3597 = unuse_way == 2'h1 ? _GEN_523 : _GEN_3213; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3598 = unuse_way == 2'h1 ? _GEN_524 : _GEN_3214; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3599 = unuse_way == 2'h1 ? _GEN_525 : _GEN_3215; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3600 = unuse_way == 2'h1 ? _GEN_526 : _GEN_3216; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3601 = unuse_way == 2'h1 ? _GEN_527 : _GEN_3217; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3602 = unuse_way == 2'h1 ? _GEN_528 : _GEN_3218; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3603 = unuse_way == 2'h1 ? _GEN_529 : _GEN_3219; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3604 = unuse_way == 2'h1 ? _GEN_530 : _GEN_3220; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3605 = unuse_way == 2'h1 ? _GEN_531 : _GEN_3221; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3606 = unuse_way == 2'h1 ? _GEN_532 : _GEN_3222; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3607 = unuse_way == 2'h1 ? _GEN_533 : _GEN_3223; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3608 = unuse_way == 2'h1 ? _GEN_534 : _GEN_3224; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3609 = unuse_way == 2'h1 ? _GEN_535 : _GEN_3225; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3610 = unuse_way == 2'h1 ? _GEN_536 : _GEN_3226; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3611 = unuse_way == 2'h1 ? _GEN_537 : _GEN_3227; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3612 = unuse_way == 2'h1 ? _GEN_538 : _GEN_3228; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3613 = unuse_way == 2'h1 ? _GEN_539 : _GEN_3229; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3614 = unuse_way == 2'h1 ? _GEN_540 : _GEN_3230; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3615 = unuse_way == 2'h1 ? _GEN_541 : _GEN_3231; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3616 = unuse_way == 2'h1 ? _GEN_542 : _GEN_3232; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3617 = unuse_way == 2'h1 ? _GEN_543 : _GEN_3233; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3618 = unuse_way == 2'h1 ? _GEN_544 : _GEN_3234; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3619 = unuse_way == 2'h1 ? _GEN_545 : _GEN_3235; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3620 = unuse_way == 2'h1 ? _GEN_546 : _GEN_3236; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3621 = unuse_way == 2'h1 ? _GEN_547 : _GEN_3237; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3622 = unuse_way == 2'h1 ? _GEN_548 : _GEN_3238; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3623 = unuse_way == 2'h1 ? _GEN_549 : _GEN_3239; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3624 = unuse_way == 2'h1 ? _GEN_550 : _GEN_3240; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3625 = unuse_way == 2'h1 ? _GEN_551 : _GEN_3241; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3626 = unuse_way == 2'h1 ? _GEN_552 : _GEN_3242; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3627 = unuse_way == 2'h1 ? _GEN_553 : _GEN_3243; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3628 = unuse_way == 2'h1 ? _GEN_554 : _GEN_3244; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3629 = unuse_way == 2'h1 ? _GEN_555 : _GEN_3245; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3630 = unuse_way == 2'h1 ? _GEN_556 : _GEN_3246; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3631 = unuse_way == 2'h1 ? _GEN_557 : _GEN_3247; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3632 = unuse_way == 2'h1 ? _GEN_558 : _GEN_3248; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3633 = unuse_way == 2'h1 ? _GEN_559 : _GEN_3249; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3634 = unuse_way == 2'h1 ? _GEN_560 : _GEN_3250; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3635 = unuse_way == 2'h1 ? _GEN_561 : _GEN_3251; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3636 = unuse_way == 2'h1 ? _GEN_562 : _GEN_3252; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3637 = unuse_way == 2'h1 ? _GEN_563 : _GEN_3253; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3638 = unuse_way == 2'h1 ? _GEN_564 : _GEN_3254; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3639 = unuse_way == 2'h1 ? _GEN_565 : _GEN_3255; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3640 = unuse_way == 2'h1 ? _GEN_566 : _GEN_3256; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3641 = unuse_way == 2'h1 ? _GEN_567 : _GEN_3257; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3642 = unuse_way == 2'h1 ? _GEN_568 : _GEN_3258; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3643 = unuse_way == 2'h1 ? _GEN_569 : _GEN_3259; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3644 = unuse_way == 2'h1 ? _GEN_570 : _GEN_3260; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3645 = unuse_way == 2'h1 ? _GEN_571 : _GEN_3261; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3646 = unuse_way == 2'h1 ? _GEN_572 : _GEN_3262; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3647 = unuse_way == 2'h1 ? _GEN_573 : _GEN_3263; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3648 = unuse_way == 2'h1 ? _GEN_574 : _GEN_3264; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3649 = unuse_way == 2'h1 ? _GEN_575 : _GEN_3265; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3650 = unuse_way == 2'h1 ? _GEN_576 : _GEN_3266; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3651 = unuse_way == 2'h1 ? _GEN_577 : _GEN_3267; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3652 = unuse_way == 2'h1 ? _GEN_578 : _GEN_3268; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3653 = unuse_way == 2'h1 ? _GEN_579 : _GEN_3269; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3654 = unuse_way == 2'h1 ? _GEN_580 : _GEN_3270; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3655 = unuse_way == 2'h1 ? _GEN_581 : _GEN_3271; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3656 = unuse_way == 2'h1 ? _GEN_582 : _GEN_3272; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3657 = unuse_way == 2'h1 ? _GEN_583 : _GEN_3273; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3658 = unuse_way == 2'h1 ? _GEN_584 : _GEN_3274; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3659 = unuse_way == 2'h1 ? _GEN_585 : _GEN_3275; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3660 = unuse_way == 2'h1 ? _GEN_586 : _GEN_3276; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3661 = unuse_way == 2'h1 ? _GEN_587 : _GEN_3277; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3662 = unuse_way == 2'h1 ? _GEN_588 : _GEN_3278; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3663 = unuse_way == 2'h1 ? _GEN_589 : _GEN_3279; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3664 = unuse_way == 2'h1 ? _GEN_590 : _GEN_3280; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3665 = unuse_way == 2'h1 ? _GEN_591 : _GEN_3281; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3666 = unuse_way == 2'h1 ? _GEN_592 : _GEN_3282; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3667 = unuse_way == 2'h1 ? _GEN_593 : _GEN_3283; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3668 = unuse_way == 2'h1 ? _GEN_594 : _GEN_3284; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3669 = unuse_way == 2'h1 ? _GEN_595 : _GEN_3285; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3670 = unuse_way == 2'h1 ? _GEN_596 : _GEN_3286; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3671 = unuse_way == 2'h1 ? _GEN_597 : _GEN_3287; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3672 = unuse_way == 2'h1 ? _GEN_598 : _GEN_3288; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3673 = unuse_way == 2'h1 ? _GEN_599 : _GEN_3289; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3674 = unuse_way == 2'h1 ? _GEN_600 : _GEN_3290; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3675 = unuse_way == 2'h1 ? _GEN_601 : _GEN_3291; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3676 = unuse_way == 2'h1 ? _GEN_602 : _GEN_3292; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3677 = unuse_way == 2'h1 ? _GEN_603 : _GEN_3293; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3678 = unuse_way == 2'h1 ? _GEN_604 : _GEN_3294; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3679 = unuse_way == 2'h1 ? _GEN_605 : _GEN_3295; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3680 = unuse_way == 2'h1 ? _GEN_606 : _GEN_3296; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3681 = unuse_way == 2'h1 ? _GEN_607 : _GEN_3297; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3682 = unuse_way == 2'h1 ? _GEN_608 : _GEN_3298; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3683 = unuse_way == 2'h1 ? _GEN_609 : _GEN_3299; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3684 = unuse_way == 2'h1 ? _GEN_610 : _GEN_3300; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3685 = unuse_way == 2'h1 ? _GEN_611 : _GEN_3301; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3686 = unuse_way == 2'h1 ? _GEN_612 : _GEN_3302; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3687 = unuse_way == 2'h1 ? _GEN_613 : _GEN_3303; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3688 = unuse_way == 2'h1 ? _GEN_614 : _GEN_3304; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3689 = unuse_way == 2'h1 ? _GEN_615 : _GEN_3305; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3690 = unuse_way == 2'h1 ? _GEN_616 : _GEN_3306; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3691 = unuse_way == 2'h1 ? _GEN_617 : _GEN_3307; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3692 = unuse_way == 2'h1 ? _GEN_618 : _GEN_3308; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3693 = unuse_way == 2'h1 ? _GEN_619 : _GEN_3309; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3694 = unuse_way == 2'h1 ? _GEN_620 : _GEN_3310; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3695 = unuse_way == 2'h1 ? _GEN_621 : _GEN_3311; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3696 = unuse_way == 2'h1 ? _GEN_622 : _GEN_3312; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3697 = unuse_way == 2'h1 ? _GEN_623 : _GEN_3313; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3698 = unuse_way == 2'h1 ? _GEN_624 : _GEN_3314; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3699 = unuse_way == 2'h1 ? _GEN_625 : _GEN_3315; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3700 = unuse_way == 2'h1 ? _GEN_626 : _GEN_3316; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3701 = unuse_way == 2'h1 ? _GEN_627 : _GEN_3317; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3702 = unuse_way == 2'h1 ? _GEN_628 : _GEN_3318; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3703 = unuse_way == 2'h1 ? _GEN_629 : _GEN_3319; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3704 = unuse_way == 2'h1 ? _GEN_630 : _GEN_3320; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3705 = unuse_way == 2'h1 ? _GEN_631 : _GEN_3321; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3706 = unuse_way == 2'h1 ? _GEN_632 : _GEN_3322; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3707 = unuse_way == 2'h1 ? _GEN_633 : _GEN_3323; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3708 = unuse_way == 2'h1 ? _GEN_634 : _GEN_3324; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3709 = unuse_way == 2'h1 ? _GEN_635 : _GEN_3325; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3710 = unuse_way == 2'h1 ? _GEN_636 : _GEN_3326; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3711 = unuse_way == 2'h1 ? _GEN_637 : _GEN_3327; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3712 = unuse_way == 2'h1 ? _GEN_638 : _GEN_3328; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3713 = unuse_way == 2'h1 ? _GEN_639 : _GEN_3329; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3714 = unuse_way == 2'h1 ? _GEN_640 : _GEN_3330; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3715 = unuse_way == 2'h1 ? _GEN_641 : _GEN_3331; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3716 = unuse_way == 2'h1 ? _GEN_642 : _GEN_3332; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3717 = unuse_way == 2'h1 ? _GEN_643 : _GEN_3333; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3718 = unuse_way == 2'h1 ? _GEN_644 : _GEN_3334; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3719 = unuse_way == 2'h1 ? _GEN_645 : _GEN_3335; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3720 = unuse_way == 2'h1 ? _GEN_646 : _GEN_3336; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3721 = unuse_way == 2'h1 ? _GEN_647 : _GEN_3337; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3722 = unuse_way == 2'h1 ? _GEN_648 : _GEN_3338; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3723 = unuse_way == 2'h1 ? _GEN_649 : _GEN_3339; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3724 = unuse_way == 2'h1 ? _GEN_650 : _GEN_3340; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3725 = unuse_way == 2'h1 ? _GEN_651 : _GEN_3341; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3726 = unuse_way == 2'h1 ? _GEN_652 : _GEN_3342; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3727 = unuse_way == 2'h1 ? _GEN_653 : _GEN_3343; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3728 = unuse_way == 2'h1 ? _GEN_654 : _GEN_3344; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3729 = unuse_way == 2'h1 ? _GEN_655 : _GEN_3345; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3730 = unuse_way == 2'h1 ? _GEN_656 : _GEN_3346; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3731 = unuse_way == 2'h1 ? _GEN_657 : _GEN_3347; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3732 = unuse_way == 2'h1 ? _GEN_658 : _GEN_3348; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3733 = unuse_way == 2'h1 ? _GEN_659 : _GEN_3349; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3734 = unuse_way == 2'h1 ? _GEN_660 : _GEN_3350; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3735 = unuse_way == 2'h1 ? _GEN_661 : _GEN_3351; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3736 = unuse_way == 2'h1 ? _GEN_662 : _GEN_3352; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3737 = unuse_way == 2'h1 ? _GEN_663 : _GEN_3353; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3738 = unuse_way == 2'h1 ? _GEN_664 : _GEN_3354; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3739 = unuse_way == 2'h1 ? _GEN_665 : _GEN_3355; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3740 = unuse_way == 2'h1 ? _GEN_666 : _GEN_3356; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3741 = unuse_way == 2'h1 ? _GEN_667 : _GEN_3357; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3742 = unuse_way == 2'h1 ? _GEN_668 : _GEN_3358; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3743 = unuse_way == 2'h1 ? _GEN_669 : _GEN_3359; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3744 = unuse_way == 2'h1 ? _GEN_670 : _GEN_3360; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3745 = unuse_way == 2'h1 ? _GEN_671 : _GEN_3361; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3746 = unuse_way == 2'h1 ? _GEN_672 : _GEN_3362; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3747 = unuse_way == 2'h1 ? _GEN_673 : _GEN_3363; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3748 = unuse_way == 2'h1 ? _GEN_674 : _GEN_3364; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3749 = unuse_way == 2'h1 ? _GEN_675 : _GEN_3365; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3750 = unuse_way == 2'h1 ? _GEN_676 : _GEN_3366; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3751 = unuse_way == 2'h1 ? _GEN_677 : _GEN_3367; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3752 = unuse_way == 2'h1 ? _GEN_678 : _GEN_3368; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3753 = unuse_way == 2'h1 ? _GEN_679 : _GEN_3369; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3754 = unuse_way == 2'h1 ? _GEN_680 : _GEN_3370; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3755 = unuse_way == 2'h1 ? _GEN_681 : _GEN_3371; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3756 = unuse_way == 2'h1 ? _GEN_682 : _GEN_3372; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3757 = unuse_way == 2'h1 ? _GEN_683 : _GEN_3373; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3758 = unuse_way == 2'h1 ? _GEN_684 : _GEN_3374; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3759 = unuse_way == 2'h1 ? _GEN_685 : _GEN_3375; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3760 = unuse_way == 2'h1 ? _GEN_686 : _GEN_3376; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3761 = unuse_way == 2'h1 ? _GEN_687 : _GEN_3377; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3762 = unuse_way == 2'h1 ? _GEN_688 : _GEN_3378; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3763 = unuse_way == 2'h1 ? _GEN_689 : _GEN_3379; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3764 = unuse_way == 2'h1 ? _GEN_690 : _GEN_3380; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3765 = unuse_way == 2'h1 ? _GEN_691 : _GEN_3381; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3766 = unuse_way == 2'h1 ? _GEN_692 : _GEN_3382; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3767 = unuse_way == 2'h1 ? _GEN_693 : _GEN_3383; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3768 = unuse_way == 2'h1 ? _GEN_694 : _GEN_3384; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3769 = unuse_way == 2'h1 ? _GEN_695 : _GEN_3385; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3770 = unuse_way == 2'h1 ? _GEN_696 : _GEN_3386; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3771 = unuse_way == 2'h1 ? _GEN_697 : _GEN_3387; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3772 = unuse_way == 2'h1 ? _GEN_698 : _GEN_3388; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3773 = unuse_way == 2'h1 ? _GEN_699 : _GEN_3389; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3774 = unuse_way == 2'h1 ? _GEN_700 : _GEN_3390; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3775 = unuse_way == 2'h1 ? _GEN_701 : _GEN_3391; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3776 = unuse_way == 2'h1 ? _GEN_702 : _GEN_3392; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3777 = unuse_way == 2'h1 ? _GEN_703 : _GEN_3393; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3778 = unuse_way == 2'h1 ? _GEN_704 : _GEN_3394; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3779 = unuse_way == 2'h1 ? _GEN_705 : _GEN_3395; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3780 = unuse_way == 2'h1 ? _GEN_706 : _GEN_3396; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3781 = unuse_way == 2'h1 ? _GEN_707 : _GEN_3397; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3782 = unuse_way == 2'h1 ? _GEN_708 : _GEN_3398; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3783 = unuse_way == 2'h1 ? _GEN_709 : _GEN_3399; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3784 = unuse_way == 2'h1 ? _GEN_710 : _GEN_3400; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3785 = unuse_way == 2'h1 ? _GEN_711 : _GEN_3401; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3786 = unuse_way == 2'h1 ? _GEN_712 : _GEN_3402; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3787 = unuse_way == 2'h1 ? _GEN_713 : _GEN_3403; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3788 = unuse_way == 2'h1 ? _GEN_714 : _GEN_3404; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3789 = unuse_way == 2'h1 ? _GEN_715 : _GEN_3405; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3790 = unuse_way == 2'h1 ? _GEN_716 : _GEN_3406; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3791 = unuse_way == 2'h1 ? _GEN_717 : _GEN_3407; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3792 = unuse_way == 2'h1 ? _GEN_718 : _GEN_3408; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3793 = unuse_way == 2'h1 ? _GEN_719 : _GEN_3409; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3794 = unuse_way == 2'h1 ? _GEN_720 : _GEN_3410; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3795 = unuse_way == 2'h1 ? _GEN_721 : _GEN_3411; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3796 = unuse_way == 2'h1 ? _GEN_722 : _GEN_3412; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3797 = unuse_way == 2'h1 ? _GEN_723 : _GEN_3413; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3798 = unuse_way == 2'h1 ? _GEN_724 : _GEN_3414; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3799 = unuse_way == 2'h1 ? _GEN_725 : _GEN_3415; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3800 = unuse_way == 2'h1 ? _GEN_726 : _GEN_3416; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3801 = unuse_way == 2'h1 ? _GEN_727 : _GEN_3417; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3802 = unuse_way == 2'h1 ? _GEN_728 : _GEN_3418; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3803 = unuse_way == 2'h1 ? _GEN_729 : _GEN_3419; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3804 = unuse_way == 2'h1 ? _GEN_730 : _GEN_3420; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3805 = unuse_way == 2'h1 ? _GEN_731 : _GEN_3421; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3806 = unuse_way == 2'h1 ? _GEN_732 : _GEN_3422; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3807 = unuse_way == 2'h1 ? _GEN_733 : _GEN_3423; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3808 = unuse_way == 2'h1 ? _GEN_734 : _GEN_3424; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3809 = unuse_way == 2'h1 ? _GEN_735 : _GEN_3425; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3810 = unuse_way == 2'h1 ? _GEN_736 : _GEN_3426; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3811 = unuse_way == 2'h1 ? _GEN_737 : _GEN_3427; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3812 = unuse_way == 2'h1 ? _GEN_738 : _GEN_3428; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3813 = unuse_way == 2'h1 ? _GEN_739 : _GEN_3429; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3814 = unuse_way == 2'h1 ? _GEN_740 : _GEN_3430; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3815 = unuse_way == 2'h1 ? _GEN_741 : _GEN_3431; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3816 = unuse_way == 2'h1 ? _GEN_742 : _GEN_3432; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3817 = unuse_way == 2'h1 ? _GEN_743 : _GEN_3433; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3818 = unuse_way == 2'h1 ? _GEN_744 : _GEN_3434; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3819 = unuse_way == 2'h1 ? _GEN_745 : _GEN_3435; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3820 = unuse_way == 2'h1 ? _GEN_746 : _GEN_3436; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3821 = unuse_way == 2'h1 ? _GEN_747 : _GEN_3437; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3822 = unuse_way == 2'h1 ? _GEN_748 : _GEN_3438; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3823 = unuse_way == 2'h1 ? _GEN_749 : _GEN_3439; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3824 = unuse_way == 2'h1 ? _GEN_750 : _GEN_3440; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3825 = unuse_way == 2'h1 ? _GEN_751 : _GEN_3441; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3826 = unuse_way == 2'h1 ? _GEN_752 : _GEN_3442; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3827 = unuse_way == 2'h1 ? _GEN_753 : _GEN_3443; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3828 = unuse_way == 2'h1 ? _GEN_754 : _GEN_3444; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3829 = unuse_way == 2'h1 ? _GEN_755 : _GEN_3445; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3830 = unuse_way == 2'h1 ? _GEN_756 : _GEN_3446; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3831 = unuse_way == 2'h1 ? _GEN_757 : _GEN_3447; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3832 = unuse_way == 2'h1 ? _GEN_758 : _GEN_3448; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3833 = unuse_way == 2'h1 ? _GEN_759 : _GEN_3449; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3834 = unuse_way == 2'h1 ? _GEN_760 : _GEN_3450; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3835 = unuse_way == 2'h1 ? _GEN_761 : _GEN_3451; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3836 = unuse_way == 2'h1 ? _GEN_762 : _GEN_3452; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3837 = unuse_way == 2'h1 ? _GEN_763 : _GEN_3453; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3838 = unuse_way == 2'h1 ? _GEN_764 : _GEN_3454; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3839 = unuse_way == 2'h1 ? _GEN_765 : _GEN_3455; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3840 = unuse_way == 2'h1 ? _GEN_766 : _GEN_3456; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3841 = unuse_way == 2'h1 ? _GEN_767 : _GEN_3457; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3842 = unuse_way == 2'h1 ? _GEN_768 : _GEN_3458; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3843 = unuse_way == 2'h1 ? _GEN_769 : _GEN_3459; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3844 = unuse_way == 2'h1 ? _GEN_770 : _GEN_3460; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3845 = unuse_way == 2'h1 ? _GEN_771 : _GEN_3461; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3846 = unuse_way == 2'h1 ? _GEN_772 : _GEN_3462; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3847 = unuse_way == 2'h1 ? _GEN_773 : _GEN_3463; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3848 = unuse_way == 2'h1 ? _GEN_774 : _GEN_3464; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3849 = unuse_way == 2'h1 ? _GEN_775 : _GEN_3465; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3850 = unuse_way == 2'h1 ? _GEN_776 : _GEN_3466; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3851 = unuse_way == 2'h1 ? _GEN_777 : _GEN_3467; // @[i_cache.scala 86:34]
  wire  _GEN_3852 = unuse_way == 2'h1 ? _GEN_778 : _GEN_3468; // @[i_cache.scala 86:34]
  wire  _GEN_3853 = unuse_way == 2'h1 ? _GEN_779 : _GEN_3469; // @[i_cache.scala 86:34]
  wire  _GEN_3854 = unuse_way == 2'h1 ? _GEN_780 : _GEN_3470; // @[i_cache.scala 86:34]
  wire  _GEN_3855 = unuse_way == 2'h1 ? _GEN_781 : _GEN_3471; // @[i_cache.scala 86:34]
  wire  _GEN_3856 = unuse_way == 2'h1 ? _GEN_782 : _GEN_3472; // @[i_cache.scala 86:34]
  wire  _GEN_3857 = unuse_way == 2'h1 ? _GEN_783 : _GEN_3473; // @[i_cache.scala 86:34]
  wire  _GEN_3858 = unuse_way == 2'h1 ? _GEN_784 : _GEN_3474; // @[i_cache.scala 86:34]
  wire  _GEN_3859 = unuse_way == 2'h1 ? _GEN_785 : _GEN_3475; // @[i_cache.scala 86:34]
  wire  _GEN_3860 = unuse_way == 2'h1 ? _GEN_786 : _GEN_3476; // @[i_cache.scala 86:34]
  wire  _GEN_3861 = unuse_way == 2'h1 ? _GEN_787 : _GEN_3477; // @[i_cache.scala 86:34]
  wire  _GEN_3862 = unuse_way == 2'h1 ? _GEN_788 : _GEN_3478; // @[i_cache.scala 86:34]
  wire  _GEN_3863 = unuse_way == 2'h1 ? _GEN_789 : _GEN_3479; // @[i_cache.scala 86:34]
  wire  _GEN_3864 = unuse_way == 2'h1 ? _GEN_790 : _GEN_3480; // @[i_cache.scala 86:34]
  wire  _GEN_3865 = unuse_way == 2'h1 ? _GEN_791 : _GEN_3481; // @[i_cache.scala 86:34]
  wire  _GEN_3866 = unuse_way == 2'h1 ? _GEN_792 : _GEN_3482; // @[i_cache.scala 86:34]
  wire  _GEN_3867 = unuse_way == 2'h1 ? _GEN_793 : _GEN_3483; // @[i_cache.scala 86:34]
  wire  _GEN_3868 = unuse_way == 2'h1 ? _GEN_794 : _GEN_3484; // @[i_cache.scala 86:34]
  wire  _GEN_3869 = unuse_way == 2'h1 ? _GEN_795 : _GEN_3485; // @[i_cache.scala 86:34]
  wire  _GEN_3870 = unuse_way == 2'h1 ? _GEN_796 : _GEN_3486; // @[i_cache.scala 86:34]
  wire  _GEN_3871 = unuse_way == 2'h1 ? _GEN_797 : _GEN_3487; // @[i_cache.scala 86:34]
  wire  _GEN_3872 = unuse_way == 2'h1 ? _GEN_798 : _GEN_3488; // @[i_cache.scala 86:34]
  wire  _GEN_3873 = unuse_way == 2'h1 ? _GEN_799 : _GEN_3489; // @[i_cache.scala 86:34]
  wire  _GEN_3874 = unuse_way == 2'h1 ? _GEN_800 : _GEN_3490; // @[i_cache.scala 86:34]
  wire  _GEN_3875 = unuse_way == 2'h1 ? _GEN_801 : _GEN_3491; // @[i_cache.scala 86:34]
  wire  _GEN_3876 = unuse_way == 2'h1 ? _GEN_802 : _GEN_3492; // @[i_cache.scala 86:34]
  wire  _GEN_3877 = unuse_way == 2'h1 ? _GEN_803 : _GEN_3493; // @[i_cache.scala 86:34]
  wire  _GEN_3878 = unuse_way == 2'h1 ? _GEN_804 : _GEN_3494; // @[i_cache.scala 86:34]
  wire  _GEN_3879 = unuse_way == 2'h1 ? _GEN_805 : _GEN_3495; // @[i_cache.scala 86:34]
  wire  _GEN_3880 = unuse_way == 2'h1 ? _GEN_806 : _GEN_3496; // @[i_cache.scala 86:34]
  wire  _GEN_3881 = unuse_way == 2'h1 ? _GEN_807 : _GEN_3497; // @[i_cache.scala 86:34]
  wire  _GEN_3882 = unuse_way == 2'h1 ? _GEN_808 : _GEN_3498; // @[i_cache.scala 86:34]
  wire  _GEN_3883 = unuse_way == 2'h1 ? _GEN_809 : _GEN_3499; // @[i_cache.scala 86:34]
  wire  _GEN_3884 = unuse_way == 2'h1 ? _GEN_810 : _GEN_3500; // @[i_cache.scala 86:34]
  wire  _GEN_3885 = unuse_way == 2'h1 ? _GEN_811 : _GEN_3501; // @[i_cache.scala 86:34]
  wire  _GEN_3886 = unuse_way == 2'h1 ? _GEN_812 : _GEN_3502; // @[i_cache.scala 86:34]
  wire  _GEN_3887 = unuse_way == 2'h1 ? _GEN_813 : _GEN_3503; // @[i_cache.scala 86:34]
  wire  _GEN_3888 = unuse_way == 2'h1 ? _GEN_814 : _GEN_3504; // @[i_cache.scala 86:34]
  wire  _GEN_3889 = unuse_way == 2'h1 ? _GEN_815 : _GEN_3505; // @[i_cache.scala 86:34]
  wire  _GEN_3890 = unuse_way == 2'h1 ? _GEN_816 : _GEN_3506; // @[i_cache.scala 86:34]
  wire  _GEN_3891 = unuse_way == 2'h1 ? _GEN_817 : _GEN_3507; // @[i_cache.scala 86:34]
  wire  _GEN_3892 = unuse_way == 2'h1 ? _GEN_818 : _GEN_3508; // @[i_cache.scala 86:34]
  wire  _GEN_3893 = unuse_way == 2'h1 ? _GEN_819 : _GEN_3509; // @[i_cache.scala 86:34]
  wire  _GEN_3894 = unuse_way == 2'h1 ? _GEN_820 : _GEN_3510; // @[i_cache.scala 86:34]
  wire  _GEN_3895 = unuse_way == 2'h1 ? _GEN_821 : _GEN_3511; // @[i_cache.scala 86:34]
  wire  _GEN_3896 = unuse_way == 2'h1 ? _GEN_822 : _GEN_3512; // @[i_cache.scala 86:34]
  wire  _GEN_3897 = unuse_way == 2'h1 ? _GEN_823 : _GEN_3513; // @[i_cache.scala 86:34]
  wire  _GEN_3898 = unuse_way == 2'h1 ? _GEN_824 : _GEN_3514; // @[i_cache.scala 86:34]
  wire  _GEN_3899 = unuse_way == 2'h1 ? _GEN_825 : _GEN_3515; // @[i_cache.scala 86:34]
  wire  _GEN_3900 = unuse_way == 2'h1 ? _GEN_826 : _GEN_3516; // @[i_cache.scala 86:34]
  wire  _GEN_3901 = unuse_way == 2'h1 ? _GEN_827 : _GEN_3517; // @[i_cache.scala 86:34]
  wire  _GEN_3902 = unuse_way == 2'h1 ? _GEN_828 : _GEN_3518; // @[i_cache.scala 86:34]
  wire  _GEN_3903 = unuse_way == 2'h1 ? _GEN_829 : _GEN_3519; // @[i_cache.scala 86:34]
  wire  _GEN_3904 = unuse_way == 2'h1 ? _GEN_830 : _GEN_3520; // @[i_cache.scala 86:34]
  wire  _GEN_3905 = unuse_way == 2'h1 ? _GEN_831 : _GEN_3521; // @[i_cache.scala 86:34]
  wire  _GEN_3906 = unuse_way == 2'h1 ? _GEN_832 : _GEN_3522; // @[i_cache.scala 86:34]
  wire  _GEN_3907 = unuse_way == 2'h1 ? _GEN_833 : _GEN_3523; // @[i_cache.scala 86:34]
  wire  _GEN_3908 = unuse_way == 2'h1 ? _GEN_834 : _GEN_3524; // @[i_cache.scala 86:34]
  wire  _GEN_3909 = unuse_way == 2'h1 ? _GEN_835 : _GEN_3525; // @[i_cache.scala 86:34]
  wire  _GEN_3910 = unuse_way == 2'h1 ? _GEN_836 : _GEN_3526; // @[i_cache.scala 86:34]
  wire  _GEN_3911 = unuse_way == 2'h1 ? _GEN_837 : _GEN_3527; // @[i_cache.scala 86:34]
  wire  _GEN_3912 = unuse_way == 2'h1 ? _GEN_838 : _GEN_3528; // @[i_cache.scala 86:34]
  wire  _GEN_3913 = unuse_way == 2'h1 ? _GEN_839 : _GEN_3529; // @[i_cache.scala 86:34]
  wire  _GEN_3914 = unuse_way == 2'h1 ? _GEN_840 : _GEN_3530; // @[i_cache.scala 86:34]
  wire  _GEN_3915 = unuse_way == 2'h1 ? _GEN_841 : _GEN_3531; // @[i_cache.scala 86:34]
  wire  _GEN_3916 = unuse_way == 2'h1 ? _GEN_842 : _GEN_3532; // @[i_cache.scala 86:34]
  wire  _GEN_3917 = unuse_way == 2'h1 ? _GEN_843 : _GEN_3533; // @[i_cache.scala 86:34]
  wire  _GEN_3918 = unuse_way == 2'h1 ? _GEN_844 : _GEN_3534; // @[i_cache.scala 86:34]
  wire  _GEN_3919 = unuse_way == 2'h1 ? _GEN_845 : _GEN_3535; // @[i_cache.scala 86:34]
  wire  _GEN_3920 = unuse_way == 2'h1 ? _GEN_846 : _GEN_3536; // @[i_cache.scala 86:34]
  wire  _GEN_3921 = unuse_way == 2'h1 ? _GEN_847 : _GEN_3537; // @[i_cache.scala 86:34]
  wire  _GEN_3922 = unuse_way == 2'h1 ? _GEN_848 : _GEN_3538; // @[i_cache.scala 86:34]
  wire  _GEN_3923 = unuse_way == 2'h1 ? _GEN_849 : _GEN_3539; // @[i_cache.scala 86:34]
  wire  _GEN_3924 = unuse_way == 2'h1 ? _GEN_850 : _GEN_3540; // @[i_cache.scala 86:34]
  wire  _GEN_3925 = unuse_way == 2'h1 ? _GEN_851 : _GEN_3541; // @[i_cache.scala 86:34]
  wire  _GEN_3926 = unuse_way == 2'h1 ? _GEN_852 : _GEN_3542; // @[i_cache.scala 86:34]
  wire  _GEN_3927 = unuse_way == 2'h1 ? _GEN_853 : _GEN_3543; // @[i_cache.scala 86:34]
  wire  _GEN_3928 = unuse_way == 2'h1 ? _GEN_854 : _GEN_3544; // @[i_cache.scala 86:34]
  wire  _GEN_3929 = unuse_way == 2'h1 ? _GEN_855 : _GEN_3545; // @[i_cache.scala 86:34]
  wire  _GEN_3930 = unuse_way == 2'h1 ? _GEN_856 : _GEN_3546; // @[i_cache.scala 86:34]
  wire  _GEN_3931 = unuse_way == 2'h1 ? _GEN_857 : _GEN_3547; // @[i_cache.scala 86:34]
  wire  _GEN_3932 = unuse_way == 2'h1 ? _GEN_858 : _GEN_3548; // @[i_cache.scala 86:34]
  wire  _GEN_3933 = unuse_way == 2'h1 ? _GEN_859 : _GEN_3549; // @[i_cache.scala 86:34]
  wire  _GEN_3934 = unuse_way == 2'h1 ? _GEN_860 : _GEN_3550; // @[i_cache.scala 86:34]
  wire  _GEN_3935 = unuse_way == 2'h1 ? _GEN_861 : _GEN_3551; // @[i_cache.scala 86:34]
  wire  _GEN_3936 = unuse_way == 2'h1 ? _GEN_862 : _GEN_3552; // @[i_cache.scala 86:34]
  wire  _GEN_3937 = unuse_way == 2'h1 ? _GEN_863 : _GEN_3553; // @[i_cache.scala 86:34]
  wire  _GEN_3938 = unuse_way == 2'h1 ? _GEN_864 : _GEN_3554; // @[i_cache.scala 86:34]
  wire  _GEN_3939 = unuse_way == 2'h1 ? _GEN_865 : _GEN_3555; // @[i_cache.scala 86:34]
  wire  _GEN_3940 = unuse_way == 2'h1 ? _GEN_866 : _GEN_3556; // @[i_cache.scala 86:34]
  wire  _GEN_3941 = unuse_way == 2'h1 ? _GEN_867 : _GEN_3557; // @[i_cache.scala 86:34]
  wire  _GEN_3942 = unuse_way == 2'h1 ? _GEN_868 : _GEN_3558; // @[i_cache.scala 86:34]
  wire  _GEN_3943 = unuse_way == 2'h1 ? _GEN_869 : _GEN_3559; // @[i_cache.scala 86:34]
  wire  _GEN_3944 = unuse_way == 2'h1 ? _GEN_870 : _GEN_3560; // @[i_cache.scala 86:34]
  wire  _GEN_3945 = unuse_way == 2'h1 ? _GEN_871 : _GEN_3561; // @[i_cache.scala 86:34]
  wire  _GEN_3946 = unuse_way == 2'h1 ? _GEN_872 : _GEN_3562; // @[i_cache.scala 86:34]
  wire  _GEN_3947 = unuse_way == 2'h1 ? _GEN_873 : _GEN_3563; // @[i_cache.scala 86:34]
  wire  _GEN_3948 = unuse_way == 2'h1 ? _GEN_874 : _GEN_3564; // @[i_cache.scala 86:34]
  wire  _GEN_3949 = unuse_way == 2'h1 ? _GEN_875 : _GEN_3565; // @[i_cache.scala 86:34]
  wire  _GEN_3950 = unuse_way == 2'h1 ? _GEN_876 : _GEN_3566; // @[i_cache.scala 86:34]
  wire  _GEN_3951 = unuse_way == 2'h1 ? _GEN_877 : _GEN_3567; // @[i_cache.scala 86:34]
  wire  _GEN_3952 = unuse_way == 2'h1 ? _GEN_878 : _GEN_3568; // @[i_cache.scala 86:34]
  wire  _GEN_3953 = unuse_way == 2'h1 ? _GEN_879 : _GEN_3569; // @[i_cache.scala 86:34]
  wire  _GEN_3954 = unuse_way == 2'h1 ? _GEN_880 : _GEN_3570; // @[i_cache.scala 86:34]
  wire  _GEN_3955 = unuse_way == 2'h1 ? _GEN_881 : _GEN_3571; // @[i_cache.scala 86:34]
  wire  _GEN_3956 = unuse_way == 2'h1 ? _GEN_882 : _GEN_3572; // @[i_cache.scala 86:34]
  wire  _GEN_3957 = unuse_way == 2'h1 ? _GEN_883 : _GEN_3573; // @[i_cache.scala 86:34]
  wire  _GEN_3958 = unuse_way == 2'h1 ? _GEN_884 : _GEN_3574; // @[i_cache.scala 86:34]
  wire  _GEN_3959 = unuse_way == 2'h1 ? _GEN_885 : _GEN_3575; // @[i_cache.scala 86:34]
  wire  _GEN_3960 = unuse_way == 2'h1 ? _GEN_886 : _GEN_3576; // @[i_cache.scala 86:34]
  wire  _GEN_3961 = unuse_way == 2'h1 ? _GEN_887 : _GEN_3577; // @[i_cache.scala 86:34]
  wire  _GEN_3962 = unuse_way == 2'h1 ? _GEN_888 : _GEN_3578; // @[i_cache.scala 86:34]
  wire  _GEN_3963 = unuse_way == 2'h1 ? _GEN_889 : _GEN_3579; // @[i_cache.scala 86:34]
  wire  _GEN_3964 = unuse_way == 2'h1 ? _GEN_890 : _GEN_3580; // @[i_cache.scala 86:34]
  wire  _GEN_3965 = unuse_way == 2'h1 ? _GEN_891 : _GEN_3581; // @[i_cache.scala 86:34]
  wire  _GEN_3966 = unuse_way == 2'h1 ? _GEN_892 : _GEN_3582; // @[i_cache.scala 86:34]
  wire  _GEN_3967 = unuse_way == 2'h1 ? _GEN_893 : _GEN_3583; // @[i_cache.scala 86:34]
  wire  _GEN_3968 = unuse_way == 2'h1 ? _GEN_894 : _GEN_3584; // @[i_cache.scala 86:34]
  wire  _GEN_3969 = unuse_way == 2'h1 ? _GEN_895 : _GEN_3585; // @[i_cache.scala 86:34]
  wire  _GEN_3970 = unuse_way == 2'h1 ? _GEN_896 : _GEN_3586; // @[i_cache.scala 86:34]
  wire  _GEN_3971 = unuse_way == 2'h1 ? _GEN_897 : _GEN_3587; // @[i_cache.scala 86:34]
  wire  _GEN_3972 = unuse_way == 2'h1 ? _GEN_898 : _GEN_3588; // @[i_cache.scala 86:34]
  wire  _GEN_3973 = unuse_way == 2'h1 ? _GEN_899 : _GEN_3589; // @[i_cache.scala 86:34]
  wire  _GEN_3974 = unuse_way == 2'h1 ? _GEN_900 : _GEN_3590; // @[i_cache.scala 86:34]
  wire  _GEN_3975 = unuse_way == 2'h1 ? _GEN_901 : _GEN_3591; // @[i_cache.scala 86:34]
  wire  _GEN_3976 = unuse_way == 2'h1 ? _GEN_902 : _GEN_3592; // @[i_cache.scala 86:34]
  wire  _GEN_3977 = unuse_way == 2'h1 ? _GEN_903 : _GEN_3593; // @[i_cache.scala 86:34]
  wire  _GEN_3978 = unuse_way == 2'h1 ? _GEN_904 : _GEN_3594; // @[i_cache.scala 86:34]
  wire  _GEN_3979 = unuse_way == 2'h1 ? _GEN_905 : _GEN_3595; // @[i_cache.scala 86:34]
  wire  _GEN_3980 = unuse_way == 2'h1 | _GEN_3211; // @[i_cache.scala 86:34 90:23]
  wire [63:0] _GEN_3981 = unuse_way == 2'h1 ? ram_1_0 : _GEN_2827; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3982 = unuse_way == 2'h1 ? ram_1_1 : _GEN_2828; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3983 = unuse_way == 2'h1 ? ram_1_2 : _GEN_2829; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3984 = unuse_way == 2'h1 ? ram_1_3 : _GEN_2830; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3985 = unuse_way == 2'h1 ? ram_1_4 : _GEN_2831; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3986 = unuse_way == 2'h1 ? ram_1_5 : _GEN_2832; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3987 = unuse_way == 2'h1 ? ram_1_6 : _GEN_2833; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3988 = unuse_way == 2'h1 ? ram_1_7 : _GEN_2834; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3989 = unuse_way == 2'h1 ? ram_1_8 : _GEN_2835; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3990 = unuse_way == 2'h1 ? ram_1_9 : _GEN_2836; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3991 = unuse_way == 2'h1 ? ram_1_10 : _GEN_2837; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3992 = unuse_way == 2'h1 ? ram_1_11 : _GEN_2838; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3993 = unuse_way == 2'h1 ? ram_1_12 : _GEN_2839; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3994 = unuse_way == 2'h1 ? ram_1_13 : _GEN_2840; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3995 = unuse_way == 2'h1 ? ram_1_14 : _GEN_2841; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3996 = unuse_way == 2'h1 ? ram_1_15 : _GEN_2842; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3997 = unuse_way == 2'h1 ? ram_1_16 : _GEN_2843; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3998 = unuse_way == 2'h1 ? ram_1_17 : _GEN_2844; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3999 = unuse_way == 2'h1 ? ram_1_18 : _GEN_2845; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4000 = unuse_way == 2'h1 ? ram_1_19 : _GEN_2846; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4001 = unuse_way == 2'h1 ? ram_1_20 : _GEN_2847; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4002 = unuse_way == 2'h1 ? ram_1_21 : _GEN_2848; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4003 = unuse_way == 2'h1 ? ram_1_22 : _GEN_2849; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4004 = unuse_way == 2'h1 ? ram_1_23 : _GEN_2850; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4005 = unuse_way == 2'h1 ? ram_1_24 : _GEN_2851; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4006 = unuse_way == 2'h1 ? ram_1_25 : _GEN_2852; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4007 = unuse_way == 2'h1 ? ram_1_26 : _GEN_2853; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4008 = unuse_way == 2'h1 ? ram_1_27 : _GEN_2854; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4009 = unuse_way == 2'h1 ? ram_1_28 : _GEN_2855; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4010 = unuse_way == 2'h1 ? ram_1_29 : _GEN_2856; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4011 = unuse_way == 2'h1 ? ram_1_30 : _GEN_2857; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4012 = unuse_way == 2'h1 ? ram_1_31 : _GEN_2858; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4013 = unuse_way == 2'h1 ? ram_1_32 : _GEN_2859; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4014 = unuse_way == 2'h1 ? ram_1_33 : _GEN_2860; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4015 = unuse_way == 2'h1 ? ram_1_34 : _GEN_2861; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4016 = unuse_way == 2'h1 ? ram_1_35 : _GEN_2862; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4017 = unuse_way == 2'h1 ? ram_1_36 : _GEN_2863; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4018 = unuse_way == 2'h1 ? ram_1_37 : _GEN_2864; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4019 = unuse_way == 2'h1 ? ram_1_38 : _GEN_2865; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4020 = unuse_way == 2'h1 ? ram_1_39 : _GEN_2866; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4021 = unuse_way == 2'h1 ? ram_1_40 : _GEN_2867; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4022 = unuse_way == 2'h1 ? ram_1_41 : _GEN_2868; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4023 = unuse_way == 2'h1 ? ram_1_42 : _GEN_2869; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4024 = unuse_way == 2'h1 ? ram_1_43 : _GEN_2870; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4025 = unuse_way == 2'h1 ? ram_1_44 : _GEN_2871; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4026 = unuse_way == 2'h1 ? ram_1_45 : _GEN_2872; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4027 = unuse_way == 2'h1 ? ram_1_46 : _GEN_2873; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4028 = unuse_way == 2'h1 ? ram_1_47 : _GEN_2874; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4029 = unuse_way == 2'h1 ? ram_1_48 : _GEN_2875; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4030 = unuse_way == 2'h1 ? ram_1_49 : _GEN_2876; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4031 = unuse_way == 2'h1 ? ram_1_50 : _GEN_2877; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4032 = unuse_way == 2'h1 ? ram_1_51 : _GEN_2878; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4033 = unuse_way == 2'h1 ? ram_1_52 : _GEN_2879; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4034 = unuse_way == 2'h1 ? ram_1_53 : _GEN_2880; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4035 = unuse_way == 2'h1 ? ram_1_54 : _GEN_2881; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4036 = unuse_way == 2'h1 ? ram_1_55 : _GEN_2882; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4037 = unuse_way == 2'h1 ? ram_1_56 : _GEN_2883; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4038 = unuse_way == 2'h1 ? ram_1_57 : _GEN_2884; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4039 = unuse_way == 2'h1 ? ram_1_58 : _GEN_2885; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4040 = unuse_way == 2'h1 ? ram_1_59 : _GEN_2886; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4041 = unuse_way == 2'h1 ? ram_1_60 : _GEN_2887; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4042 = unuse_way == 2'h1 ? ram_1_61 : _GEN_2888; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4043 = unuse_way == 2'h1 ? ram_1_62 : _GEN_2889; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4044 = unuse_way == 2'h1 ? ram_1_63 : _GEN_2890; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4045 = unuse_way == 2'h1 ? ram_1_64 : _GEN_2891; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4046 = unuse_way == 2'h1 ? ram_1_65 : _GEN_2892; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4047 = unuse_way == 2'h1 ? ram_1_66 : _GEN_2893; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4048 = unuse_way == 2'h1 ? ram_1_67 : _GEN_2894; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4049 = unuse_way == 2'h1 ? ram_1_68 : _GEN_2895; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4050 = unuse_way == 2'h1 ? ram_1_69 : _GEN_2896; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4051 = unuse_way == 2'h1 ? ram_1_70 : _GEN_2897; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4052 = unuse_way == 2'h1 ? ram_1_71 : _GEN_2898; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4053 = unuse_way == 2'h1 ? ram_1_72 : _GEN_2899; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4054 = unuse_way == 2'h1 ? ram_1_73 : _GEN_2900; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4055 = unuse_way == 2'h1 ? ram_1_74 : _GEN_2901; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4056 = unuse_way == 2'h1 ? ram_1_75 : _GEN_2902; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4057 = unuse_way == 2'h1 ? ram_1_76 : _GEN_2903; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4058 = unuse_way == 2'h1 ? ram_1_77 : _GEN_2904; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4059 = unuse_way == 2'h1 ? ram_1_78 : _GEN_2905; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4060 = unuse_way == 2'h1 ? ram_1_79 : _GEN_2906; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4061 = unuse_way == 2'h1 ? ram_1_80 : _GEN_2907; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4062 = unuse_way == 2'h1 ? ram_1_81 : _GEN_2908; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4063 = unuse_way == 2'h1 ? ram_1_82 : _GEN_2909; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4064 = unuse_way == 2'h1 ? ram_1_83 : _GEN_2910; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4065 = unuse_way == 2'h1 ? ram_1_84 : _GEN_2911; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4066 = unuse_way == 2'h1 ? ram_1_85 : _GEN_2912; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4067 = unuse_way == 2'h1 ? ram_1_86 : _GEN_2913; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4068 = unuse_way == 2'h1 ? ram_1_87 : _GEN_2914; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4069 = unuse_way == 2'h1 ? ram_1_88 : _GEN_2915; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4070 = unuse_way == 2'h1 ? ram_1_89 : _GEN_2916; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4071 = unuse_way == 2'h1 ? ram_1_90 : _GEN_2917; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4072 = unuse_way == 2'h1 ? ram_1_91 : _GEN_2918; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4073 = unuse_way == 2'h1 ? ram_1_92 : _GEN_2919; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4074 = unuse_way == 2'h1 ? ram_1_93 : _GEN_2920; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4075 = unuse_way == 2'h1 ? ram_1_94 : _GEN_2921; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4076 = unuse_way == 2'h1 ? ram_1_95 : _GEN_2922; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4077 = unuse_way == 2'h1 ? ram_1_96 : _GEN_2923; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4078 = unuse_way == 2'h1 ? ram_1_97 : _GEN_2924; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4079 = unuse_way == 2'h1 ? ram_1_98 : _GEN_2925; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4080 = unuse_way == 2'h1 ? ram_1_99 : _GEN_2926; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4081 = unuse_way == 2'h1 ? ram_1_100 : _GEN_2927; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4082 = unuse_way == 2'h1 ? ram_1_101 : _GEN_2928; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4083 = unuse_way == 2'h1 ? ram_1_102 : _GEN_2929; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4084 = unuse_way == 2'h1 ? ram_1_103 : _GEN_2930; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4085 = unuse_way == 2'h1 ? ram_1_104 : _GEN_2931; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4086 = unuse_way == 2'h1 ? ram_1_105 : _GEN_2932; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4087 = unuse_way == 2'h1 ? ram_1_106 : _GEN_2933; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4088 = unuse_way == 2'h1 ? ram_1_107 : _GEN_2934; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4089 = unuse_way == 2'h1 ? ram_1_108 : _GEN_2935; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4090 = unuse_way == 2'h1 ? ram_1_109 : _GEN_2936; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4091 = unuse_way == 2'h1 ? ram_1_110 : _GEN_2937; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4092 = unuse_way == 2'h1 ? ram_1_111 : _GEN_2938; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4093 = unuse_way == 2'h1 ? ram_1_112 : _GEN_2939; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4094 = unuse_way == 2'h1 ? ram_1_113 : _GEN_2940; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4095 = unuse_way == 2'h1 ? ram_1_114 : _GEN_2941; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4096 = unuse_way == 2'h1 ? ram_1_115 : _GEN_2942; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4097 = unuse_way == 2'h1 ? ram_1_116 : _GEN_2943; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4098 = unuse_way == 2'h1 ? ram_1_117 : _GEN_2944; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4099 = unuse_way == 2'h1 ? ram_1_118 : _GEN_2945; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4100 = unuse_way == 2'h1 ? ram_1_119 : _GEN_2946; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4101 = unuse_way == 2'h1 ? ram_1_120 : _GEN_2947; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4102 = unuse_way == 2'h1 ? ram_1_121 : _GEN_2948; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4103 = unuse_way == 2'h1 ? ram_1_122 : _GEN_2949; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4104 = unuse_way == 2'h1 ? ram_1_123 : _GEN_2950; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4105 = unuse_way == 2'h1 ? ram_1_124 : _GEN_2951; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4106 = unuse_way == 2'h1 ? ram_1_125 : _GEN_2952; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4107 = unuse_way == 2'h1 ? ram_1_126 : _GEN_2953; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4108 = unuse_way == 2'h1 ? ram_1_127 : _GEN_2954; // @[i_cache.scala 18:24 86:34]
  wire [31:0] _GEN_4109 = unuse_way == 2'h1 ? tag_1_0 : _GEN_2955; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4110 = unuse_way == 2'h1 ? tag_1_1 : _GEN_2956; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4111 = unuse_way == 2'h1 ? tag_1_2 : _GEN_2957; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4112 = unuse_way == 2'h1 ? tag_1_3 : _GEN_2958; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4113 = unuse_way == 2'h1 ? tag_1_4 : _GEN_2959; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4114 = unuse_way == 2'h1 ? tag_1_5 : _GEN_2960; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4115 = unuse_way == 2'h1 ? tag_1_6 : _GEN_2961; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4116 = unuse_way == 2'h1 ? tag_1_7 : _GEN_2962; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4117 = unuse_way == 2'h1 ? tag_1_8 : _GEN_2963; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4118 = unuse_way == 2'h1 ? tag_1_9 : _GEN_2964; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4119 = unuse_way == 2'h1 ? tag_1_10 : _GEN_2965; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4120 = unuse_way == 2'h1 ? tag_1_11 : _GEN_2966; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4121 = unuse_way == 2'h1 ? tag_1_12 : _GEN_2967; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4122 = unuse_way == 2'h1 ? tag_1_13 : _GEN_2968; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4123 = unuse_way == 2'h1 ? tag_1_14 : _GEN_2969; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4124 = unuse_way == 2'h1 ? tag_1_15 : _GEN_2970; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4125 = unuse_way == 2'h1 ? tag_1_16 : _GEN_2971; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4126 = unuse_way == 2'h1 ? tag_1_17 : _GEN_2972; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4127 = unuse_way == 2'h1 ? tag_1_18 : _GEN_2973; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4128 = unuse_way == 2'h1 ? tag_1_19 : _GEN_2974; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4129 = unuse_way == 2'h1 ? tag_1_20 : _GEN_2975; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4130 = unuse_way == 2'h1 ? tag_1_21 : _GEN_2976; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4131 = unuse_way == 2'h1 ? tag_1_22 : _GEN_2977; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4132 = unuse_way == 2'h1 ? tag_1_23 : _GEN_2978; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4133 = unuse_way == 2'h1 ? tag_1_24 : _GEN_2979; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4134 = unuse_way == 2'h1 ? tag_1_25 : _GEN_2980; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4135 = unuse_way == 2'h1 ? tag_1_26 : _GEN_2981; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4136 = unuse_way == 2'h1 ? tag_1_27 : _GEN_2982; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4137 = unuse_way == 2'h1 ? tag_1_28 : _GEN_2983; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4138 = unuse_way == 2'h1 ? tag_1_29 : _GEN_2984; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4139 = unuse_way == 2'h1 ? tag_1_30 : _GEN_2985; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4140 = unuse_way == 2'h1 ? tag_1_31 : _GEN_2986; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4141 = unuse_way == 2'h1 ? tag_1_32 : _GEN_2987; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4142 = unuse_way == 2'h1 ? tag_1_33 : _GEN_2988; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4143 = unuse_way == 2'h1 ? tag_1_34 : _GEN_2989; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4144 = unuse_way == 2'h1 ? tag_1_35 : _GEN_2990; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4145 = unuse_way == 2'h1 ? tag_1_36 : _GEN_2991; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4146 = unuse_way == 2'h1 ? tag_1_37 : _GEN_2992; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4147 = unuse_way == 2'h1 ? tag_1_38 : _GEN_2993; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4148 = unuse_way == 2'h1 ? tag_1_39 : _GEN_2994; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4149 = unuse_way == 2'h1 ? tag_1_40 : _GEN_2995; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4150 = unuse_way == 2'h1 ? tag_1_41 : _GEN_2996; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4151 = unuse_way == 2'h1 ? tag_1_42 : _GEN_2997; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4152 = unuse_way == 2'h1 ? tag_1_43 : _GEN_2998; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4153 = unuse_way == 2'h1 ? tag_1_44 : _GEN_2999; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4154 = unuse_way == 2'h1 ? tag_1_45 : _GEN_3000; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4155 = unuse_way == 2'h1 ? tag_1_46 : _GEN_3001; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4156 = unuse_way == 2'h1 ? tag_1_47 : _GEN_3002; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4157 = unuse_way == 2'h1 ? tag_1_48 : _GEN_3003; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4158 = unuse_way == 2'h1 ? tag_1_49 : _GEN_3004; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4159 = unuse_way == 2'h1 ? tag_1_50 : _GEN_3005; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4160 = unuse_way == 2'h1 ? tag_1_51 : _GEN_3006; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4161 = unuse_way == 2'h1 ? tag_1_52 : _GEN_3007; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4162 = unuse_way == 2'h1 ? tag_1_53 : _GEN_3008; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4163 = unuse_way == 2'h1 ? tag_1_54 : _GEN_3009; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4164 = unuse_way == 2'h1 ? tag_1_55 : _GEN_3010; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4165 = unuse_way == 2'h1 ? tag_1_56 : _GEN_3011; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4166 = unuse_way == 2'h1 ? tag_1_57 : _GEN_3012; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4167 = unuse_way == 2'h1 ? tag_1_58 : _GEN_3013; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4168 = unuse_way == 2'h1 ? tag_1_59 : _GEN_3014; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4169 = unuse_way == 2'h1 ? tag_1_60 : _GEN_3015; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4170 = unuse_way == 2'h1 ? tag_1_61 : _GEN_3016; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4171 = unuse_way == 2'h1 ? tag_1_62 : _GEN_3017; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4172 = unuse_way == 2'h1 ? tag_1_63 : _GEN_3018; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4173 = unuse_way == 2'h1 ? tag_1_64 : _GEN_3019; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4174 = unuse_way == 2'h1 ? tag_1_65 : _GEN_3020; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4175 = unuse_way == 2'h1 ? tag_1_66 : _GEN_3021; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4176 = unuse_way == 2'h1 ? tag_1_67 : _GEN_3022; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4177 = unuse_way == 2'h1 ? tag_1_68 : _GEN_3023; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4178 = unuse_way == 2'h1 ? tag_1_69 : _GEN_3024; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4179 = unuse_way == 2'h1 ? tag_1_70 : _GEN_3025; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4180 = unuse_way == 2'h1 ? tag_1_71 : _GEN_3026; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4181 = unuse_way == 2'h1 ? tag_1_72 : _GEN_3027; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4182 = unuse_way == 2'h1 ? tag_1_73 : _GEN_3028; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4183 = unuse_way == 2'h1 ? tag_1_74 : _GEN_3029; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4184 = unuse_way == 2'h1 ? tag_1_75 : _GEN_3030; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4185 = unuse_way == 2'h1 ? tag_1_76 : _GEN_3031; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4186 = unuse_way == 2'h1 ? tag_1_77 : _GEN_3032; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4187 = unuse_way == 2'h1 ? tag_1_78 : _GEN_3033; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4188 = unuse_way == 2'h1 ? tag_1_79 : _GEN_3034; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4189 = unuse_way == 2'h1 ? tag_1_80 : _GEN_3035; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4190 = unuse_way == 2'h1 ? tag_1_81 : _GEN_3036; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4191 = unuse_way == 2'h1 ? tag_1_82 : _GEN_3037; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4192 = unuse_way == 2'h1 ? tag_1_83 : _GEN_3038; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4193 = unuse_way == 2'h1 ? tag_1_84 : _GEN_3039; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4194 = unuse_way == 2'h1 ? tag_1_85 : _GEN_3040; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4195 = unuse_way == 2'h1 ? tag_1_86 : _GEN_3041; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4196 = unuse_way == 2'h1 ? tag_1_87 : _GEN_3042; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4197 = unuse_way == 2'h1 ? tag_1_88 : _GEN_3043; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4198 = unuse_way == 2'h1 ? tag_1_89 : _GEN_3044; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4199 = unuse_way == 2'h1 ? tag_1_90 : _GEN_3045; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4200 = unuse_way == 2'h1 ? tag_1_91 : _GEN_3046; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4201 = unuse_way == 2'h1 ? tag_1_92 : _GEN_3047; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4202 = unuse_way == 2'h1 ? tag_1_93 : _GEN_3048; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4203 = unuse_way == 2'h1 ? tag_1_94 : _GEN_3049; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4204 = unuse_way == 2'h1 ? tag_1_95 : _GEN_3050; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4205 = unuse_way == 2'h1 ? tag_1_96 : _GEN_3051; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4206 = unuse_way == 2'h1 ? tag_1_97 : _GEN_3052; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4207 = unuse_way == 2'h1 ? tag_1_98 : _GEN_3053; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4208 = unuse_way == 2'h1 ? tag_1_99 : _GEN_3054; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4209 = unuse_way == 2'h1 ? tag_1_100 : _GEN_3055; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4210 = unuse_way == 2'h1 ? tag_1_101 : _GEN_3056; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4211 = unuse_way == 2'h1 ? tag_1_102 : _GEN_3057; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4212 = unuse_way == 2'h1 ? tag_1_103 : _GEN_3058; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4213 = unuse_way == 2'h1 ? tag_1_104 : _GEN_3059; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4214 = unuse_way == 2'h1 ? tag_1_105 : _GEN_3060; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4215 = unuse_way == 2'h1 ? tag_1_106 : _GEN_3061; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4216 = unuse_way == 2'h1 ? tag_1_107 : _GEN_3062; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4217 = unuse_way == 2'h1 ? tag_1_108 : _GEN_3063; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4218 = unuse_way == 2'h1 ? tag_1_109 : _GEN_3064; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4219 = unuse_way == 2'h1 ? tag_1_110 : _GEN_3065; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4220 = unuse_way == 2'h1 ? tag_1_111 : _GEN_3066; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4221 = unuse_way == 2'h1 ? tag_1_112 : _GEN_3067; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4222 = unuse_way == 2'h1 ? tag_1_113 : _GEN_3068; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4223 = unuse_way == 2'h1 ? tag_1_114 : _GEN_3069; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4224 = unuse_way == 2'h1 ? tag_1_115 : _GEN_3070; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4225 = unuse_way == 2'h1 ? tag_1_116 : _GEN_3071; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4226 = unuse_way == 2'h1 ? tag_1_117 : _GEN_3072; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4227 = unuse_way == 2'h1 ? tag_1_118 : _GEN_3073; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4228 = unuse_way == 2'h1 ? tag_1_119 : _GEN_3074; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4229 = unuse_way == 2'h1 ? tag_1_120 : _GEN_3075; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4230 = unuse_way == 2'h1 ? tag_1_121 : _GEN_3076; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4231 = unuse_way == 2'h1 ? tag_1_122 : _GEN_3077; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4232 = unuse_way == 2'h1 ? tag_1_123 : _GEN_3078; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4233 = unuse_way == 2'h1 ? tag_1_124 : _GEN_3079; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4234 = unuse_way == 2'h1 ? tag_1_125 : _GEN_3080; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4235 = unuse_way == 2'h1 ? tag_1_126 : _GEN_3081; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4236 = unuse_way == 2'h1 ? tag_1_127 : _GEN_3082; // @[i_cache.scala 20:24 86:34]
  wire  _GEN_4237 = unuse_way == 2'h1 ? valid_1_0 : _GEN_3083; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4238 = unuse_way == 2'h1 ? valid_1_1 : _GEN_3084; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4239 = unuse_way == 2'h1 ? valid_1_2 : _GEN_3085; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4240 = unuse_way == 2'h1 ? valid_1_3 : _GEN_3086; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4241 = unuse_way == 2'h1 ? valid_1_4 : _GEN_3087; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4242 = unuse_way == 2'h1 ? valid_1_5 : _GEN_3088; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4243 = unuse_way == 2'h1 ? valid_1_6 : _GEN_3089; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4244 = unuse_way == 2'h1 ? valid_1_7 : _GEN_3090; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4245 = unuse_way == 2'h1 ? valid_1_8 : _GEN_3091; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4246 = unuse_way == 2'h1 ? valid_1_9 : _GEN_3092; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4247 = unuse_way == 2'h1 ? valid_1_10 : _GEN_3093; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4248 = unuse_way == 2'h1 ? valid_1_11 : _GEN_3094; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4249 = unuse_way == 2'h1 ? valid_1_12 : _GEN_3095; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4250 = unuse_way == 2'h1 ? valid_1_13 : _GEN_3096; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4251 = unuse_way == 2'h1 ? valid_1_14 : _GEN_3097; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4252 = unuse_way == 2'h1 ? valid_1_15 : _GEN_3098; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4253 = unuse_way == 2'h1 ? valid_1_16 : _GEN_3099; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4254 = unuse_way == 2'h1 ? valid_1_17 : _GEN_3100; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4255 = unuse_way == 2'h1 ? valid_1_18 : _GEN_3101; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4256 = unuse_way == 2'h1 ? valid_1_19 : _GEN_3102; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4257 = unuse_way == 2'h1 ? valid_1_20 : _GEN_3103; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4258 = unuse_way == 2'h1 ? valid_1_21 : _GEN_3104; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4259 = unuse_way == 2'h1 ? valid_1_22 : _GEN_3105; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4260 = unuse_way == 2'h1 ? valid_1_23 : _GEN_3106; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4261 = unuse_way == 2'h1 ? valid_1_24 : _GEN_3107; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4262 = unuse_way == 2'h1 ? valid_1_25 : _GEN_3108; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4263 = unuse_way == 2'h1 ? valid_1_26 : _GEN_3109; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4264 = unuse_way == 2'h1 ? valid_1_27 : _GEN_3110; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4265 = unuse_way == 2'h1 ? valid_1_28 : _GEN_3111; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4266 = unuse_way == 2'h1 ? valid_1_29 : _GEN_3112; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4267 = unuse_way == 2'h1 ? valid_1_30 : _GEN_3113; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4268 = unuse_way == 2'h1 ? valid_1_31 : _GEN_3114; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4269 = unuse_way == 2'h1 ? valid_1_32 : _GEN_3115; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4270 = unuse_way == 2'h1 ? valid_1_33 : _GEN_3116; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4271 = unuse_way == 2'h1 ? valid_1_34 : _GEN_3117; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4272 = unuse_way == 2'h1 ? valid_1_35 : _GEN_3118; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4273 = unuse_way == 2'h1 ? valid_1_36 : _GEN_3119; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4274 = unuse_way == 2'h1 ? valid_1_37 : _GEN_3120; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4275 = unuse_way == 2'h1 ? valid_1_38 : _GEN_3121; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4276 = unuse_way == 2'h1 ? valid_1_39 : _GEN_3122; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4277 = unuse_way == 2'h1 ? valid_1_40 : _GEN_3123; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4278 = unuse_way == 2'h1 ? valid_1_41 : _GEN_3124; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4279 = unuse_way == 2'h1 ? valid_1_42 : _GEN_3125; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4280 = unuse_way == 2'h1 ? valid_1_43 : _GEN_3126; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4281 = unuse_way == 2'h1 ? valid_1_44 : _GEN_3127; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4282 = unuse_way == 2'h1 ? valid_1_45 : _GEN_3128; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4283 = unuse_way == 2'h1 ? valid_1_46 : _GEN_3129; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4284 = unuse_way == 2'h1 ? valid_1_47 : _GEN_3130; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4285 = unuse_way == 2'h1 ? valid_1_48 : _GEN_3131; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4286 = unuse_way == 2'h1 ? valid_1_49 : _GEN_3132; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4287 = unuse_way == 2'h1 ? valid_1_50 : _GEN_3133; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4288 = unuse_way == 2'h1 ? valid_1_51 : _GEN_3134; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4289 = unuse_way == 2'h1 ? valid_1_52 : _GEN_3135; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4290 = unuse_way == 2'h1 ? valid_1_53 : _GEN_3136; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4291 = unuse_way == 2'h1 ? valid_1_54 : _GEN_3137; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4292 = unuse_way == 2'h1 ? valid_1_55 : _GEN_3138; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4293 = unuse_way == 2'h1 ? valid_1_56 : _GEN_3139; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4294 = unuse_way == 2'h1 ? valid_1_57 : _GEN_3140; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4295 = unuse_way == 2'h1 ? valid_1_58 : _GEN_3141; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4296 = unuse_way == 2'h1 ? valid_1_59 : _GEN_3142; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4297 = unuse_way == 2'h1 ? valid_1_60 : _GEN_3143; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4298 = unuse_way == 2'h1 ? valid_1_61 : _GEN_3144; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4299 = unuse_way == 2'h1 ? valid_1_62 : _GEN_3145; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4300 = unuse_way == 2'h1 ? valid_1_63 : _GEN_3146; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4301 = unuse_way == 2'h1 ? valid_1_64 : _GEN_3147; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4302 = unuse_way == 2'h1 ? valid_1_65 : _GEN_3148; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4303 = unuse_way == 2'h1 ? valid_1_66 : _GEN_3149; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4304 = unuse_way == 2'h1 ? valid_1_67 : _GEN_3150; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4305 = unuse_way == 2'h1 ? valid_1_68 : _GEN_3151; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4306 = unuse_way == 2'h1 ? valid_1_69 : _GEN_3152; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4307 = unuse_way == 2'h1 ? valid_1_70 : _GEN_3153; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4308 = unuse_way == 2'h1 ? valid_1_71 : _GEN_3154; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4309 = unuse_way == 2'h1 ? valid_1_72 : _GEN_3155; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4310 = unuse_way == 2'h1 ? valid_1_73 : _GEN_3156; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4311 = unuse_way == 2'h1 ? valid_1_74 : _GEN_3157; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4312 = unuse_way == 2'h1 ? valid_1_75 : _GEN_3158; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4313 = unuse_way == 2'h1 ? valid_1_76 : _GEN_3159; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4314 = unuse_way == 2'h1 ? valid_1_77 : _GEN_3160; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4315 = unuse_way == 2'h1 ? valid_1_78 : _GEN_3161; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4316 = unuse_way == 2'h1 ? valid_1_79 : _GEN_3162; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4317 = unuse_way == 2'h1 ? valid_1_80 : _GEN_3163; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4318 = unuse_way == 2'h1 ? valid_1_81 : _GEN_3164; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4319 = unuse_way == 2'h1 ? valid_1_82 : _GEN_3165; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4320 = unuse_way == 2'h1 ? valid_1_83 : _GEN_3166; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4321 = unuse_way == 2'h1 ? valid_1_84 : _GEN_3167; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4322 = unuse_way == 2'h1 ? valid_1_85 : _GEN_3168; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4323 = unuse_way == 2'h1 ? valid_1_86 : _GEN_3169; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4324 = unuse_way == 2'h1 ? valid_1_87 : _GEN_3170; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4325 = unuse_way == 2'h1 ? valid_1_88 : _GEN_3171; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4326 = unuse_way == 2'h1 ? valid_1_89 : _GEN_3172; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4327 = unuse_way == 2'h1 ? valid_1_90 : _GEN_3173; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4328 = unuse_way == 2'h1 ? valid_1_91 : _GEN_3174; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4329 = unuse_way == 2'h1 ? valid_1_92 : _GEN_3175; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4330 = unuse_way == 2'h1 ? valid_1_93 : _GEN_3176; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4331 = unuse_way == 2'h1 ? valid_1_94 : _GEN_3177; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4332 = unuse_way == 2'h1 ? valid_1_95 : _GEN_3178; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4333 = unuse_way == 2'h1 ? valid_1_96 : _GEN_3179; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4334 = unuse_way == 2'h1 ? valid_1_97 : _GEN_3180; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4335 = unuse_way == 2'h1 ? valid_1_98 : _GEN_3181; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4336 = unuse_way == 2'h1 ? valid_1_99 : _GEN_3182; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4337 = unuse_way == 2'h1 ? valid_1_100 : _GEN_3183; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4338 = unuse_way == 2'h1 ? valid_1_101 : _GEN_3184; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4339 = unuse_way == 2'h1 ? valid_1_102 : _GEN_3185; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4340 = unuse_way == 2'h1 ? valid_1_103 : _GEN_3186; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4341 = unuse_way == 2'h1 ? valid_1_104 : _GEN_3187; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4342 = unuse_way == 2'h1 ? valid_1_105 : _GEN_3188; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4343 = unuse_way == 2'h1 ? valid_1_106 : _GEN_3189; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4344 = unuse_way == 2'h1 ? valid_1_107 : _GEN_3190; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4345 = unuse_way == 2'h1 ? valid_1_108 : _GEN_3191; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4346 = unuse_way == 2'h1 ? valid_1_109 : _GEN_3192; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4347 = unuse_way == 2'h1 ? valid_1_110 : _GEN_3193; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4348 = unuse_way == 2'h1 ? valid_1_111 : _GEN_3194; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4349 = unuse_way == 2'h1 ? valid_1_112 : _GEN_3195; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4350 = unuse_way == 2'h1 ? valid_1_113 : _GEN_3196; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4351 = unuse_way == 2'h1 ? valid_1_114 : _GEN_3197; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4352 = unuse_way == 2'h1 ? valid_1_115 : _GEN_3198; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4353 = unuse_way == 2'h1 ? valid_1_116 : _GEN_3199; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4354 = unuse_way == 2'h1 ? valid_1_117 : _GEN_3200; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4355 = unuse_way == 2'h1 ? valid_1_118 : _GEN_3201; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4356 = unuse_way == 2'h1 ? valid_1_119 : _GEN_3202; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4357 = unuse_way == 2'h1 ? valid_1_120 : _GEN_3203; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4358 = unuse_way == 2'h1 ? valid_1_121 : _GEN_3204; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4359 = unuse_way == 2'h1 ? valid_1_122 : _GEN_3205; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4360 = unuse_way == 2'h1 ? valid_1_123 : _GEN_3206; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4361 = unuse_way == 2'h1 ? valid_1_124 : _GEN_3207; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4362 = unuse_way == 2'h1 ? valid_1_125 : _GEN_3208; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4363 = unuse_way == 2'h1 ? valid_1_126 : _GEN_3209; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4364 = unuse_way == 2'h1 ? valid_1_127 : _GEN_3210; // @[i_cache.scala 22:26 86:34]
  wire [2:0] _GEN_4365 = 3'h4 == state ? 3'h1 : state; // @[i_cache.scala 55:18 111:19 53:24]
  wire [2:0] _GEN_4366 = 3'h3 == state ? 3'h4 : _GEN_4365; // @[i_cache.scala 55:18 85:19]
  wire [63:0] _GEN_4367 = 3'h3 == state ? _GEN_3596 : ram_0_0; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4368 = 3'h3 == state ? _GEN_3597 : ram_0_1; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4369 = 3'h3 == state ? _GEN_3598 : ram_0_2; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4370 = 3'h3 == state ? _GEN_3599 : ram_0_3; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4371 = 3'h3 == state ? _GEN_3600 : ram_0_4; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4372 = 3'h3 == state ? _GEN_3601 : ram_0_5; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4373 = 3'h3 == state ? _GEN_3602 : ram_0_6; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4374 = 3'h3 == state ? _GEN_3603 : ram_0_7; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4375 = 3'h3 == state ? _GEN_3604 : ram_0_8; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4376 = 3'h3 == state ? _GEN_3605 : ram_0_9; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4377 = 3'h3 == state ? _GEN_3606 : ram_0_10; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4378 = 3'h3 == state ? _GEN_3607 : ram_0_11; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4379 = 3'h3 == state ? _GEN_3608 : ram_0_12; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4380 = 3'h3 == state ? _GEN_3609 : ram_0_13; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4381 = 3'h3 == state ? _GEN_3610 : ram_0_14; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4382 = 3'h3 == state ? _GEN_3611 : ram_0_15; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4383 = 3'h3 == state ? _GEN_3612 : ram_0_16; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4384 = 3'h3 == state ? _GEN_3613 : ram_0_17; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4385 = 3'h3 == state ? _GEN_3614 : ram_0_18; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4386 = 3'h3 == state ? _GEN_3615 : ram_0_19; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4387 = 3'h3 == state ? _GEN_3616 : ram_0_20; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4388 = 3'h3 == state ? _GEN_3617 : ram_0_21; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4389 = 3'h3 == state ? _GEN_3618 : ram_0_22; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4390 = 3'h3 == state ? _GEN_3619 : ram_0_23; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4391 = 3'h3 == state ? _GEN_3620 : ram_0_24; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4392 = 3'h3 == state ? _GEN_3621 : ram_0_25; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4393 = 3'h3 == state ? _GEN_3622 : ram_0_26; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4394 = 3'h3 == state ? _GEN_3623 : ram_0_27; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4395 = 3'h3 == state ? _GEN_3624 : ram_0_28; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4396 = 3'h3 == state ? _GEN_3625 : ram_0_29; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4397 = 3'h3 == state ? _GEN_3626 : ram_0_30; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4398 = 3'h3 == state ? _GEN_3627 : ram_0_31; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4399 = 3'h3 == state ? _GEN_3628 : ram_0_32; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4400 = 3'h3 == state ? _GEN_3629 : ram_0_33; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4401 = 3'h3 == state ? _GEN_3630 : ram_0_34; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4402 = 3'h3 == state ? _GEN_3631 : ram_0_35; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4403 = 3'h3 == state ? _GEN_3632 : ram_0_36; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4404 = 3'h3 == state ? _GEN_3633 : ram_0_37; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4405 = 3'h3 == state ? _GEN_3634 : ram_0_38; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4406 = 3'h3 == state ? _GEN_3635 : ram_0_39; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4407 = 3'h3 == state ? _GEN_3636 : ram_0_40; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4408 = 3'h3 == state ? _GEN_3637 : ram_0_41; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4409 = 3'h3 == state ? _GEN_3638 : ram_0_42; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4410 = 3'h3 == state ? _GEN_3639 : ram_0_43; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4411 = 3'h3 == state ? _GEN_3640 : ram_0_44; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4412 = 3'h3 == state ? _GEN_3641 : ram_0_45; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4413 = 3'h3 == state ? _GEN_3642 : ram_0_46; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4414 = 3'h3 == state ? _GEN_3643 : ram_0_47; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4415 = 3'h3 == state ? _GEN_3644 : ram_0_48; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4416 = 3'h3 == state ? _GEN_3645 : ram_0_49; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4417 = 3'h3 == state ? _GEN_3646 : ram_0_50; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4418 = 3'h3 == state ? _GEN_3647 : ram_0_51; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4419 = 3'h3 == state ? _GEN_3648 : ram_0_52; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4420 = 3'h3 == state ? _GEN_3649 : ram_0_53; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4421 = 3'h3 == state ? _GEN_3650 : ram_0_54; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4422 = 3'h3 == state ? _GEN_3651 : ram_0_55; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4423 = 3'h3 == state ? _GEN_3652 : ram_0_56; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4424 = 3'h3 == state ? _GEN_3653 : ram_0_57; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4425 = 3'h3 == state ? _GEN_3654 : ram_0_58; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4426 = 3'h3 == state ? _GEN_3655 : ram_0_59; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4427 = 3'h3 == state ? _GEN_3656 : ram_0_60; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4428 = 3'h3 == state ? _GEN_3657 : ram_0_61; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4429 = 3'h3 == state ? _GEN_3658 : ram_0_62; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4430 = 3'h3 == state ? _GEN_3659 : ram_0_63; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4431 = 3'h3 == state ? _GEN_3660 : ram_0_64; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4432 = 3'h3 == state ? _GEN_3661 : ram_0_65; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4433 = 3'h3 == state ? _GEN_3662 : ram_0_66; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4434 = 3'h3 == state ? _GEN_3663 : ram_0_67; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4435 = 3'h3 == state ? _GEN_3664 : ram_0_68; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4436 = 3'h3 == state ? _GEN_3665 : ram_0_69; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4437 = 3'h3 == state ? _GEN_3666 : ram_0_70; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4438 = 3'h3 == state ? _GEN_3667 : ram_0_71; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4439 = 3'h3 == state ? _GEN_3668 : ram_0_72; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4440 = 3'h3 == state ? _GEN_3669 : ram_0_73; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4441 = 3'h3 == state ? _GEN_3670 : ram_0_74; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4442 = 3'h3 == state ? _GEN_3671 : ram_0_75; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4443 = 3'h3 == state ? _GEN_3672 : ram_0_76; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4444 = 3'h3 == state ? _GEN_3673 : ram_0_77; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4445 = 3'h3 == state ? _GEN_3674 : ram_0_78; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4446 = 3'h3 == state ? _GEN_3675 : ram_0_79; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4447 = 3'h3 == state ? _GEN_3676 : ram_0_80; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4448 = 3'h3 == state ? _GEN_3677 : ram_0_81; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4449 = 3'h3 == state ? _GEN_3678 : ram_0_82; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4450 = 3'h3 == state ? _GEN_3679 : ram_0_83; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4451 = 3'h3 == state ? _GEN_3680 : ram_0_84; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4452 = 3'h3 == state ? _GEN_3681 : ram_0_85; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4453 = 3'h3 == state ? _GEN_3682 : ram_0_86; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4454 = 3'h3 == state ? _GEN_3683 : ram_0_87; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4455 = 3'h3 == state ? _GEN_3684 : ram_0_88; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4456 = 3'h3 == state ? _GEN_3685 : ram_0_89; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4457 = 3'h3 == state ? _GEN_3686 : ram_0_90; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4458 = 3'h3 == state ? _GEN_3687 : ram_0_91; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4459 = 3'h3 == state ? _GEN_3688 : ram_0_92; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4460 = 3'h3 == state ? _GEN_3689 : ram_0_93; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4461 = 3'h3 == state ? _GEN_3690 : ram_0_94; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4462 = 3'h3 == state ? _GEN_3691 : ram_0_95; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4463 = 3'h3 == state ? _GEN_3692 : ram_0_96; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4464 = 3'h3 == state ? _GEN_3693 : ram_0_97; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4465 = 3'h3 == state ? _GEN_3694 : ram_0_98; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4466 = 3'h3 == state ? _GEN_3695 : ram_0_99; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4467 = 3'h3 == state ? _GEN_3696 : ram_0_100; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4468 = 3'h3 == state ? _GEN_3697 : ram_0_101; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4469 = 3'h3 == state ? _GEN_3698 : ram_0_102; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4470 = 3'h3 == state ? _GEN_3699 : ram_0_103; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4471 = 3'h3 == state ? _GEN_3700 : ram_0_104; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4472 = 3'h3 == state ? _GEN_3701 : ram_0_105; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4473 = 3'h3 == state ? _GEN_3702 : ram_0_106; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4474 = 3'h3 == state ? _GEN_3703 : ram_0_107; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4475 = 3'h3 == state ? _GEN_3704 : ram_0_108; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4476 = 3'h3 == state ? _GEN_3705 : ram_0_109; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4477 = 3'h3 == state ? _GEN_3706 : ram_0_110; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4478 = 3'h3 == state ? _GEN_3707 : ram_0_111; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4479 = 3'h3 == state ? _GEN_3708 : ram_0_112; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4480 = 3'h3 == state ? _GEN_3709 : ram_0_113; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4481 = 3'h3 == state ? _GEN_3710 : ram_0_114; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4482 = 3'h3 == state ? _GEN_3711 : ram_0_115; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4483 = 3'h3 == state ? _GEN_3712 : ram_0_116; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4484 = 3'h3 == state ? _GEN_3713 : ram_0_117; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4485 = 3'h3 == state ? _GEN_3714 : ram_0_118; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4486 = 3'h3 == state ? _GEN_3715 : ram_0_119; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4487 = 3'h3 == state ? _GEN_3716 : ram_0_120; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4488 = 3'h3 == state ? _GEN_3717 : ram_0_121; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4489 = 3'h3 == state ? _GEN_3718 : ram_0_122; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4490 = 3'h3 == state ? _GEN_3719 : ram_0_123; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4491 = 3'h3 == state ? _GEN_3720 : ram_0_124; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4492 = 3'h3 == state ? _GEN_3721 : ram_0_125; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4493 = 3'h3 == state ? _GEN_3722 : ram_0_126; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4494 = 3'h3 == state ? _GEN_3723 : ram_0_127; // @[i_cache.scala 55:18 17:24]
  wire [31:0] _GEN_4495 = 3'h3 == state ? _GEN_3724 : tag_0_0; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4496 = 3'h3 == state ? _GEN_3725 : tag_0_1; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4497 = 3'h3 == state ? _GEN_3726 : tag_0_2; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4498 = 3'h3 == state ? _GEN_3727 : tag_0_3; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4499 = 3'h3 == state ? _GEN_3728 : tag_0_4; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4500 = 3'h3 == state ? _GEN_3729 : tag_0_5; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4501 = 3'h3 == state ? _GEN_3730 : tag_0_6; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4502 = 3'h3 == state ? _GEN_3731 : tag_0_7; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4503 = 3'h3 == state ? _GEN_3732 : tag_0_8; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4504 = 3'h3 == state ? _GEN_3733 : tag_0_9; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4505 = 3'h3 == state ? _GEN_3734 : tag_0_10; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4506 = 3'h3 == state ? _GEN_3735 : tag_0_11; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4507 = 3'h3 == state ? _GEN_3736 : tag_0_12; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4508 = 3'h3 == state ? _GEN_3737 : tag_0_13; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4509 = 3'h3 == state ? _GEN_3738 : tag_0_14; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4510 = 3'h3 == state ? _GEN_3739 : tag_0_15; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4511 = 3'h3 == state ? _GEN_3740 : tag_0_16; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4512 = 3'h3 == state ? _GEN_3741 : tag_0_17; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4513 = 3'h3 == state ? _GEN_3742 : tag_0_18; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4514 = 3'h3 == state ? _GEN_3743 : tag_0_19; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4515 = 3'h3 == state ? _GEN_3744 : tag_0_20; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4516 = 3'h3 == state ? _GEN_3745 : tag_0_21; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4517 = 3'h3 == state ? _GEN_3746 : tag_0_22; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4518 = 3'h3 == state ? _GEN_3747 : tag_0_23; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4519 = 3'h3 == state ? _GEN_3748 : tag_0_24; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4520 = 3'h3 == state ? _GEN_3749 : tag_0_25; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4521 = 3'h3 == state ? _GEN_3750 : tag_0_26; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4522 = 3'h3 == state ? _GEN_3751 : tag_0_27; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4523 = 3'h3 == state ? _GEN_3752 : tag_0_28; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4524 = 3'h3 == state ? _GEN_3753 : tag_0_29; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4525 = 3'h3 == state ? _GEN_3754 : tag_0_30; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4526 = 3'h3 == state ? _GEN_3755 : tag_0_31; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4527 = 3'h3 == state ? _GEN_3756 : tag_0_32; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4528 = 3'h3 == state ? _GEN_3757 : tag_0_33; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4529 = 3'h3 == state ? _GEN_3758 : tag_0_34; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4530 = 3'h3 == state ? _GEN_3759 : tag_0_35; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4531 = 3'h3 == state ? _GEN_3760 : tag_0_36; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4532 = 3'h3 == state ? _GEN_3761 : tag_0_37; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4533 = 3'h3 == state ? _GEN_3762 : tag_0_38; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4534 = 3'h3 == state ? _GEN_3763 : tag_0_39; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4535 = 3'h3 == state ? _GEN_3764 : tag_0_40; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4536 = 3'h3 == state ? _GEN_3765 : tag_0_41; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4537 = 3'h3 == state ? _GEN_3766 : tag_0_42; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4538 = 3'h3 == state ? _GEN_3767 : tag_0_43; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4539 = 3'h3 == state ? _GEN_3768 : tag_0_44; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4540 = 3'h3 == state ? _GEN_3769 : tag_0_45; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4541 = 3'h3 == state ? _GEN_3770 : tag_0_46; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4542 = 3'h3 == state ? _GEN_3771 : tag_0_47; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4543 = 3'h3 == state ? _GEN_3772 : tag_0_48; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4544 = 3'h3 == state ? _GEN_3773 : tag_0_49; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4545 = 3'h3 == state ? _GEN_3774 : tag_0_50; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4546 = 3'h3 == state ? _GEN_3775 : tag_0_51; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4547 = 3'h3 == state ? _GEN_3776 : tag_0_52; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4548 = 3'h3 == state ? _GEN_3777 : tag_0_53; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4549 = 3'h3 == state ? _GEN_3778 : tag_0_54; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4550 = 3'h3 == state ? _GEN_3779 : tag_0_55; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4551 = 3'h3 == state ? _GEN_3780 : tag_0_56; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4552 = 3'h3 == state ? _GEN_3781 : tag_0_57; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4553 = 3'h3 == state ? _GEN_3782 : tag_0_58; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4554 = 3'h3 == state ? _GEN_3783 : tag_0_59; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4555 = 3'h3 == state ? _GEN_3784 : tag_0_60; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4556 = 3'h3 == state ? _GEN_3785 : tag_0_61; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4557 = 3'h3 == state ? _GEN_3786 : tag_0_62; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4558 = 3'h3 == state ? _GEN_3787 : tag_0_63; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4559 = 3'h3 == state ? _GEN_3788 : tag_0_64; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4560 = 3'h3 == state ? _GEN_3789 : tag_0_65; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4561 = 3'h3 == state ? _GEN_3790 : tag_0_66; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4562 = 3'h3 == state ? _GEN_3791 : tag_0_67; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4563 = 3'h3 == state ? _GEN_3792 : tag_0_68; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4564 = 3'h3 == state ? _GEN_3793 : tag_0_69; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4565 = 3'h3 == state ? _GEN_3794 : tag_0_70; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4566 = 3'h3 == state ? _GEN_3795 : tag_0_71; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4567 = 3'h3 == state ? _GEN_3796 : tag_0_72; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4568 = 3'h3 == state ? _GEN_3797 : tag_0_73; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4569 = 3'h3 == state ? _GEN_3798 : tag_0_74; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4570 = 3'h3 == state ? _GEN_3799 : tag_0_75; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4571 = 3'h3 == state ? _GEN_3800 : tag_0_76; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4572 = 3'h3 == state ? _GEN_3801 : tag_0_77; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4573 = 3'h3 == state ? _GEN_3802 : tag_0_78; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4574 = 3'h3 == state ? _GEN_3803 : tag_0_79; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4575 = 3'h3 == state ? _GEN_3804 : tag_0_80; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4576 = 3'h3 == state ? _GEN_3805 : tag_0_81; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4577 = 3'h3 == state ? _GEN_3806 : tag_0_82; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4578 = 3'h3 == state ? _GEN_3807 : tag_0_83; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4579 = 3'h3 == state ? _GEN_3808 : tag_0_84; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4580 = 3'h3 == state ? _GEN_3809 : tag_0_85; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4581 = 3'h3 == state ? _GEN_3810 : tag_0_86; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4582 = 3'h3 == state ? _GEN_3811 : tag_0_87; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4583 = 3'h3 == state ? _GEN_3812 : tag_0_88; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4584 = 3'h3 == state ? _GEN_3813 : tag_0_89; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4585 = 3'h3 == state ? _GEN_3814 : tag_0_90; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4586 = 3'h3 == state ? _GEN_3815 : tag_0_91; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4587 = 3'h3 == state ? _GEN_3816 : tag_0_92; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4588 = 3'h3 == state ? _GEN_3817 : tag_0_93; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4589 = 3'h3 == state ? _GEN_3818 : tag_0_94; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4590 = 3'h3 == state ? _GEN_3819 : tag_0_95; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4591 = 3'h3 == state ? _GEN_3820 : tag_0_96; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4592 = 3'h3 == state ? _GEN_3821 : tag_0_97; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4593 = 3'h3 == state ? _GEN_3822 : tag_0_98; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4594 = 3'h3 == state ? _GEN_3823 : tag_0_99; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4595 = 3'h3 == state ? _GEN_3824 : tag_0_100; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4596 = 3'h3 == state ? _GEN_3825 : tag_0_101; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4597 = 3'h3 == state ? _GEN_3826 : tag_0_102; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4598 = 3'h3 == state ? _GEN_3827 : tag_0_103; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4599 = 3'h3 == state ? _GEN_3828 : tag_0_104; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4600 = 3'h3 == state ? _GEN_3829 : tag_0_105; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4601 = 3'h3 == state ? _GEN_3830 : tag_0_106; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4602 = 3'h3 == state ? _GEN_3831 : tag_0_107; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4603 = 3'h3 == state ? _GEN_3832 : tag_0_108; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4604 = 3'h3 == state ? _GEN_3833 : tag_0_109; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4605 = 3'h3 == state ? _GEN_3834 : tag_0_110; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4606 = 3'h3 == state ? _GEN_3835 : tag_0_111; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4607 = 3'h3 == state ? _GEN_3836 : tag_0_112; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4608 = 3'h3 == state ? _GEN_3837 : tag_0_113; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4609 = 3'h3 == state ? _GEN_3838 : tag_0_114; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4610 = 3'h3 == state ? _GEN_3839 : tag_0_115; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4611 = 3'h3 == state ? _GEN_3840 : tag_0_116; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4612 = 3'h3 == state ? _GEN_3841 : tag_0_117; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4613 = 3'h3 == state ? _GEN_3842 : tag_0_118; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4614 = 3'h3 == state ? _GEN_3843 : tag_0_119; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4615 = 3'h3 == state ? _GEN_3844 : tag_0_120; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4616 = 3'h3 == state ? _GEN_3845 : tag_0_121; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4617 = 3'h3 == state ? _GEN_3846 : tag_0_122; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4618 = 3'h3 == state ? _GEN_3847 : tag_0_123; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4619 = 3'h3 == state ? _GEN_3848 : tag_0_124; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4620 = 3'h3 == state ? _GEN_3849 : tag_0_125; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4621 = 3'h3 == state ? _GEN_3850 : tag_0_126; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4622 = 3'h3 == state ? _GEN_3851 : tag_0_127; // @[i_cache.scala 55:18 19:24]
  wire  _GEN_4623 = 3'h3 == state ? _GEN_3852 : valid_0_0; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4624 = 3'h3 == state ? _GEN_3853 : valid_0_1; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4625 = 3'h3 == state ? _GEN_3854 : valid_0_2; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4626 = 3'h3 == state ? _GEN_3855 : valid_0_3; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4627 = 3'h3 == state ? _GEN_3856 : valid_0_4; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4628 = 3'h3 == state ? _GEN_3857 : valid_0_5; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4629 = 3'h3 == state ? _GEN_3858 : valid_0_6; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4630 = 3'h3 == state ? _GEN_3859 : valid_0_7; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4631 = 3'h3 == state ? _GEN_3860 : valid_0_8; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4632 = 3'h3 == state ? _GEN_3861 : valid_0_9; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4633 = 3'h3 == state ? _GEN_3862 : valid_0_10; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4634 = 3'h3 == state ? _GEN_3863 : valid_0_11; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4635 = 3'h3 == state ? _GEN_3864 : valid_0_12; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4636 = 3'h3 == state ? _GEN_3865 : valid_0_13; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4637 = 3'h3 == state ? _GEN_3866 : valid_0_14; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4638 = 3'h3 == state ? _GEN_3867 : valid_0_15; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4639 = 3'h3 == state ? _GEN_3868 : valid_0_16; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4640 = 3'h3 == state ? _GEN_3869 : valid_0_17; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4641 = 3'h3 == state ? _GEN_3870 : valid_0_18; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4642 = 3'h3 == state ? _GEN_3871 : valid_0_19; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4643 = 3'h3 == state ? _GEN_3872 : valid_0_20; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4644 = 3'h3 == state ? _GEN_3873 : valid_0_21; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4645 = 3'h3 == state ? _GEN_3874 : valid_0_22; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4646 = 3'h3 == state ? _GEN_3875 : valid_0_23; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4647 = 3'h3 == state ? _GEN_3876 : valid_0_24; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4648 = 3'h3 == state ? _GEN_3877 : valid_0_25; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4649 = 3'h3 == state ? _GEN_3878 : valid_0_26; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4650 = 3'h3 == state ? _GEN_3879 : valid_0_27; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4651 = 3'h3 == state ? _GEN_3880 : valid_0_28; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4652 = 3'h3 == state ? _GEN_3881 : valid_0_29; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4653 = 3'h3 == state ? _GEN_3882 : valid_0_30; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4654 = 3'h3 == state ? _GEN_3883 : valid_0_31; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4655 = 3'h3 == state ? _GEN_3884 : valid_0_32; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4656 = 3'h3 == state ? _GEN_3885 : valid_0_33; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4657 = 3'h3 == state ? _GEN_3886 : valid_0_34; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4658 = 3'h3 == state ? _GEN_3887 : valid_0_35; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4659 = 3'h3 == state ? _GEN_3888 : valid_0_36; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4660 = 3'h3 == state ? _GEN_3889 : valid_0_37; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4661 = 3'h3 == state ? _GEN_3890 : valid_0_38; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4662 = 3'h3 == state ? _GEN_3891 : valid_0_39; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4663 = 3'h3 == state ? _GEN_3892 : valid_0_40; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4664 = 3'h3 == state ? _GEN_3893 : valid_0_41; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4665 = 3'h3 == state ? _GEN_3894 : valid_0_42; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4666 = 3'h3 == state ? _GEN_3895 : valid_0_43; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4667 = 3'h3 == state ? _GEN_3896 : valid_0_44; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4668 = 3'h3 == state ? _GEN_3897 : valid_0_45; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4669 = 3'h3 == state ? _GEN_3898 : valid_0_46; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4670 = 3'h3 == state ? _GEN_3899 : valid_0_47; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4671 = 3'h3 == state ? _GEN_3900 : valid_0_48; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4672 = 3'h3 == state ? _GEN_3901 : valid_0_49; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4673 = 3'h3 == state ? _GEN_3902 : valid_0_50; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4674 = 3'h3 == state ? _GEN_3903 : valid_0_51; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4675 = 3'h3 == state ? _GEN_3904 : valid_0_52; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4676 = 3'h3 == state ? _GEN_3905 : valid_0_53; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4677 = 3'h3 == state ? _GEN_3906 : valid_0_54; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4678 = 3'h3 == state ? _GEN_3907 : valid_0_55; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4679 = 3'h3 == state ? _GEN_3908 : valid_0_56; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4680 = 3'h3 == state ? _GEN_3909 : valid_0_57; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4681 = 3'h3 == state ? _GEN_3910 : valid_0_58; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4682 = 3'h3 == state ? _GEN_3911 : valid_0_59; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4683 = 3'h3 == state ? _GEN_3912 : valid_0_60; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4684 = 3'h3 == state ? _GEN_3913 : valid_0_61; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4685 = 3'h3 == state ? _GEN_3914 : valid_0_62; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4686 = 3'h3 == state ? _GEN_3915 : valid_0_63; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4687 = 3'h3 == state ? _GEN_3916 : valid_0_64; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4688 = 3'h3 == state ? _GEN_3917 : valid_0_65; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4689 = 3'h3 == state ? _GEN_3918 : valid_0_66; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4690 = 3'h3 == state ? _GEN_3919 : valid_0_67; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4691 = 3'h3 == state ? _GEN_3920 : valid_0_68; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4692 = 3'h3 == state ? _GEN_3921 : valid_0_69; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4693 = 3'h3 == state ? _GEN_3922 : valid_0_70; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4694 = 3'h3 == state ? _GEN_3923 : valid_0_71; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4695 = 3'h3 == state ? _GEN_3924 : valid_0_72; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4696 = 3'h3 == state ? _GEN_3925 : valid_0_73; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4697 = 3'h3 == state ? _GEN_3926 : valid_0_74; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4698 = 3'h3 == state ? _GEN_3927 : valid_0_75; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4699 = 3'h3 == state ? _GEN_3928 : valid_0_76; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4700 = 3'h3 == state ? _GEN_3929 : valid_0_77; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4701 = 3'h3 == state ? _GEN_3930 : valid_0_78; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4702 = 3'h3 == state ? _GEN_3931 : valid_0_79; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4703 = 3'h3 == state ? _GEN_3932 : valid_0_80; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4704 = 3'h3 == state ? _GEN_3933 : valid_0_81; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4705 = 3'h3 == state ? _GEN_3934 : valid_0_82; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4706 = 3'h3 == state ? _GEN_3935 : valid_0_83; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4707 = 3'h3 == state ? _GEN_3936 : valid_0_84; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4708 = 3'h3 == state ? _GEN_3937 : valid_0_85; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4709 = 3'h3 == state ? _GEN_3938 : valid_0_86; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4710 = 3'h3 == state ? _GEN_3939 : valid_0_87; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4711 = 3'h3 == state ? _GEN_3940 : valid_0_88; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4712 = 3'h3 == state ? _GEN_3941 : valid_0_89; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4713 = 3'h3 == state ? _GEN_3942 : valid_0_90; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4714 = 3'h3 == state ? _GEN_3943 : valid_0_91; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4715 = 3'h3 == state ? _GEN_3944 : valid_0_92; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4716 = 3'h3 == state ? _GEN_3945 : valid_0_93; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4717 = 3'h3 == state ? _GEN_3946 : valid_0_94; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4718 = 3'h3 == state ? _GEN_3947 : valid_0_95; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4719 = 3'h3 == state ? _GEN_3948 : valid_0_96; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4720 = 3'h3 == state ? _GEN_3949 : valid_0_97; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4721 = 3'h3 == state ? _GEN_3950 : valid_0_98; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4722 = 3'h3 == state ? _GEN_3951 : valid_0_99; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4723 = 3'h3 == state ? _GEN_3952 : valid_0_100; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4724 = 3'h3 == state ? _GEN_3953 : valid_0_101; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4725 = 3'h3 == state ? _GEN_3954 : valid_0_102; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4726 = 3'h3 == state ? _GEN_3955 : valid_0_103; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4727 = 3'h3 == state ? _GEN_3956 : valid_0_104; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4728 = 3'h3 == state ? _GEN_3957 : valid_0_105; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4729 = 3'h3 == state ? _GEN_3958 : valid_0_106; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4730 = 3'h3 == state ? _GEN_3959 : valid_0_107; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4731 = 3'h3 == state ? _GEN_3960 : valid_0_108; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4732 = 3'h3 == state ? _GEN_3961 : valid_0_109; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4733 = 3'h3 == state ? _GEN_3962 : valid_0_110; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4734 = 3'h3 == state ? _GEN_3963 : valid_0_111; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4735 = 3'h3 == state ? _GEN_3964 : valid_0_112; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4736 = 3'h3 == state ? _GEN_3965 : valid_0_113; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4737 = 3'h3 == state ? _GEN_3966 : valid_0_114; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4738 = 3'h3 == state ? _GEN_3967 : valid_0_115; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4739 = 3'h3 == state ? _GEN_3968 : valid_0_116; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4740 = 3'h3 == state ? _GEN_3969 : valid_0_117; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4741 = 3'h3 == state ? _GEN_3970 : valid_0_118; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4742 = 3'h3 == state ? _GEN_3971 : valid_0_119; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4743 = 3'h3 == state ? _GEN_3972 : valid_0_120; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4744 = 3'h3 == state ? _GEN_3973 : valid_0_121; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4745 = 3'h3 == state ? _GEN_3974 : valid_0_122; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4746 = 3'h3 == state ? _GEN_3975 : valid_0_123; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4747 = 3'h3 == state ? _GEN_3976 : valid_0_124; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4748 = 3'h3 == state ? _GEN_3977 : valid_0_125; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4749 = 3'h3 == state ? _GEN_3978 : valid_0_126; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4750 = 3'h3 == state ? _GEN_3979 : valid_0_127; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4751 = 3'h3 == state ? _GEN_3980 : quene; // @[i_cache.scala 55:18 28:24]
  wire [63:0] _GEN_4752 = 3'h3 == state ? _GEN_3981 : ram_1_0; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4753 = 3'h3 == state ? _GEN_3982 : ram_1_1; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4754 = 3'h3 == state ? _GEN_3983 : ram_1_2; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4755 = 3'h3 == state ? _GEN_3984 : ram_1_3; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4756 = 3'h3 == state ? _GEN_3985 : ram_1_4; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4757 = 3'h3 == state ? _GEN_3986 : ram_1_5; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4758 = 3'h3 == state ? _GEN_3987 : ram_1_6; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4759 = 3'h3 == state ? _GEN_3988 : ram_1_7; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4760 = 3'h3 == state ? _GEN_3989 : ram_1_8; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4761 = 3'h3 == state ? _GEN_3990 : ram_1_9; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4762 = 3'h3 == state ? _GEN_3991 : ram_1_10; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4763 = 3'h3 == state ? _GEN_3992 : ram_1_11; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4764 = 3'h3 == state ? _GEN_3993 : ram_1_12; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4765 = 3'h3 == state ? _GEN_3994 : ram_1_13; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4766 = 3'h3 == state ? _GEN_3995 : ram_1_14; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4767 = 3'h3 == state ? _GEN_3996 : ram_1_15; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4768 = 3'h3 == state ? _GEN_3997 : ram_1_16; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4769 = 3'h3 == state ? _GEN_3998 : ram_1_17; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4770 = 3'h3 == state ? _GEN_3999 : ram_1_18; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4771 = 3'h3 == state ? _GEN_4000 : ram_1_19; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4772 = 3'h3 == state ? _GEN_4001 : ram_1_20; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4773 = 3'h3 == state ? _GEN_4002 : ram_1_21; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4774 = 3'h3 == state ? _GEN_4003 : ram_1_22; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4775 = 3'h3 == state ? _GEN_4004 : ram_1_23; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4776 = 3'h3 == state ? _GEN_4005 : ram_1_24; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4777 = 3'h3 == state ? _GEN_4006 : ram_1_25; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4778 = 3'h3 == state ? _GEN_4007 : ram_1_26; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4779 = 3'h3 == state ? _GEN_4008 : ram_1_27; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4780 = 3'h3 == state ? _GEN_4009 : ram_1_28; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4781 = 3'h3 == state ? _GEN_4010 : ram_1_29; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4782 = 3'h3 == state ? _GEN_4011 : ram_1_30; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4783 = 3'h3 == state ? _GEN_4012 : ram_1_31; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4784 = 3'h3 == state ? _GEN_4013 : ram_1_32; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4785 = 3'h3 == state ? _GEN_4014 : ram_1_33; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4786 = 3'h3 == state ? _GEN_4015 : ram_1_34; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4787 = 3'h3 == state ? _GEN_4016 : ram_1_35; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4788 = 3'h3 == state ? _GEN_4017 : ram_1_36; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4789 = 3'h3 == state ? _GEN_4018 : ram_1_37; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4790 = 3'h3 == state ? _GEN_4019 : ram_1_38; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4791 = 3'h3 == state ? _GEN_4020 : ram_1_39; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4792 = 3'h3 == state ? _GEN_4021 : ram_1_40; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4793 = 3'h3 == state ? _GEN_4022 : ram_1_41; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4794 = 3'h3 == state ? _GEN_4023 : ram_1_42; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4795 = 3'h3 == state ? _GEN_4024 : ram_1_43; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4796 = 3'h3 == state ? _GEN_4025 : ram_1_44; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4797 = 3'h3 == state ? _GEN_4026 : ram_1_45; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4798 = 3'h3 == state ? _GEN_4027 : ram_1_46; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4799 = 3'h3 == state ? _GEN_4028 : ram_1_47; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4800 = 3'h3 == state ? _GEN_4029 : ram_1_48; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4801 = 3'h3 == state ? _GEN_4030 : ram_1_49; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4802 = 3'h3 == state ? _GEN_4031 : ram_1_50; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4803 = 3'h3 == state ? _GEN_4032 : ram_1_51; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4804 = 3'h3 == state ? _GEN_4033 : ram_1_52; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4805 = 3'h3 == state ? _GEN_4034 : ram_1_53; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4806 = 3'h3 == state ? _GEN_4035 : ram_1_54; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4807 = 3'h3 == state ? _GEN_4036 : ram_1_55; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4808 = 3'h3 == state ? _GEN_4037 : ram_1_56; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4809 = 3'h3 == state ? _GEN_4038 : ram_1_57; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4810 = 3'h3 == state ? _GEN_4039 : ram_1_58; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4811 = 3'h3 == state ? _GEN_4040 : ram_1_59; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4812 = 3'h3 == state ? _GEN_4041 : ram_1_60; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4813 = 3'h3 == state ? _GEN_4042 : ram_1_61; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4814 = 3'h3 == state ? _GEN_4043 : ram_1_62; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4815 = 3'h3 == state ? _GEN_4044 : ram_1_63; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4816 = 3'h3 == state ? _GEN_4045 : ram_1_64; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4817 = 3'h3 == state ? _GEN_4046 : ram_1_65; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4818 = 3'h3 == state ? _GEN_4047 : ram_1_66; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4819 = 3'h3 == state ? _GEN_4048 : ram_1_67; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4820 = 3'h3 == state ? _GEN_4049 : ram_1_68; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4821 = 3'h3 == state ? _GEN_4050 : ram_1_69; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4822 = 3'h3 == state ? _GEN_4051 : ram_1_70; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4823 = 3'h3 == state ? _GEN_4052 : ram_1_71; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4824 = 3'h3 == state ? _GEN_4053 : ram_1_72; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4825 = 3'h3 == state ? _GEN_4054 : ram_1_73; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4826 = 3'h3 == state ? _GEN_4055 : ram_1_74; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4827 = 3'h3 == state ? _GEN_4056 : ram_1_75; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4828 = 3'h3 == state ? _GEN_4057 : ram_1_76; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4829 = 3'h3 == state ? _GEN_4058 : ram_1_77; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4830 = 3'h3 == state ? _GEN_4059 : ram_1_78; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4831 = 3'h3 == state ? _GEN_4060 : ram_1_79; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4832 = 3'h3 == state ? _GEN_4061 : ram_1_80; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4833 = 3'h3 == state ? _GEN_4062 : ram_1_81; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4834 = 3'h3 == state ? _GEN_4063 : ram_1_82; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4835 = 3'h3 == state ? _GEN_4064 : ram_1_83; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4836 = 3'h3 == state ? _GEN_4065 : ram_1_84; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4837 = 3'h3 == state ? _GEN_4066 : ram_1_85; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4838 = 3'h3 == state ? _GEN_4067 : ram_1_86; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4839 = 3'h3 == state ? _GEN_4068 : ram_1_87; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4840 = 3'h3 == state ? _GEN_4069 : ram_1_88; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4841 = 3'h3 == state ? _GEN_4070 : ram_1_89; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4842 = 3'h3 == state ? _GEN_4071 : ram_1_90; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4843 = 3'h3 == state ? _GEN_4072 : ram_1_91; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4844 = 3'h3 == state ? _GEN_4073 : ram_1_92; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4845 = 3'h3 == state ? _GEN_4074 : ram_1_93; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4846 = 3'h3 == state ? _GEN_4075 : ram_1_94; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4847 = 3'h3 == state ? _GEN_4076 : ram_1_95; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4848 = 3'h3 == state ? _GEN_4077 : ram_1_96; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4849 = 3'h3 == state ? _GEN_4078 : ram_1_97; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4850 = 3'h3 == state ? _GEN_4079 : ram_1_98; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4851 = 3'h3 == state ? _GEN_4080 : ram_1_99; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4852 = 3'h3 == state ? _GEN_4081 : ram_1_100; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4853 = 3'h3 == state ? _GEN_4082 : ram_1_101; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4854 = 3'h3 == state ? _GEN_4083 : ram_1_102; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4855 = 3'h3 == state ? _GEN_4084 : ram_1_103; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4856 = 3'h3 == state ? _GEN_4085 : ram_1_104; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4857 = 3'h3 == state ? _GEN_4086 : ram_1_105; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4858 = 3'h3 == state ? _GEN_4087 : ram_1_106; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4859 = 3'h3 == state ? _GEN_4088 : ram_1_107; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4860 = 3'h3 == state ? _GEN_4089 : ram_1_108; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4861 = 3'h3 == state ? _GEN_4090 : ram_1_109; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4862 = 3'h3 == state ? _GEN_4091 : ram_1_110; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4863 = 3'h3 == state ? _GEN_4092 : ram_1_111; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4864 = 3'h3 == state ? _GEN_4093 : ram_1_112; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4865 = 3'h3 == state ? _GEN_4094 : ram_1_113; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4866 = 3'h3 == state ? _GEN_4095 : ram_1_114; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4867 = 3'h3 == state ? _GEN_4096 : ram_1_115; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4868 = 3'h3 == state ? _GEN_4097 : ram_1_116; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4869 = 3'h3 == state ? _GEN_4098 : ram_1_117; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4870 = 3'h3 == state ? _GEN_4099 : ram_1_118; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4871 = 3'h3 == state ? _GEN_4100 : ram_1_119; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4872 = 3'h3 == state ? _GEN_4101 : ram_1_120; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4873 = 3'h3 == state ? _GEN_4102 : ram_1_121; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4874 = 3'h3 == state ? _GEN_4103 : ram_1_122; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4875 = 3'h3 == state ? _GEN_4104 : ram_1_123; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4876 = 3'h3 == state ? _GEN_4105 : ram_1_124; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4877 = 3'h3 == state ? _GEN_4106 : ram_1_125; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4878 = 3'h3 == state ? _GEN_4107 : ram_1_126; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4879 = 3'h3 == state ? _GEN_4108 : ram_1_127; // @[i_cache.scala 55:18 18:24]
  wire [31:0] _GEN_4880 = 3'h3 == state ? _GEN_4109 : tag_1_0; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4881 = 3'h3 == state ? _GEN_4110 : tag_1_1; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4882 = 3'h3 == state ? _GEN_4111 : tag_1_2; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4883 = 3'h3 == state ? _GEN_4112 : tag_1_3; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4884 = 3'h3 == state ? _GEN_4113 : tag_1_4; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4885 = 3'h3 == state ? _GEN_4114 : tag_1_5; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4886 = 3'h3 == state ? _GEN_4115 : tag_1_6; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4887 = 3'h3 == state ? _GEN_4116 : tag_1_7; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4888 = 3'h3 == state ? _GEN_4117 : tag_1_8; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4889 = 3'h3 == state ? _GEN_4118 : tag_1_9; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4890 = 3'h3 == state ? _GEN_4119 : tag_1_10; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4891 = 3'h3 == state ? _GEN_4120 : tag_1_11; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4892 = 3'h3 == state ? _GEN_4121 : tag_1_12; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4893 = 3'h3 == state ? _GEN_4122 : tag_1_13; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4894 = 3'h3 == state ? _GEN_4123 : tag_1_14; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4895 = 3'h3 == state ? _GEN_4124 : tag_1_15; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4896 = 3'h3 == state ? _GEN_4125 : tag_1_16; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4897 = 3'h3 == state ? _GEN_4126 : tag_1_17; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4898 = 3'h3 == state ? _GEN_4127 : tag_1_18; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4899 = 3'h3 == state ? _GEN_4128 : tag_1_19; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4900 = 3'h3 == state ? _GEN_4129 : tag_1_20; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4901 = 3'h3 == state ? _GEN_4130 : tag_1_21; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4902 = 3'h3 == state ? _GEN_4131 : tag_1_22; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4903 = 3'h3 == state ? _GEN_4132 : tag_1_23; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4904 = 3'h3 == state ? _GEN_4133 : tag_1_24; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4905 = 3'h3 == state ? _GEN_4134 : tag_1_25; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4906 = 3'h3 == state ? _GEN_4135 : tag_1_26; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4907 = 3'h3 == state ? _GEN_4136 : tag_1_27; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4908 = 3'h3 == state ? _GEN_4137 : tag_1_28; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4909 = 3'h3 == state ? _GEN_4138 : tag_1_29; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4910 = 3'h3 == state ? _GEN_4139 : tag_1_30; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4911 = 3'h3 == state ? _GEN_4140 : tag_1_31; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4912 = 3'h3 == state ? _GEN_4141 : tag_1_32; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4913 = 3'h3 == state ? _GEN_4142 : tag_1_33; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4914 = 3'h3 == state ? _GEN_4143 : tag_1_34; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4915 = 3'h3 == state ? _GEN_4144 : tag_1_35; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4916 = 3'h3 == state ? _GEN_4145 : tag_1_36; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4917 = 3'h3 == state ? _GEN_4146 : tag_1_37; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4918 = 3'h3 == state ? _GEN_4147 : tag_1_38; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4919 = 3'h3 == state ? _GEN_4148 : tag_1_39; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4920 = 3'h3 == state ? _GEN_4149 : tag_1_40; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4921 = 3'h3 == state ? _GEN_4150 : tag_1_41; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4922 = 3'h3 == state ? _GEN_4151 : tag_1_42; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4923 = 3'h3 == state ? _GEN_4152 : tag_1_43; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4924 = 3'h3 == state ? _GEN_4153 : tag_1_44; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4925 = 3'h3 == state ? _GEN_4154 : tag_1_45; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4926 = 3'h3 == state ? _GEN_4155 : tag_1_46; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4927 = 3'h3 == state ? _GEN_4156 : tag_1_47; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4928 = 3'h3 == state ? _GEN_4157 : tag_1_48; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4929 = 3'h3 == state ? _GEN_4158 : tag_1_49; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4930 = 3'h3 == state ? _GEN_4159 : tag_1_50; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4931 = 3'h3 == state ? _GEN_4160 : tag_1_51; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4932 = 3'h3 == state ? _GEN_4161 : tag_1_52; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4933 = 3'h3 == state ? _GEN_4162 : tag_1_53; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4934 = 3'h3 == state ? _GEN_4163 : tag_1_54; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4935 = 3'h3 == state ? _GEN_4164 : tag_1_55; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4936 = 3'h3 == state ? _GEN_4165 : tag_1_56; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4937 = 3'h3 == state ? _GEN_4166 : tag_1_57; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4938 = 3'h3 == state ? _GEN_4167 : tag_1_58; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4939 = 3'h3 == state ? _GEN_4168 : tag_1_59; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4940 = 3'h3 == state ? _GEN_4169 : tag_1_60; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4941 = 3'h3 == state ? _GEN_4170 : tag_1_61; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4942 = 3'h3 == state ? _GEN_4171 : tag_1_62; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4943 = 3'h3 == state ? _GEN_4172 : tag_1_63; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4944 = 3'h3 == state ? _GEN_4173 : tag_1_64; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4945 = 3'h3 == state ? _GEN_4174 : tag_1_65; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4946 = 3'h3 == state ? _GEN_4175 : tag_1_66; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4947 = 3'h3 == state ? _GEN_4176 : tag_1_67; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4948 = 3'h3 == state ? _GEN_4177 : tag_1_68; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4949 = 3'h3 == state ? _GEN_4178 : tag_1_69; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4950 = 3'h3 == state ? _GEN_4179 : tag_1_70; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4951 = 3'h3 == state ? _GEN_4180 : tag_1_71; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4952 = 3'h3 == state ? _GEN_4181 : tag_1_72; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4953 = 3'h3 == state ? _GEN_4182 : tag_1_73; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4954 = 3'h3 == state ? _GEN_4183 : tag_1_74; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4955 = 3'h3 == state ? _GEN_4184 : tag_1_75; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4956 = 3'h3 == state ? _GEN_4185 : tag_1_76; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4957 = 3'h3 == state ? _GEN_4186 : tag_1_77; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4958 = 3'h3 == state ? _GEN_4187 : tag_1_78; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4959 = 3'h3 == state ? _GEN_4188 : tag_1_79; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4960 = 3'h3 == state ? _GEN_4189 : tag_1_80; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4961 = 3'h3 == state ? _GEN_4190 : tag_1_81; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4962 = 3'h3 == state ? _GEN_4191 : tag_1_82; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4963 = 3'h3 == state ? _GEN_4192 : tag_1_83; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4964 = 3'h3 == state ? _GEN_4193 : tag_1_84; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4965 = 3'h3 == state ? _GEN_4194 : tag_1_85; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4966 = 3'h3 == state ? _GEN_4195 : tag_1_86; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4967 = 3'h3 == state ? _GEN_4196 : tag_1_87; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4968 = 3'h3 == state ? _GEN_4197 : tag_1_88; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4969 = 3'h3 == state ? _GEN_4198 : tag_1_89; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4970 = 3'h3 == state ? _GEN_4199 : tag_1_90; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4971 = 3'h3 == state ? _GEN_4200 : tag_1_91; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4972 = 3'h3 == state ? _GEN_4201 : tag_1_92; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4973 = 3'h3 == state ? _GEN_4202 : tag_1_93; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4974 = 3'h3 == state ? _GEN_4203 : tag_1_94; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4975 = 3'h3 == state ? _GEN_4204 : tag_1_95; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4976 = 3'h3 == state ? _GEN_4205 : tag_1_96; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4977 = 3'h3 == state ? _GEN_4206 : tag_1_97; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4978 = 3'h3 == state ? _GEN_4207 : tag_1_98; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4979 = 3'h3 == state ? _GEN_4208 : tag_1_99; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4980 = 3'h3 == state ? _GEN_4209 : tag_1_100; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4981 = 3'h3 == state ? _GEN_4210 : tag_1_101; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4982 = 3'h3 == state ? _GEN_4211 : tag_1_102; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4983 = 3'h3 == state ? _GEN_4212 : tag_1_103; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4984 = 3'h3 == state ? _GEN_4213 : tag_1_104; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4985 = 3'h3 == state ? _GEN_4214 : tag_1_105; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4986 = 3'h3 == state ? _GEN_4215 : tag_1_106; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4987 = 3'h3 == state ? _GEN_4216 : tag_1_107; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4988 = 3'h3 == state ? _GEN_4217 : tag_1_108; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4989 = 3'h3 == state ? _GEN_4218 : tag_1_109; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4990 = 3'h3 == state ? _GEN_4219 : tag_1_110; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4991 = 3'h3 == state ? _GEN_4220 : tag_1_111; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4992 = 3'h3 == state ? _GEN_4221 : tag_1_112; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4993 = 3'h3 == state ? _GEN_4222 : tag_1_113; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4994 = 3'h3 == state ? _GEN_4223 : tag_1_114; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4995 = 3'h3 == state ? _GEN_4224 : tag_1_115; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4996 = 3'h3 == state ? _GEN_4225 : tag_1_116; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4997 = 3'h3 == state ? _GEN_4226 : tag_1_117; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4998 = 3'h3 == state ? _GEN_4227 : tag_1_118; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4999 = 3'h3 == state ? _GEN_4228 : tag_1_119; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5000 = 3'h3 == state ? _GEN_4229 : tag_1_120; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5001 = 3'h3 == state ? _GEN_4230 : tag_1_121; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5002 = 3'h3 == state ? _GEN_4231 : tag_1_122; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5003 = 3'h3 == state ? _GEN_4232 : tag_1_123; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5004 = 3'h3 == state ? _GEN_4233 : tag_1_124; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5005 = 3'h3 == state ? _GEN_4234 : tag_1_125; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5006 = 3'h3 == state ? _GEN_4235 : tag_1_126; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5007 = 3'h3 == state ? _GEN_4236 : tag_1_127; // @[i_cache.scala 55:18 20:24]
  wire  _GEN_5008 = 3'h3 == state ? _GEN_4237 : valid_1_0; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5009 = 3'h3 == state ? _GEN_4238 : valid_1_1; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5010 = 3'h3 == state ? _GEN_4239 : valid_1_2; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5011 = 3'h3 == state ? _GEN_4240 : valid_1_3; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5012 = 3'h3 == state ? _GEN_4241 : valid_1_4; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5013 = 3'h3 == state ? _GEN_4242 : valid_1_5; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5014 = 3'h3 == state ? _GEN_4243 : valid_1_6; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5015 = 3'h3 == state ? _GEN_4244 : valid_1_7; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5016 = 3'h3 == state ? _GEN_4245 : valid_1_8; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5017 = 3'h3 == state ? _GEN_4246 : valid_1_9; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5018 = 3'h3 == state ? _GEN_4247 : valid_1_10; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5019 = 3'h3 == state ? _GEN_4248 : valid_1_11; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5020 = 3'h3 == state ? _GEN_4249 : valid_1_12; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5021 = 3'h3 == state ? _GEN_4250 : valid_1_13; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5022 = 3'h3 == state ? _GEN_4251 : valid_1_14; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5023 = 3'h3 == state ? _GEN_4252 : valid_1_15; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5024 = 3'h3 == state ? _GEN_4253 : valid_1_16; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5025 = 3'h3 == state ? _GEN_4254 : valid_1_17; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5026 = 3'h3 == state ? _GEN_4255 : valid_1_18; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5027 = 3'h3 == state ? _GEN_4256 : valid_1_19; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5028 = 3'h3 == state ? _GEN_4257 : valid_1_20; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5029 = 3'h3 == state ? _GEN_4258 : valid_1_21; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5030 = 3'h3 == state ? _GEN_4259 : valid_1_22; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5031 = 3'h3 == state ? _GEN_4260 : valid_1_23; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5032 = 3'h3 == state ? _GEN_4261 : valid_1_24; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5033 = 3'h3 == state ? _GEN_4262 : valid_1_25; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5034 = 3'h3 == state ? _GEN_4263 : valid_1_26; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5035 = 3'h3 == state ? _GEN_4264 : valid_1_27; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5036 = 3'h3 == state ? _GEN_4265 : valid_1_28; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5037 = 3'h3 == state ? _GEN_4266 : valid_1_29; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5038 = 3'h3 == state ? _GEN_4267 : valid_1_30; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5039 = 3'h3 == state ? _GEN_4268 : valid_1_31; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5040 = 3'h3 == state ? _GEN_4269 : valid_1_32; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5041 = 3'h3 == state ? _GEN_4270 : valid_1_33; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5042 = 3'h3 == state ? _GEN_4271 : valid_1_34; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5043 = 3'h3 == state ? _GEN_4272 : valid_1_35; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5044 = 3'h3 == state ? _GEN_4273 : valid_1_36; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5045 = 3'h3 == state ? _GEN_4274 : valid_1_37; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5046 = 3'h3 == state ? _GEN_4275 : valid_1_38; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5047 = 3'h3 == state ? _GEN_4276 : valid_1_39; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5048 = 3'h3 == state ? _GEN_4277 : valid_1_40; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5049 = 3'h3 == state ? _GEN_4278 : valid_1_41; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5050 = 3'h3 == state ? _GEN_4279 : valid_1_42; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5051 = 3'h3 == state ? _GEN_4280 : valid_1_43; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5052 = 3'h3 == state ? _GEN_4281 : valid_1_44; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5053 = 3'h3 == state ? _GEN_4282 : valid_1_45; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5054 = 3'h3 == state ? _GEN_4283 : valid_1_46; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5055 = 3'h3 == state ? _GEN_4284 : valid_1_47; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5056 = 3'h3 == state ? _GEN_4285 : valid_1_48; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5057 = 3'h3 == state ? _GEN_4286 : valid_1_49; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5058 = 3'h3 == state ? _GEN_4287 : valid_1_50; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5059 = 3'h3 == state ? _GEN_4288 : valid_1_51; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5060 = 3'h3 == state ? _GEN_4289 : valid_1_52; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5061 = 3'h3 == state ? _GEN_4290 : valid_1_53; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5062 = 3'h3 == state ? _GEN_4291 : valid_1_54; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5063 = 3'h3 == state ? _GEN_4292 : valid_1_55; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5064 = 3'h3 == state ? _GEN_4293 : valid_1_56; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5065 = 3'h3 == state ? _GEN_4294 : valid_1_57; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5066 = 3'h3 == state ? _GEN_4295 : valid_1_58; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5067 = 3'h3 == state ? _GEN_4296 : valid_1_59; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5068 = 3'h3 == state ? _GEN_4297 : valid_1_60; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5069 = 3'h3 == state ? _GEN_4298 : valid_1_61; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5070 = 3'h3 == state ? _GEN_4299 : valid_1_62; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5071 = 3'h3 == state ? _GEN_4300 : valid_1_63; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5072 = 3'h3 == state ? _GEN_4301 : valid_1_64; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5073 = 3'h3 == state ? _GEN_4302 : valid_1_65; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5074 = 3'h3 == state ? _GEN_4303 : valid_1_66; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5075 = 3'h3 == state ? _GEN_4304 : valid_1_67; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5076 = 3'h3 == state ? _GEN_4305 : valid_1_68; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5077 = 3'h3 == state ? _GEN_4306 : valid_1_69; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5078 = 3'h3 == state ? _GEN_4307 : valid_1_70; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5079 = 3'h3 == state ? _GEN_4308 : valid_1_71; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5080 = 3'h3 == state ? _GEN_4309 : valid_1_72; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5081 = 3'h3 == state ? _GEN_4310 : valid_1_73; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5082 = 3'h3 == state ? _GEN_4311 : valid_1_74; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5083 = 3'h3 == state ? _GEN_4312 : valid_1_75; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5084 = 3'h3 == state ? _GEN_4313 : valid_1_76; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5085 = 3'h3 == state ? _GEN_4314 : valid_1_77; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5086 = 3'h3 == state ? _GEN_4315 : valid_1_78; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5087 = 3'h3 == state ? _GEN_4316 : valid_1_79; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5088 = 3'h3 == state ? _GEN_4317 : valid_1_80; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5089 = 3'h3 == state ? _GEN_4318 : valid_1_81; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5090 = 3'h3 == state ? _GEN_4319 : valid_1_82; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5091 = 3'h3 == state ? _GEN_4320 : valid_1_83; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5092 = 3'h3 == state ? _GEN_4321 : valid_1_84; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5093 = 3'h3 == state ? _GEN_4322 : valid_1_85; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5094 = 3'h3 == state ? _GEN_4323 : valid_1_86; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5095 = 3'h3 == state ? _GEN_4324 : valid_1_87; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5096 = 3'h3 == state ? _GEN_4325 : valid_1_88; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5097 = 3'h3 == state ? _GEN_4326 : valid_1_89; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5098 = 3'h3 == state ? _GEN_4327 : valid_1_90; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5099 = 3'h3 == state ? _GEN_4328 : valid_1_91; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5100 = 3'h3 == state ? _GEN_4329 : valid_1_92; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5101 = 3'h3 == state ? _GEN_4330 : valid_1_93; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5102 = 3'h3 == state ? _GEN_4331 : valid_1_94; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5103 = 3'h3 == state ? _GEN_4332 : valid_1_95; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5104 = 3'h3 == state ? _GEN_4333 : valid_1_96; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5105 = 3'h3 == state ? _GEN_4334 : valid_1_97; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5106 = 3'h3 == state ? _GEN_4335 : valid_1_98; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5107 = 3'h3 == state ? _GEN_4336 : valid_1_99; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5108 = 3'h3 == state ? _GEN_4337 : valid_1_100; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5109 = 3'h3 == state ? _GEN_4338 : valid_1_101; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5110 = 3'h3 == state ? _GEN_4339 : valid_1_102; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5111 = 3'h3 == state ? _GEN_4340 : valid_1_103; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5112 = 3'h3 == state ? _GEN_4341 : valid_1_104; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5113 = 3'h3 == state ? _GEN_4342 : valid_1_105; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5114 = 3'h3 == state ? _GEN_4343 : valid_1_106; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5115 = 3'h3 == state ? _GEN_4344 : valid_1_107; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5116 = 3'h3 == state ? _GEN_4345 : valid_1_108; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5117 = 3'h3 == state ? _GEN_4346 : valid_1_109; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5118 = 3'h3 == state ? _GEN_4347 : valid_1_110; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5119 = 3'h3 == state ? _GEN_4348 : valid_1_111; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5120 = 3'h3 == state ? _GEN_4349 : valid_1_112; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5121 = 3'h3 == state ? _GEN_4350 : valid_1_113; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5122 = 3'h3 == state ? _GEN_4351 : valid_1_114; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5123 = 3'h3 == state ? _GEN_4352 : valid_1_115; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5124 = 3'h3 == state ? _GEN_4353 : valid_1_116; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5125 = 3'h3 == state ? _GEN_4354 : valid_1_117; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5126 = 3'h3 == state ? _GEN_4355 : valid_1_118; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5127 = 3'h3 == state ? _GEN_4356 : valid_1_119; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5128 = 3'h3 == state ? _GEN_4357 : valid_1_120; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5129 = 3'h3 == state ? _GEN_4358 : valid_1_121; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5130 = 3'h3 == state ? _GEN_4359 : valid_1_122; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5131 = 3'h3 == state ? _GEN_4360 : valid_1_123; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5132 = 3'h3 == state ? _GEN_4361 : valid_1_124; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5133 = 3'h3 == state ? _GEN_4362 : valid_1_125; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5134 = 3'h3 == state ? _GEN_4363 : valid_1_126; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5135 = 3'h3 == state ? _GEN_4364 : valid_1_127; // @[i_cache.scala 55:18 22:26]
  wire [63:0] _GEN_7450 = 7'h1 == index ? ram_0_1 : ram_0_0; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7451 = 7'h2 == index ? ram_0_2 : _GEN_7450; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7452 = 7'h3 == index ? ram_0_3 : _GEN_7451; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7453 = 7'h4 == index ? ram_0_4 : _GEN_7452; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7454 = 7'h5 == index ? ram_0_5 : _GEN_7453; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7455 = 7'h6 == index ? ram_0_6 : _GEN_7454; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7456 = 7'h7 == index ? ram_0_7 : _GEN_7455; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7457 = 7'h8 == index ? ram_0_8 : _GEN_7456; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7458 = 7'h9 == index ? ram_0_9 : _GEN_7457; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7459 = 7'ha == index ? ram_0_10 : _GEN_7458; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7460 = 7'hb == index ? ram_0_11 : _GEN_7459; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7461 = 7'hc == index ? ram_0_12 : _GEN_7460; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7462 = 7'hd == index ? ram_0_13 : _GEN_7461; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7463 = 7'he == index ? ram_0_14 : _GEN_7462; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7464 = 7'hf == index ? ram_0_15 : _GEN_7463; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7465 = 7'h10 == index ? ram_0_16 : _GEN_7464; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7466 = 7'h11 == index ? ram_0_17 : _GEN_7465; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7467 = 7'h12 == index ? ram_0_18 : _GEN_7466; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7468 = 7'h13 == index ? ram_0_19 : _GEN_7467; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7469 = 7'h14 == index ? ram_0_20 : _GEN_7468; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7470 = 7'h15 == index ? ram_0_21 : _GEN_7469; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7471 = 7'h16 == index ? ram_0_22 : _GEN_7470; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7472 = 7'h17 == index ? ram_0_23 : _GEN_7471; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7473 = 7'h18 == index ? ram_0_24 : _GEN_7472; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7474 = 7'h19 == index ? ram_0_25 : _GEN_7473; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7475 = 7'h1a == index ? ram_0_26 : _GEN_7474; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7476 = 7'h1b == index ? ram_0_27 : _GEN_7475; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7477 = 7'h1c == index ? ram_0_28 : _GEN_7476; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7478 = 7'h1d == index ? ram_0_29 : _GEN_7477; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7479 = 7'h1e == index ? ram_0_30 : _GEN_7478; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7480 = 7'h1f == index ? ram_0_31 : _GEN_7479; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7481 = 7'h20 == index ? ram_0_32 : _GEN_7480; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7482 = 7'h21 == index ? ram_0_33 : _GEN_7481; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7483 = 7'h22 == index ? ram_0_34 : _GEN_7482; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7484 = 7'h23 == index ? ram_0_35 : _GEN_7483; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7485 = 7'h24 == index ? ram_0_36 : _GEN_7484; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7486 = 7'h25 == index ? ram_0_37 : _GEN_7485; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7487 = 7'h26 == index ? ram_0_38 : _GEN_7486; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7488 = 7'h27 == index ? ram_0_39 : _GEN_7487; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7489 = 7'h28 == index ? ram_0_40 : _GEN_7488; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7490 = 7'h29 == index ? ram_0_41 : _GEN_7489; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7491 = 7'h2a == index ? ram_0_42 : _GEN_7490; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7492 = 7'h2b == index ? ram_0_43 : _GEN_7491; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7493 = 7'h2c == index ? ram_0_44 : _GEN_7492; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7494 = 7'h2d == index ? ram_0_45 : _GEN_7493; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7495 = 7'h2e == index ? ram_0_46 : _GEN_7494; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7496 = 7'h2f == index ? ram_0_47 : _GEN_7495; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7497 = 7'h30 == index ? ram_0_48 : _GEN_7496; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7498 = 7'h31 == index ? ram_0_49 : _GEN_7497; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7499 = 7'h32 == index ? ram_0_50 : _GEN_7498; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7500 = 7'h33 == index ? ram_0_51 : _GEN_7499; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7501 = 7'h34 == index ? ram_0_52 : _GEN_7500; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7502 = 7'h35 == index ? ram_0_53 : _GEN_7501; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7503 = 7'h36 == index ? ram_0_54 : _GEN_7502; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7504 = 7'h37 == index ? ram_0_55 : _GEN_7503; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7505 = 7'h38 == index ? ram_0_56 : _GEN_7504; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7506 = 7'h39 == index ? ram_0_57 : _GEN_7505; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7507 = 7'h3a == index ? ram_0_58 : _GEN_7506; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7508 = 7'h3b == index ? ram_0_59 : _GEN_7507; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7509 = 7'h3c == index ? ram_0_60 : _GEN_7508; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7510 = 7'h3d == index ? ram_0_61 : _GEN_7509; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7511 = 7'h3e == index ? ram_0_62 : _GEN_7510; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7512 = 7'h3f == index ? ram_0_63 : _GEN_7511; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7513 = 7'h40 == index ? ram_0_64 : _GEN_7512; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7514 = 7'h41 == index ? ram_0_65 : _GEN_7513; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7515 = 7'h42 == index ? ram_0_66 : _GEN_7514; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7516 = 7'h43 == index ? ram_0_67 : _GEN_7515; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7517 = 7'h44 == index ? ram_0_68 : _GEN_7516; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7518 = 7'h45 == index ? ram_0_69 : _GEN_7517; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7519 = 7'h46 == index ? ram_0_70 : _GEN_7518; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7520 = 7'h47 == index ? ram_0_71 : _GEN_7519; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7521 = 7'h48 == index ? ram_0_72 : _GEN_7520; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7522 = 7'h49 == index ? ram_0_73 : _GEN_7521; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7523 = 7'h4a == index ? ram_0_74 : _GEN_7522; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7524 = 7'h4b == index ? ram_0_75 : _GEN_7523; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7525 = 7'h4c == index ? ram_0_76 : _GEN_7524; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7526 = 7'h4d == index ? ram_0_77 : _GEN_7525; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7527 = 7'h4e == index ? ram_0_78 : _GEN_7526; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7528 = 7'h4f == index ? ram_0_79 : _GEN_7527; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7529 = 7'h50 == index ? ram_0_80 : _GEN_7528; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7530 = 7'h51 == index ? ram_0_81 : _GEN_7529; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7531 = 7'h52 == index ? ram_0_82 : _GEN_7530; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7532 = 7'h53 == index ? ram_0_83 : _GEN_7531; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7533 = 7'h54 == index ? ram_0_84 : _GEN_7532; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7534 = 7'h55 == index ? ram_0_85 : _GEN_7533; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7535 = 7'h56 == index ? ram_0_86 : _GEN_7534; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7536 = 7'h57 == index ? ram_0_87 : _GEN_7535; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7537 = 7'h58 == index ? ram_0_88 : _GEN_7536; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7538 = 7'h59 == index ? ram_0_89 : _GEN_7537; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7539 = 7'h5a == index ? ram_0_90 : _GEN_7538; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7540 = 7'h5b == index ? ram_0_91 : _GEN_7539; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7541 = 7'h5c == index ? ram_0_92 : _GEN_7540; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7542 = 7'h5d == index ? ram_0_93 : _GEN_7541; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7543 = 7'h5e == index ? ram_0_94 : _GEN_7542; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7544 = 7'h5f == index ? ram_0_95 : _GEN_7543; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7545 = 7'h60 == index ? ram_0_96 : _GEN_7544; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7546 = 7'h61 == index ? ram_0_97 : _GEN_7545; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7547 = 7'h62 == index ? ram_0_98 : _GEN_7546; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7548 = 7'h63 == index ? ram_0_99 : _GEN_7547; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7549 = 7'h64 == index ? ram_0_100 : _GEN_7548; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7550 = 7'h65 == index ? ram_0_101 : _GEN_7549; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7551 = 7'h66 == index ? ram_0_102 : _GEN_7550; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7552 = 7'h67 == index ? ram_0_103 : _GEN_7551; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7553 = 7'h68 == index ? ram_0_104 : _GEN_7552; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7554 = 7'h69 == index ? ram_0_105 : _GEN_7553; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7555 = 7'h6a == index ? ram_0_106 : _GEN_7554; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7556 = 7'h6b == index ? ram_0_107 : _GEN_7555; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7557 = 7'h6c == index ? ram_0_108 : _GEN_7556; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7558 = 7'h6d == index ? ram_0_109 : _GEN_7557; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7559 = 7'h6e == index ? ram_0_110 : _GEN_7558; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7560 = 7'h6f == index ? ram_0_111 : _GEN_7559; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7561 = 7'h70 == index ? ram_0_112 : _GEN_7560; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7562 = 7'h71 == index ? ram_0_113 : _GEN_7561; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7563 = 7'h72 == index ? ram_0_114 : _GEN_7562; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7564 = 7'h73 == index ? ram_0_115 : _GEN_7563; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7565 = 7'h74 == index ? ram_0_116 : _GEN_7564; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7566 = 7'h75 == index ? ram_0_117 : _GEN_7565; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7567 = 7'h76 == index ? ram_0_118 : _GEN_7566; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7568 = 7'h77 == index ? ram_0_119 : _GEN_7567; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7569 = 7'h78 == index ? ram_0_120 : _GEN_7568; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7570 = 7'h79 == index ? ram_0_121 : _GEN_7569; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7571 = 7'h7a == index ? ram_0_122 : _GEN_7570; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7572 = 7'h7b == index ? ram_0_123 : _GEN_7571; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7573 = 7'h7c == index ? ram_0_124 : _GEN_7572; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7574 = 7'h7d == index ? ram_0_125 : _GEN_7573; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7575 = 7'h7e == index ? ram_0_126 : _GEN_7574; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7576 = 7'h7f == index ? ram_0_127 : _GEN_7575; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7578 = 7'h1 == index ? ram_1_1 : ram_1_0; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7579 = 7'h2 == index ? ram_1_2 : _GEN_7578; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7580 = 7'h3 == index ? ram_1_3 : _GEN_7579; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7581 = 7'h4 == index ? ram_1_4 : _GEN_7580; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7582 = 7'h5 == index ? ram_1_5 : _GEN_7581; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7583 = 7'h6 == index ? ram_1_6 : _GEN_7582; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7584 = 7'h7 == index ? ram_1_7 : _GEN_7583; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7585 = 7'h8 == index ? ram_1_8 : _GEN_7584; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7586 = 7'h9 == index ? ram_1_9 : _GEN_7585; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7587 = 7'ha == index ? ram_1_10 : _GEN_7586; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7588 = 7'hb == index ? ram_1_11 : _GEN_7587; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7589 = 7'hc == index ? ram_1_12 : _GEN_7588; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7590 = 7'hd == index ? ram_1_13 : _GEN_7589; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7591 = 7'he == index ? ram_1_14 : _GEN_7590; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7592 = 7'hf == index ? ram_1_15 : _GEN_7591; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7593 = 7'h10 == index ? ram_1_16 : _GEN_7592; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7594 = 7'h11 == index ? ram_1_17 : _GEN_7593; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7595 = 7'h12 == index ? ram_1_18 : _GEN_7594; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7596 = 7'h13 == index ? ram_1_19 : _GEN_7595; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7597 = 7'h14 == index ? ram_1_20 : _GEN_7596; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7598 = 7'h15 == index ? ram_1_21 : _GEN_7597; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7599 = 7'h16 == index ? ram_1_22 : _GEN_7598; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7600 = 7'h17 == index ? ram_1_23 : _GEN_7599; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7601 = 7'h18 == index ? ram_1_24 : _GEN_7600; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7602 = 7'h19 == index ? ram_1_25 : _GEN_7601; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7603 = 7'h1a == index ? ram_1_26 : _GEN_7602; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7604 = 7'h1b == index ? ram_1_27 : _GEN_7603; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7605 = 7'h1c == index ? ram_1_28 : _GEN_7604; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7606 = 7'h1d == index ? ram_1_29 : _GEN_7605; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7607 = 7'h1e == index ? ram_1_30 : _GEN_7606; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7608 = 7'h1f == index ? ram_1_31 : _GEN_7607; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7609 = 7'h20 == index ? ram_1_32 : _GEN_7608; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7610 = 7'h21 == index ? ram_1_33 : _GEN_7609; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7611 = 7'h22 == index ? ram_1_34 : _GEN_7610; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7612 = 7'h23 == index ? ram_1_35 : _GEN_7611; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7613 = 7'h24 == index ? ram_1_36 : _GEN_7612; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7614 = 7'h25 == index ? ram_1_37 : _GEN_7613; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7615 = 7'h26 == index ? ram_1_38 : _GEN_7614; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7616 = 7'h27 == index ? ram_1_39 : _GEN_7615; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7617 = 7'h28 == index ? ram_1_40 : _GEN_7616; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7618 = 7'h29 == index ? ram_1_41 : _GEN_7617; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7619 = 7'h2a == index ? ram_1_42 : _GEN_7618; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7620 = 7'h2b == index ? ram_1_43 : _GEN_7619; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7621 = 7'h2c == index ? ram_1_44 : _GEN_7620; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7622 = 7'h2d == index ? ram_1_45 : _GEN_7621; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7623 = 7'h2e == index ? ram_1_46 : _GEN_7622; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7624 = 7'h2f == index ? ram_1_47 : _GEN_7623; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7625 = 7'h30 == index ? ram_1_48 : _GEN_7624; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7626 = 7'h31 == index ? ram_1_49 : _GEN_7625; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7627 = 7'h32 == index ? ram_1_50 : _GEN_7626; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7628 = 7'h33 == index ? ram_1_51 : _GEN_7627; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7629 = 7'h34 == index ? ram_1_52 : _GEN_7628; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7630 = 7'h35 == index ? ram_1_53 : _GEN_7629; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7631 = 7'h36 == index ? ram_1_54 : _GEN_7630; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7632 = 7'h37 == index ? ram_1_55 : _GEN_7631; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7633 = 7'h38 == index ? ram_1_56 : _GEN_7632; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7634 = 7'h39 == index ? ram_1_57 : _GEN_7633; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7635 = 7'h3a == index ? ram_1_58 : _GEN_7634; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7636 = 7'h3b == index ? ram_1_59 : _GEN_7635; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7637 = 7'h3c == index ? ram_1_60 : _GEN_7636; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7638 = 7'h3d == index ? ram_1_61 : _GEN_7637; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7639 = 7'h3e == index ? ram_1_62 : _GEN_7638; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7640 = 7'h3f == index ? ram_1_63 : _GEN_7639; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7641 = 7'h40 == index ? ram_1_64 : _GEN_7640; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7642 = 7'h41 == index ? ram_1_65 : _GEN_7641; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7643 = 7'h42 == index ? ram_1_66 : _GEN_7642; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7644 = 7'h43 == index ? ram_1_67 : _GEN_7643; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7645 = 7'h44 == index ? ram_1_68 : _GEN_7644; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7646 = 7'h45 == index ? ram_1_69 : _GEN_7645; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7647 = 7'h46 == index ? ram_1_70 : _GEN_7646; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7648 = 7'h47 == index ? ram_1_71 : _GEN_7647; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7649 = 7'h48 == index ? ram_1_72 : _GEN_7648; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7650 = 7'h49 == index ? ram_1_73 : _GEN_7649; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7651 = 7'h4a == index ? ram_1_74 : _GEN_7650; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7652 = 7'h4b == index ? ram_1_75 : _GEN_7651; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7653 = 7'h4c == index ? ram_1_76 : _GEN_7652; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7654 = 7'h4d == index ? ram_1_77 : _GEN_7653; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7655 = 7'h4e == index ? ram_1_78 : _GEN_7654; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7656 = 7'h4f == index ? ram_1_79 : _GEN_7655; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7657 = 7'h50 == index ? ram_1_80 : _GEN_7656; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7658 = 7'h51 == index ? ram_1_81 : _GEN_7657; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7659 = 7'h52 == index ? ram_1_82 : _GEN_7658; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7660 = 7'h53 == index ? ram_1_83 : _GEN_7659; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7661 = 7'h54 == index ? ram_1_84 : _GEN_7660; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7662 = 7'h55 == index ? ram_1_85 : _GEN_7661; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7663 = 7'h56 == index ? ram_1_86 : _GEN_7662; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7664 = 7'h57 == index ? ram_1_87 : _GEN_7663; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7665 = 7'h58 == index ? ram_1_88 : _GEN_7664; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7666 = 7'h59 == index ? ram_1_89 : _GEN_7665; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7667 = 7'h5a == index ? ram_1_90 : _GEN_7666; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7668 = 7'h5b == index ? ram_1_91 : _GEN_7667; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7669 = 7'h5c == index ? ram_1_92 : _GEN_7668; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7670 = 7'h5d == index ? ram_1_93 : _GEN_7669; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7671 = 7'h5e == index ? ram_1_94 : _GEN_7670; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7672 = 7'h5f == index ? ram_1_95 : _GEN_7671; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7673 = 7'h60 == index ? ram_1_96 : _GEN_7672; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7674 = 7'h61 == index ? ram_1_97 : _GEN_7673; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7675 = 7'h62 == index ? ram_1_98 : _GEN_7674; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7676 = 7'h63 == index ? ram_1_99 : _GEN_7675; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7677 = 7'h64 == index ? ram_1_100 : _GEN_7676; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7678 = 7'h65 == index ? ram_1_101 : _GEN_7677; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7679 = 7'h66 == index ? ram_1_102 : _GEN_7678; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7680 = 7'h67 == index ? ram_1_103 : _GEN_7679; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7681 = 7'h68 == index ? ram_1_104 : _GEN_7680; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7682 = 7'h69 == index ? ram_1_105 : _GEN_7681; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7683 = 7'h6a == index ? ram_1_106 : _GEN_7682; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7684 = 7'h6b == index ? ram_1_107 : _GEN_7683; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7685 = 7'h6c == index ? ram_1_108 : _GEN_7684; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7686 = 7'h6d == index ? ram_1_109 : _GEN_7685; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7687 = 7'h6e == index ? ram_1_110 : _GEN_7686; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7688 = 7'h6f == index ? ram_1_111 : _GEN_7687; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7689 = 7'h70 == index ? ram_1_112 : _GEN_7688; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7690 = 7'h71 == index ? ram_1_113 : _GEN_7689; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7691 = 7'h72 == index ? ram_1_114 : _GEN_7690; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7692 = 7'h73 == index ? ram_1_115 : _GEN_7691; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7693 = 7'h74 == index ? ram_1_116 : _GEN_7692; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7694 = 7'h75 == index ? ram_1_117 : _GEN_7693; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7695 = 7'h76 == index ? ram_1_118 : _GEN_7694; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7696 = 7'h77 == index ? ram_1_119 : _GEN_7695; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7697 = 7'h78 == index ? ram_1_120 : _GEN_7696; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7698 = 7'h79 == index ? ram_1_121 : _GEN_7697; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7699 = 7'h7a == index ? ram_1_122 : _GEN_7698; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7700 = 7'h7b == index ? ram_1_123 : _GEN_7699; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7701 = 7'h7c == index ? ram_1_124 : _GEN_7700; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7702 = 7'h7d == index ? ram_1_125 : _GEN_7701; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7703 = 7'h7e == index ? ram_1_126 : _GEN_7702; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7704 = 7'h7f == index ? ram_1_127 : _GEN_7703; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7705 = way1_hit ? _GEN_7704 : 64'h0; // @[i_cache.scala 148:33 149:33 156:33]
  wire [63:0] _GEN_7709 = way0_hit ? _GEN_7576 : _GEN_7705; // @[i_cache.scala 140:23 141:33]
  wire  _GEN_7711 = way0_hit | way1_hit; // @[i_cache.scala 140:23 143:34]
  wire  _T_18 = state == 3'h2; // @[i_cache.scala 163:21]
  wire  _GEN_7722 = state == 3'h1 ? 1'h0 : _T_18; // @[i_cache.scala 130:31 131:27]
  wire  _GEN_7724 = state == 3'h1 ? 1'h0 : io_from_ifu_rready; // @[i_cache.scala 130:31 133:26]
  wire [63:0] _GEN_7726 = state == 3'h1 ? _GEN_7709 : 64'h0; // @[i_cache.scala 130:31]
  wire  _GEN_7728 = state == 3'h1 & _GEN_7711; // @[i_cache.scala 130:31]
  assign io_to_ifu_rdata = state == 3'h0 ? 64'h0 : _GEN_7726; // @[i_cache.scala 114:23 115:25]
  assign io_to_ifu_rvalid = state == 3'h0 ? 1'h0 : _GEN_7728; // @[i_cache.scala 114:23 117:26]
  assign io_to_axi_araddr = io_from_ifu_araddr; // @[i_cache.scala 114:23 122:26]
  assign io_to_axi_arvalid = state == 3'h0 ? 1'h0 : _GEN_7722; // @[i_cache.scala 114:23 121:27]
  assign io_to_axi_rready = state == 3'h0 ? io_from_ifu_rready : _GEN_7724; // @[i_cache.scala 114:23 123:26]
  always @(posedge clock) begin
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_0 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_0 <= _GEN_4367;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_1 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_1 <= _GEN_4368;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_2 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_2 <= _GEN_4369;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_3 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_3 <= _GEN_4370;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_4 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_4 <= _GEN_4371;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_5 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_5 <= _GEN_4372;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_6 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_6 <= _GEN_4373;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_7 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_7 <= _GEN_4374;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_8 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_8 <= _GEN_4375;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_9 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_9 <= _GEN_4376;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_10 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_10 <= _GEN_4377;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_11 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_11 <= _GEN_4378;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_12 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_12 <= _GEN_4379;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_13 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_13 <= _GEN_4380;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_14 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_14 <= _GEN_4381;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_15 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_15 <= _GEN_4382;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_16 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_16 <= _GEN_4383;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_17 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_17 <= _GEN_4384;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_18 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_18 <= _GEN_4385;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_19 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_19 <= _GEN_4386;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_20 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_20 <= _GEN_4387;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_21 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_21 <= _GEN_4388;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_22 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_22 <= _GEN_4389;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_23 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_23 <= _GEN_4390;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_24 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_24 <= _GEN_4391;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_25 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_25 <= _GEN_4392;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_26 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_26 <= _GEN_4393;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_27 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_27 <= _GEN_4394;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_28 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_28 <= _GEN_4395;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_29 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_29 <= _GEN_4396;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_30 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_30 <= _GEN_4397;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_31 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_31 <= _GEN_4398;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_32 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_32 <= _GEN_4399;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_33 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_33 <= _GEN_4400;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_34 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_34 <= _GEN_4401;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_35 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_35 <= _GEN_4402;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_36 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_36 <= _GEN_4403;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_37 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_37 <= _GEN_4404;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_38 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_38 <= _GEN_4405;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_39 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_39 <= _GEN_4406;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_40 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_40 <= _GEN_4407;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_41 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_41 <= _GEN_4408;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_42 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_42 <= _GEN_4409;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_43 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_43 <= _GEN_4410;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_44 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_44 <= _GEN_4411;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_45 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_45 <= _GEN_4412;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_46 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_46 <= _GEN_4413;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_47 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_47 <= _GEN_4414;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_48 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_48 <= _GEN_4415;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_49 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_49 <= _GEN_4416;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_50 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_50 <= _GEN_4417;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_51 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_51 <= _GEN_4418;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_52 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_52 <= _GEN_4419;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_53 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_53 <= _GEN_4420;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_54 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_54 <= _GEN_4421;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_55 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_55 <= _GEN_4422;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_56 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_56 <= _GEN_4423;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_57 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_57 <= _GEN_4424;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_58 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_58 <= _GEN_4425;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_59 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_59 <= _GEN_4426;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_60 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_60 <= _GEN_4427;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_61 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_61 <= _GEN_4428;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_62 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_62 <= _GEN_4429;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_63 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_63 <= _GEN_4430;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_64 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_64 <= _GEN_4431;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_65 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_65 <= _GEN_4432;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_66 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_66 <= _GEN_4433;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_67 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_67 <= _GEN_4434;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_68 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_68 <= _GEN_4435;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_69 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_69 <= _GEN_4436;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_70 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_70 <= _GEN_4437;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_71 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_71 <= _GEN_4438;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_72 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_72 <= _GEN_4439;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_73 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_73 <= _GEN_4440;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_74 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_74 <= _GEN_4441;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_75 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_75 <= _GEN_4442;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_76 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_76 <= _GEN_4443;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_77 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_77 <= _GEN_4444;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_78 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_78 <= _GEN_4445;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_79 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_79 <= _GEN_4446;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_80 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_80 <= _GEN_4447;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_81 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_81 <= _GEN_4448;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_82 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_82 <= _GEN_4449;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_83 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_83 <= _GEN_4450;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_84 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_84 <= _GEN_4451;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_85 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_85 <= _GEN_4452;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_86 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_86 <= _GEN_4453;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_87 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_87 <= _GEN_4454;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_88 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_88 <= _GEN_4455;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_89 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_89 <= _GEN_4456;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_90 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_90 <= _GEN_4457;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_91 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_91 <= _GEN_4458;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_92 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_92 <= _GEN_4459;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_93 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_93 <= _GEN_4460;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_94 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_94 <= _GEN_4461;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_95 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_95 <= _GEN_4462;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_96 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_96 <= _GEN_4463;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_97 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_97 <= _GEN_4464;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_98 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_98 <= _GEN_4465;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_99 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_99 <= _GEN_4466;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_100 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_100 <= _GEN_4467;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_101 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_101 <= _GEN_4468;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_102 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_102 <= _GEN_4469;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_103 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_103 <= _GEN_4470;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_104 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_104 <= _GEN_4471;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_105 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_105 <= _GEN_4472;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_106 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_106 <= _GEN_4473;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_107 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_107 <= _GEN_4474;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_108 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_108 <= _GEN_4475;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_109 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_109 <= _GEN_4476;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_110 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_110 <= _GEN_4477;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_111 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_111 <= _GEN_4478;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_112 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_112 <= _GEN_4479;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_113 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_113 <= _GEN_4480;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_114 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_114 <= _GEN_4481;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_115 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_115 <= _GEN_4482;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_116 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_116 <= _GEN_4483;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_117 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_117 <= _GEN_4484;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_118 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_118 <= _GEN_4485;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_119 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_119 <= _GEN_4486;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_120 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_120 <= _GEN_4487;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_121 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_121 <= _GEN_4488;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_122 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_122 <= _GEN_4489;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_123 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_123 <= _GEN_4490;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_124 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_124 <= _GEN_4491;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_125 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_125 <= _GEN_4492;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_126 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_126 <= _GEN_4493;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_127 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_127 <= _GEN_4494;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_0 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_0 <= _GEN_4752;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_1 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_1 <= _GEN_4753;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_2 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_2 <= _GEN_4754;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_3 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_3 <= _GEN_4755;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_4 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_4 <= _GEN_4756;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_5 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_5 <= _GEN_4757;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_6 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_6 <= _GEN_4758;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_7 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_7 <= _GEN_4759;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_8 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_8 <= _GEN_4760;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_9 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_9 <= _GEN_4761;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_10 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_10 <= _GEN_4762;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_11 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_11 <= _GEN_4763;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_12 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_12 <= _GEN_4764;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_13 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_13 <= _GEN_4765;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_14 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_14 <= _GEN_4766;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_15 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_15 <= _GEN_4767;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_16 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_16 <= _GEN_4768;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_17 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_17 <= _GEN_4769;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_18 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_18 <= _GEN_4770;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_19 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_19 <= _GEN_4771;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_20 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_20 <= _GEN_4772;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_21 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_21 <= _GEN_4773;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_22 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_22 <= _GEN_4774;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_23 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_23 <= _GEN_4775;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_24 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_24 <= _GEN_4776;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_25 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_25 <= _GEN_4777;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_26 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_26 <= _GEN_4778;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_27 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_27 <= _GEN_4779;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_28 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_28 <= _GEN_4780;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_29 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_29 <= _GEN_4781;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_30 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_30 <= _GEN_4782;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_31 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_31 <= _GEN_4783;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_32 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_32 <= _GEN_4784;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_33 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_33 <= _GEN_4785;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_34 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_34 <= _GEN_4786;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_35 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_35 <= _GEN_4787;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_36 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_36 <= _GEN_4788;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_37 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_37 <= _GEN_4789;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_38 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_38 <= _GEN_4790;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_39 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_39 <= _GEN_4791;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_40 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_40 <= _GEN_4792;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_41 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_41 <= _GEN_4793;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_42 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_42 <= _GEN_4794;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_43 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_43 <= _GEN_4795;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_44 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_44 <= _GEN_4796;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_45 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_45 <= _GEN_4797;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_46 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_46 <= _GEN_4798;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_47 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_47 <= _GEN_4799;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_48 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_48 <= _GEN_4800;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_49 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_49 <= _GEN_4801;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_50 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_50 <= _GEN_4802;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_51 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_51 <= _GEN_4803;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_52 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_52 <= _GEN_4804;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_53 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_53 <= _GEN_4805;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_54 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_54 <= _GEN_4806;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_55 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_55 <= _GEN_4807;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_56 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_56 <= _GEN_4808;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_57 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_57 <= _GEN_4809;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_58 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_58 <= _GEN_4810;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_59 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_59 <= _GEN_4811;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_60 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_60 <= _GEN_4812;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_61 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_61 <= _GEN_4813;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_62 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_62 <= _GEN_4814;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_63 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_63 <= _GEN_4815;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_64 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_64 <= _GEN_4816;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_65 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_65 <= _GEN_4817;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_66 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_66 <= _GEN_4818;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_67 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_67 <= _GEN_4819;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_68 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_68 <= _GEN_4820;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_69 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_69 <= _GEN_4821;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_70 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_70 <= _GEN_4822;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_71 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_71 <= _GEN_4823;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_72 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_72 <= _GEN_4824;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_73 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_73 <= _GEN_4825;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_74 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_74 <= _GEN_4826;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_75 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_75 <= _GEN_4827;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_76 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_76 <= _GEN_4828;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_77 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_77 <= _GEN_4829;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_78 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_78 <= _GEN_4830;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_79 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_79 <= _GEN_4831;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_80 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_80 <= _GEN_4832;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_81 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_81 <= _GEN_4833;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_82 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_82 <= _GEN_4834;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_83 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_83 <= _GEN_4835;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_84 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_84 <= _GEN_4836;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_85 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_85 <= _GEN_4837;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_86 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_86 <= _GEN_4838;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_87 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_87 <= _GEN_4839;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_88 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_88 <= _GEN_4840;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_89 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_89 <= _GEN_4841;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_90 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_90 <= _GEN_4842;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_91 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_91 <= _GEN_4843;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_92 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_92 <= _GEN_4844;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_93 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_93 <= _GEN_4845;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_94 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_94 <= _GEN_4846;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_95 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_95 <= _GEN_4847;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_96 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_96 <= _GEN_4848;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_97 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_97 <= _GEN_4849;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_98 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_98 <= _GEN_4850;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_99 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_99 <= _GEN_4851;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_100 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_100 <= _GEN_4852;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_101 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_101 <= _GEN_4853;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_102 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_102 <= _GEN_4854;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_103 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_103 <= _GEN_4855;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_104 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_104 <= _GEN_4856;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_105 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_105 <= _GEN_4857;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_106 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_106 <= _GEN_4858;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_107 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_107 <= _GEN_4859;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_108 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_108 <= _GEN_4860;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_109 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_109 <= _GEN_4861;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_110 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_110 <= _GEN_4862;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_111 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_111 <= _GEN_4863;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_112 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_112 <= _GEN_4864;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_113 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_113 <= _GEN_4865;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_114 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_114 <= _GEN_4866;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_115 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_115 <= _GEN_4867;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_116 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_116 <= _GEN_4868;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_117 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_117 <= _GEN_4869;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_118 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_118 <= _GEN_4870;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_119 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_119 <= _GEN_4871;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_120 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_120 <= _GEN_4872;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_121 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_121 <= _GEN_4873;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_122 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_122 <= _GEN_4874;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_123 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_123 <= _GEN_4875;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_124 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_124 <= _GEN_4876;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_125 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_125 <= _GEN_4877;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_126 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_126 <= _GEN_4878;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_127 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_127 <= _GEN_4879;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_0 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_0 <= _GEN_4495;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_1 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_1 <= _GEN_4496;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_2 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_2 <= _GEN_4497;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_3 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_3 <= _GEN_4498;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_4 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_4 <= _GEN_4499;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_5 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_5 <= _GEN_4500;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_6 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_6 <= _GEN_4501;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_7 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_7 <= _GEN_4502;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_8 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_8 <= _GEN_4503;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_9 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_9 <= _GEN_4504;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_10 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_10 <= _GEN_4505;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_11 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_11 <= _GEN_4506;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_12 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_12 <= _GEN_4507;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_13 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_13 <= _GEN_4508;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_14 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_14 <= _GEN_4509;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_15 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_15 <= _GEN_4510;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_16 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_16 <= _GEN_4511;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_17 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_17 <= _GEN_4512;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_18 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_18 <= _GEN_4513;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_19 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_19 <= _GEN_4514;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_20 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_20 <= _GEN_4515;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_21 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_21 <= _GEN_4516;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_22 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_22 <= _GEN_4517;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_23 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_23 <= _GEN_4518;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_24 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_24 <= _GEN_4519;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_25 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_25 <= _GEN_4520;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_26 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_26 <= _GEN_4521;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_27 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_27 <= _GEN_4522;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_28 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_28 <= _GEN_4523;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_29 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_29 <= _GEN_4524;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_30 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_30 <= _GEN_4525;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_31 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_31 <= _GEN_4526;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_32 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_32 <= _GEN_4527;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_33 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_33 <= _GEN_4528;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_34 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_34 <= _GEN_4529;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_35 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_35 <= _GEN_4530;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_36 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_36 <= _GEN_4531;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_37 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_37 <= _GEN_4532;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_38 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_38 <= _GEN_4533;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_39 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_39 <= _GEN_4534;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_40 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_40 <= _GEN_4535;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_41 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_41 <= _GEN_4536;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_42 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_42 <= _GEN_4537;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_43 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_43 <= _GEN_4538;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_44 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_44 <= _GEN_4539;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_45 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_45 <= _GEN_4540;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_46 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_46 <= _GEN_4541;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_47 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_47 <= _GEN_4542;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_48 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_48 <= _GEN_4543;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_49 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_49 <= _GEN_4544;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_50 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_50 <= _GEN_4545;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_51 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_51 <= _GEN_4546;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_52 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_52 <= _GEN_4547;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_53 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_53 <= _GEN_4548;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_54 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_54 <= _GEN_4549;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_55 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_55 <= _GEN_4550;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_56 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_56 <= _GEN_4551;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_57 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_57 <= _GEN_4552;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_58 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_58 <= _GEN_4553;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_59 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_59 <= _GEN_4554;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_60 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_60 <= _GEN_4555;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_61 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_61 <= _GEN_4556;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_62 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_62 <= _GEN_4557;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_63 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_63 <= _GEN_4558;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_64 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_64 <= _GEN_4559;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_65 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_65 <= _GEN_4560;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_66 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_66 <= _GEN_4561;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_67 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_67 <= _GEN_4562;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_68 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_68 <= _GEN_4563;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_69 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_69 <= _GEN_4564;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_70 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_70 <= _GEN_4565;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_71 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_71 <= _GEN_4566;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_72 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_72 <= _GEN_4567;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_73 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_73 <= _GEN_4568;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_74 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_74 <= _GEN_4569;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_75 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_75 <= _GEN_4570;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_76 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_76 <= _GEN_4571;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_77 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_77 <= _GEN_4572;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_78 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_78 <= _GEN_4573;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_79 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_79 <= _GEN_4574;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_80 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_80 <= _GEN_4575;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_81 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_81 <= _GEN_4576;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_82 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_82 <= _GEN_4577;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_83 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_83 <= _GEN_4578;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_84 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_84 <= _GEN_4579;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_85 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_85 <= _GEN_4580;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_86 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_86 <= _GEN_4581;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_87 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_87 <= _GEN_4582;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_88 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_88 <= _GEN_4583;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_89 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_89 <= _GEN_4584;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_90 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_90 <= _GEN_4585;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_91 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_91 <= _GEN_4586;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_92 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_92 <= _GEN_4587;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_93 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_93 <= _GEN_4588;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_94 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_94 <= _GEN_4589;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_95 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_95 <= _GEN_4590;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_96 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_96 <= _GEN_4591;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_97 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_97 <= _GEN_4592;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_98 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_98 <= _GEN_4593;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_99 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_99 <= _GEN_4594;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_100 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_100 <= _GEN_4595;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_101 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_101 <= _GEN_4596;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_102 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_102 <= _GEN_4597;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_103 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_103 <= _GEN_4598;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_104 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_104 <= _GEN_4599;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_105 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_105 <= _GEN_4600;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_106 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_106 <= _GEN_4601;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_107 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_107 <= _GEN_4602;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_108 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_108 <= _GEN_4603;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_109 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_109 <= _GEN_4604;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_110 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_110 <= _GEN_4605;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_111 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_111 <= _GEN_4606;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_112 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_112 <= _GEN_4607;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_113 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_113 <= _GEN_4608;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_114 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_114 <= _GEN_4609;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_115 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_115 <= _GEN_4610;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_116 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_116 <= _GEN_4611;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_117 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_117 <= _GEN_4612;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_118 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_118 <= _GEN_4613;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_119 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_119 <= _GEN_4614;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_120 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_120 <= _GEN_4615;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_121 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_121 <= _GEN_4616;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_122 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_122 <= _GEN_4617;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_123 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_123 <= _GEN_4618;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_124 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_124 <= _GEN_4619;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_125 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_125 <= _GEN_4620;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_126 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_126 <= _GEN_4621;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_127 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_127 <= _GEN_4622;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_0 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_0 <= _GEN_4880;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_1 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_1 <= _GEN_4881;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_2 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_2 <= _GEN_4882;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_3 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_3 <= _GEN_4883;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_4 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_4 <= _GEN_4884;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_5 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_5 <= _GEN_4885;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_6 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_6 <= _GEN_4886;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_7 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_7 <= _GEN_4887;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_8 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_8 <= _GEN_4888;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_9 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_9 <= _GEN_4889;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_10 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_10 <= _GEN_4890;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_11 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_11 <= _GEN_4891;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_12 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_12 <= _GEN_4892;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_13 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_13 <= _GEN_4893;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_14 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_14 <= _GEN_4894;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_15 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_15 <= _GEN_4895;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_16 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_16 <= _GEN_4896;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_17 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_17 <= _GEN_4897;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_18 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_18 <= _GEN_4898;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_19 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_19 <= _GEN_4899;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_20 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_20 <= _GEN_4900;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_21 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_21 <= _GEN_4901;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_22 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_22 <= _GEN_4902;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_23 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_23 <= _GEN_4903;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_24 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_24 <= _GEN_4904;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_25 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_25 <= _GEN_4905;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_26 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_26 <= _GEN_4906;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_27 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_27 <= _GEN_4907;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_28 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_28 <= _GEN_4908;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_29 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_29 <= _GEN_4909;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_30 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_30 <= _GEN_4910;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_31 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_31 <= _GEN_4911;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_32 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_32 <= _GEN_4912;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_33 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_33 <= _GEN_4913;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_34 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_34 <= _GEN_4914;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_35 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_35 <= _GEN_4915;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_36 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_36 <= _GEN_4916;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_37 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_37 <= _GEN_4917;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_38 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_38 <= _GEN_4918;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_39 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_39 <= _GEN_4919;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_40 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_40 <= _GEN_4920;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_41 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_41 <= _GEN_4921;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_42 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_42 <= _GEN_4922;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_43 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_43 <= _GEN_4923;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_44 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_44 <= _GEN_4924;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_45 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_45 <= _GEN_4925;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_46 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_46 <= _GEN_4926;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_47 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_47 <= _GEN_4927;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_48 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_48 <= _GEN_4928;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_49 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_49 <= _GEN_4929;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_50 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_50 <= _GEN_4930;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_51 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_51 <= _GEN_4931;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_52 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_52 <= _GEN_4932;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_53 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_53 <= _GEN_4933;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_54 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_54 <= _GEN_4934;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_55 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_55 <= _GEN_4935;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_56 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_56 <= _GEN_4936;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_57 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_57 <= _GEN_4937;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_58 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_58 <= _GEN_4938;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_59 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_59 <= _GEN_4939;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_60 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_60 <= _GEN_4940;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_61 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_61 <= _GEN_4941;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_62 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_62 <= _GEN_4942;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_63 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_63 <= _GEN_4943;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_64 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_64 <= _GEN_4944;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_65 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_65 <= _GEN_4945;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_66 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_66 <= _GEN_4946;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_67 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_67 <= _GEN_4947;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_68 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_68 <= _GEN_4948;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_69 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_69 <= _GEN_4949;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_70 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_70 <= _GEN_4950;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_71 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_71 <= _GEN_4951;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_72 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_72 <= _GEN_4952;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_73 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_73 <= _GEN_4953;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_74 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_74 <= _GEN_4954;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_75 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_75 <= _GEN_4955;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_76 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_76 <= _GEN_4956;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_77 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_77 <= _GEN_4957;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_78 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_78 <= _GEN_4958;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_79 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_79 <= _GEN_4959;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_80 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_80 <= _GEN_4960;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_81 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_81 <= _GEN_4961;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_82 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_82 <= _GEN_4962;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_83 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_83 <= _GEN_4963;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_84 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_84 <= _GEN_4964;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_85 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_85 <= _GEN_4965;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_86 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_86 <= _GEN_4966;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_87 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_87 <= _GEN_4967;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_88 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_88 <= _GEN_4968;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_89 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_89 <= _GEN_4969;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_90 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_90 <= _GEN_4970;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_91 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_91 <= _GEN_4971;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_92 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_92 <= _GEN_4972;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_93 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_93 <= _GEN_4973;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_94 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_94 <= _GEN_4974;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_95 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_95 <= _GEN_4975;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_96 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_96 <= _GEN_4976;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_97 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_97 <= _GEN_4977;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_98 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_98 <= _GEN_4978;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_99 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_99 <= _GEN_4979;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_100 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_100 <= _GEN_4980;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_101 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_101 <= _GEN_4981;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_102 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_102 <= _GEN_4982;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_103 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_103 <= _GEN_4983;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_104 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_104 <= _GEN_4984;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_105 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_105 <= _GEN_4985;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_106 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_106 <= _GEN_4986;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_107 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_107 <= _GEN_4987;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_108 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_108 <= _GEN_4988;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_109 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_109 <= _GEN_4989;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_110 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_110 <= _GEN_4990;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_111 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_111 <= _GEN_4991;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_112 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_112 <= _GEN_4992;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_113 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_113 <= _GEN_4993;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_114 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_114 <= _GEN_4994;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_115 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_115 <= _GEN_4995;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_116 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_116 <= _GEN_4996;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_117 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_117 <= _GEN_4997;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_118 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_118 <= _GEN_4998;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_119 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_119 <= _GEN_4999;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_120 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_120 <= _GEN_5000;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_121 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_121 <= _GEN_5001;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_122 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_122 <= _GEN_5002;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_123 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_123 <= _GEN_5003;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_124 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_124 <= _GEN_5004;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_125 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_125 <= _GEN_5005;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_126 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_126 <= _GEN_5006;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_127 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_127 <= _GEN_5007;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_0 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_0 <= _GEN_4623;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_1 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_1 <= _GEN_4624;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_2 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_2 <= _GEN_4625;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_3 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_3 <= _GEN_4626;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_4 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_4 <= _GEN_4627;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_5 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_5 <= _GEN_4628;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_6 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_6 <= _GEN_4629;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_7 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_7 <= _GEN_4630;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_8 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_8 <= _GEN_4631;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_9 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_9 <= _GEN_4632;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_10 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_10 <= _GEN_4633;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_11 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_11 <= _GEN_4634;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_12 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_12 <= _GEN_4635;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_13 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_13 <= _GEN_4636;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_14 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_14 <= _GEN_4637;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_15 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_15 <= _GEN_4638;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_16 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_16 <= _GEN_4639;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_17 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_17 <= _GEN_4640;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_18 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_18 <= _GEN_4641;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_19 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_19 <= _GEN_4642;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_20 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_20 <= _GEN_4643;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_21 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_21 <= _GEN_4644;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_22 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_22 <= _GEN_4645;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_23 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_23 <= _GEN_4646;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_24 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_24 <= _GEN_4647;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_25 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_25 <= _GEN_4648;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_26 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_26 <= _GEN_4649;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_27 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_27 <= _GEN_4650;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_28 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_28 <= _GEN_4651;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_29 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_29 <= _GEN_4652;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_30 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_30 <= _GEN_4653;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_31 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_31 <= _GEN_4654;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_32 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_32 <= _GEN_4655;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_33 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_33 <= _GEN_4656;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_34 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_34 <= _GEN_4657;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_35 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_35 <= _GEN_4658;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_36 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_36 <= _GEN_4659;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_37 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_37 <= _GEN_4660;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_38 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_38 <= _GEN_4661;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_39 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_39 <= _GEN_4662;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_40 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_40 <= _GEN_4663;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_41 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_41 <= _GEN_4664;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_42 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_42 <= _GEN_4665;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_43 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_43 <= _GEN_4666;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_44 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_44 <= _GEN_4667;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_45 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_45 <= _GEN_4668;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_46 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_46 <= _GEN_4669;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_47 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_47 <= _GEN_4670;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_48 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_48 <= _GEN_4671;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_49 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_49 <= _GEN_4672;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_50 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_50 <= _GEN_4673;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_51 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_51 <= _GEN_4674;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_52 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_52 <= _GEN_4675;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_53 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_53 <= _GEN_4676;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_54 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_54 <= _GEN_4677;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_55 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_55 <= _GEN_4678;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_56 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_56 <= _GEN_4679;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_57 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_57 <= _GEN_4680;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_58 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_58 <= _GEN_4681;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_59 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_59 <= _GEN_4682;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_60 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_60 <= _GEN_4683;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_61 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_61 <= _GEN_4684;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_62 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_62 <= _GEN_4685;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_63 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_63 <= _GEN_4686;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_64 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_64 <= _GEN_4687;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_65 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_65 <= _GEN_4688;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_66 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_66 <= _GEN_4689;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_67 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_67 <= _GEN_4690;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_68 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_68 <= _GEN_4691;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_69 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_69 <= _GEN_4692;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_70 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_70 <= _GEN_4693;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_71 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_71 <= _GEN_4694;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_72 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_72 <= _GEN_4695;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_73 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_73 <= _GEN_4696;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_74 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_74 <= _GEN_4697;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_75 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_75 <= _GEN_4698;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_76 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_76 <= _GEN_4699;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_77 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_77 <= _GEN_4700;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_78 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_78 <= _GEN_4701;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_79 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_79 <= _GEN_4702;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_80 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_80 <= _GEN_4703;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_81 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_81 <= _GEN_4704;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_82 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_82 <= _GEN_4705;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_83 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_83 <= _GEN_4706;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_84 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_84 <= _GEN_4707;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_85 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_85 <= _GEN_4708;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_86 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_86 <= _GEN_4709;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_87 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_87 <= _GEN_4710;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_88 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_88 <= _GEN_4711;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_89 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_89 <= _GEN_4712;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_90 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_90 <= _GEN_4713;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_91 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_91 <= _GEN_4714;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_92 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_92 <= _GEN_4715;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_93 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_93 <= _GEN_4716;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_94 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_94 <= _GEN_4717;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_95 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_95 <= _GEN_4718;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_96 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_96 <= _GEN_4719;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_97 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_97 <= _GEN_4720;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_98 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_98 <= _GEN_4721;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_99 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_99 <= _GEN_4722;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_100 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_100 <= _GEN_4723;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_101 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_101 <= _GEN_4724;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_102 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_102 <= _GEN_4725;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_103 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_103 <= _GEN_4726;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_104 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_104 <= _GEN_4727;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_105 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_105 <= _GEN_4728;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_106 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_106 <= _GEN_4729;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_107 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_107 <= _GEN_4730;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_108 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_108 <= _GEN_4731;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_109 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_109 <= _GEN_4732;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_110 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_110 <= _GEN_4733;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_111 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_111 <= _GEN_4734;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_112 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_112 <= _GEN_4735;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_113 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_113 <= _GEN_4736;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_114 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_114 <= _GEN_4737;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_115 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_115 <= _GEN_4738;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_116 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_116 <= _GEN_4739;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_117 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_117 <= _GEN_4740;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_118 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_118 <= _GEN_4741;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_119 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_119 <= _GEN_4742;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_120 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_120 <= _GEN_4743;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_121 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_121 <= _GEN_4744;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_122 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_122 <= _GEN_4745;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_123 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_123 <= _GEN_4746;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_124 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_124 <= _GEN_4747;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_125 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_125 <= _GEN_4748;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_126 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_126 <= _GEN_4749;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_127 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_127 <= _GEN_4750;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_0 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_0 <= _GEN_5008;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_1 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_1 <= _GEN_5009;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_2 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_2 <= _GEN_5010;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_3 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_3 <= _GEN_5011;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_4 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_4 <= _GEN_5012;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_5 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_5 <= _GEN_5013;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_6 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_6 <= _GEN_5014;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_7 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_7 <= _GEN_5015;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_8 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_8 <= _GEN_5016;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_9 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_9 <= _GEN_5017;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_10 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_10 <= _GEN_5018;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_11 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_11 <= _GEN_5019;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_12 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_12 <= _GEN_5020;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_13 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_13 <= _GEN_5021;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_14 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_14 <= _GEN_5022;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_15 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_15 <= _GEN_5023;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_16 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_16 <= _GEN_5024;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_17 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_17 <= _GEN_5025;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_18 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_18 <= _GEN_5026;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_19 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_19 <= _GEN_5027;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_20 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_20 <= _GEN_5028;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_21 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_21 <= _GEN_5029;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_22 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_22 <= _GEN_5030;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_23 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_23 <= _GEN_5031;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_24 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_24 <= _GEN_5032;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_25 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_25 <= _GEN_5033;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_26 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_26 <= _GEN_5034;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_27 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_27 <= _GEN_5035;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_28 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_28 <= _GEN_5036;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_29 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_29 <= _GEN_5037;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_30 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_30 <= _GEN_5038;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_31 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_31 <= _GEN_5039;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_32 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_32 <= _GEN_5040;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_33 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_33 <= _GEN_5041;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_34 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_34 <= _GEN_5042;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_35 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_35 <= _GEN_5043;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_36 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_36 <= _GEN_5044;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_37 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_37 <= _GEN_5045;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_38 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_38 <= _GEN_5046;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_39 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_39 <= _GEN_5047;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_40 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_40 <= _GEN_5048;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_41 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_41 <= _GEN_5049;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_42 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_42 <= _GEN_5050;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_43 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_43 <= _GEN_5051;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_44 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_44 <= _GEN_5052;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_45 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_45 <= _GEN_5053;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_46 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_46 <= _GEN_5054;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_47 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_47 <= _GEN_5055;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_48 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_48 <= _GEN_5056;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_49 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_49 <= _GEN_5057;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_50 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_50 <= _GEN_5058;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_51 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_51 <= _GEN_5059;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_52 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_52 <= _GEN_5060;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_53 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_53 <= _GEN_5061;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_54 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_54 <= _GEN_5062;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_55 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_55 <= _GEN_5063;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_56 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_56 <= _GEN_5064;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_57 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_57 <= _GEN_5065;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_58 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_58 <= _GEN_5066;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_59 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_59 <= _GEN_5067;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_60 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_60 <= _GEN_5068;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_61 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_61 <= _GEN_5069;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_62 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_62 <= _GEN_5070;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_63 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_63 <= _GEN_5071;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_64 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_64 <= _GEN_5072;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_65 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_65 <= _GEN_5073;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_66 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_66 <= _GEN_5074;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_67 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_67 <= _GEN_5075;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_68 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_68 <= _GEN_5076;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_69 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_69 <= _GEN_5077;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_70 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_70 <= _GEN_5078;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_71 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_71 <= _GEN_5079;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_72 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_72 <= _GEN_5080;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_73 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_73 <= _GEN_5081;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_74 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_74 <= _GEN_5082;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_75 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_75 <= _GEN_5083;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_76 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_76 <= _GEN_5084;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_77 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_77 <= _GEN_5085;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_78 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_78 <= _GEN_5086;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_79 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_79 <= _GEN_5087;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_80 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_80 <= _GEN_5088;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_81 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_81 <= _GEN_5089;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_82 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_82 <= _GEN_5090;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_83 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_83 <= _GEN_5091;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_84 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_84 <= _GEN_5092;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_85 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_85 <= _GEN_5093;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_86 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_86 <= _GEN_5094;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_87 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_87 <= _GEN_5095;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_88 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_88 <= _GEN_5096;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_89 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_89 <= _GEN_5097;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_90 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_90 <= _GEN_5098;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_91 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_91 <= _GEN_5099;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_92 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_92 <= _GEN_5100;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_93 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_93 <= _GEN_5101;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_94 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_94 <= _GEN_5102;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_95 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_95 <= _GEN_5103;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_96 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_96 <= _GEN_5104;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_97 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_97 <= _GEN_5105;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_98 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_98 <= _GEN_5106;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_99 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_99 <= _GEN_5107;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_100 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_100 <= _GEN_5108;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_101 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_101 <= _GEN_5109;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_102 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_102 <= _GEN_5110;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_103 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_103 <= _GEN_5111;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_104 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_104 <= _GEN_5112;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_105 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_105 <= _GEN_5113;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_106 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_106 <= _GEN_5114;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_107 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_107 <= _GEN_5115;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_108 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_108 <= _GEN_5116;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_109 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_109 <= _GEN_5117;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_110 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_110 <= _GEN_5118;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_111 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_111 <= _GEN_5119;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_112 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_112 <= _GEN_5120;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_113 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_113 <= _GEN_5121;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_114 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_114 <= _GEN_5122;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_115 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_115 <= _GEN_5123;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_116 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_116 <= _GEN_5124;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_117 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_117 <= _GEN_5125;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_118 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_118 <= _GEN_5126;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_119 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_119 <= _GEN_5127;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_120 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_120 <= _GEN_5128;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_121 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_121 <= _GEN_5129;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_122 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_122 <= _GEN_5130;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_123 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_123 <= _GEN_5131;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_124 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_124 <= _GEN_5132;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_125 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_125 <= _GEN_5133;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_126 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_126 <= _GEN_5134;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_127 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_127 <= _GEN_5135;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:27]
      way0_hit <= 1'h0; // @[i_cache.scala 23:27]
    end else begin
      way0_hit <= _T_2;
    end
    if (reset) begin // @[i_cache.scala 24:27]
      way1_hit <= 1'h0; // @[i_cache.scala 24:27]
    end else begin
      way1_hit <= _T_5;
    end
    if (reset) begin // @[i_cache.scala 26:28]
      unuse_way <= 2'h0; // @[i_cache.scala 26:28]
    end else if (~_GEN_255) begin // @[i_cache.scala 45:31]
      unuse_way <= 2'h1; // @[i_cache.scala 46:19]
    end else if (~_GEN_512) begin // @[i_cache.scala 47:37]
      unuse_way <= 2'h2; // @[i_cache.scala 48:19]
    end else begin
      unuse_way <= 2'h0; // @[i_cache.scala 50:19]
    end
    if (reset) begin // @[i_cache.scala 27:31]
      receive_data <= 64'h0; // @[i_cache.scala 27:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (3'h2 == state) begin // @[i_cache.scala 55:18]
          receive_data <= _GEN_521;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:24]
      quene <= 1'h0; // @[i_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          quene <= _GEN_4751;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 53:24]
      state <= 3'h0; // @[i_cache.scala 53:24]
    end else if (3'h0 == state) begin // @[i_cache.scala 55:18]
      if (io_from_ifu_arvalid) begin // @[i_cache.scala 57:38]
        state <= 3'h1; // @[i_cache.scala 58:23]
      end
    end else if (3'h1 == state) begin // @[i_cache.scala 55:18]
      if (way0_hit) begin // @[i_cache.scala 63:27]
        state <= _GEN_517;
      end else begin
        state <= _GEN_518;
      end
    end else if (3'h2 == state) begin // @[i_cache.scala 55:18]
      state <= _GEN_520;
    end else begin
      state <= _GEN_4366;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ram_0_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ram_0_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ram_0_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ram_0_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ram_0_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ram_0_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ram_0_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ram_0_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  ram_0_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  ram_0_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  ram_0_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  ram_0_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  ram_0_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  ram_0_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  ram_0_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  ram_0_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  ram_0_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  ram_0_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  ram_0_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  ram_0_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  ram_0_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  ram_0_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  ram_0_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  ram_0_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  ram_0_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  ram_0_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  ram_0_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  ram_0_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  ram_0_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  ram_0_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  ram_0_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  ram_0_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  ram_0_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  ram_0_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  ram_0_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  ram_0_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  ram_0_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  ram_0_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  ram_0_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  ram_0_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  ram_0_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  ram_0_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  ram_0_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  ram_0_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  ram_0_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  ram_0_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  ram_0_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  ram_0_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  ram_0_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  ram_0_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  ram_0_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  ram_0_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  ram_0_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  ram_0_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  ram_0_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  ram_0_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  ram_0_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  ram_0_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  ram_0_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  ram_0_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  ram_0_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  ram_0_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  ram_0_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  ram_0_63 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  ram_0_64 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  ram_0_65 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  ram_0_66 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  ram_0_67 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  ram_0_68 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  ram_0_69 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  ram_0_70 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  ram_0_71 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  ram_0_72 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  ram_0_73 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  ram_0_74 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  ram_0_75 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  ram_0_76 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  ram_0_77 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  ram_0_78 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  ram_0_79 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  ram_0_80 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  ram_0_81 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  ram_0_82 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  ram_0_83 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  ram_0_84 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  ram_0_85 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  ram_0_86 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  ram_0_87 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  ram_0_88 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  ram_0_89 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  ram_0_90 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  ram_0_91 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  ram_0_92 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  ram_0_93 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  ram_0_94 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  ram_0_95 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  ram_0_96 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  ram_0_97 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  ram_0_98 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  ram_0_99 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  ram_0_100 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  ram_0_101 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  ram_0_102 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  ram_0_103 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  ram_0_104 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  ram_0_105 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  ram_0_106 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  ram_0_107 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  ram_0_108 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  ram_0_109 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  ram_0_110 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  ram_0_111 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  ram_0_112 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  ram_0_113 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  ram_0_114 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  ram_0_115 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  ram_0_116 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  ram_0_117 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  ram_0_118 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  ram_0_119 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  ram_0_120 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  ram_0_121 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  ram_0_122 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  ram_0_123 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  ram_0_124 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  ram_0_125 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  ram_0_126 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  ram_0_127 = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  ram_1_0 = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  ram_1_1 = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  ram_1_2 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  ram_1_3 = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  ram_1_4 = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  ram_1_5 = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  ram_1_6 = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  ram_1_7 = _RAND_135[63:0];
  _RAND_136 = {2{`RANDOM}};
  ram_1_8 = _RAND_136[63:0];
  _RAND_137 = {2{`RANDOM}};
  ram_1_9 = _RAND_137[63:0];
  _RAND_138 = {2{`RANDOM}};
  ram_1_10 = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  ram_1_11 = _RAND_139[63:0];
  _RAND_140 = {2{`RANDOM}};
  ram_1_12 = _RAND_140[63:0];
  _RAND_141 = {2{`RANDOM}};
  ram_1_13 = _RAND_141[63:0];
  _RAND_142 = {2{`RANDOM}};
  ram_1_14 = _RAND_142[63:0];
  _RAND_143 = {2{`RANDOM}};
  ram_1_15 = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  ram_1_16 = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  ram_1_17 = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  ram_1_18 = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  ram_1_19 = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  ram_1_20 = _RAND_148[63:0];
  _RAND_149 = {2{`RANDOM}};
  ram_1_21 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  ram_1_22 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  ram_1_23 = _RAND_151[63:0];
  _RAND_152 = {2{`RANDOM}};
  ram_1_24 = _RAND_152[63:0];
  _RAND_153 = {2{`RANDOM}};
  ram_1_25 = _RAND_153[63:0];
  _RAND_154 = {2{`RANDOM}};
  ram_1_26 = _RAND_154[63:0];
  _RAND_155 = {2{`RANDOM}};
  ram_1_27 = _RAND_155[63:0];
  _RAND_156 = {2{`RANDOM}};
  ram_1_28 = _RAND_156[63:0];
  _RAND_157 = {2{`RANDOM}};
  ram_1_29 = _RAND_157[63:0];
  _RAND_158 = {2{`RANDOM}};
  ram_1_30 = _RAND_158[63:0];
  _RAND_159 = {2{`RANDOM}};
  ram_1_31 = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  ram_1_32 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  ram_1_33 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  ram_1_34 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  ram_1_35 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  ram_1_36 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  ram_1_37 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  ram_1_38 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  ram_1_39 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  ram_1_40 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  ram_1_41 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  ram_1_42 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  ram_1_43 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  ram_1_44 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  ram_1_45 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  ram_1_46 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  ram_1_47 = _RAND_175[63:0];
  _RAND_176 = {2{`RANDOM}};
  ram_1_48 = _RAND_176[63:0];
  _RAND_177 = {2{`RANDOM}};
  ram_1_49 = _RAND_177[63:0];
  _RAND_178 = {2{`RANDOM}};
  ram_1_50 = _RAND_178[63:0];
  _RAND_179 = {2{`RANDOM}};
  ram_1_51 = _RAND_179[63:0];
  _RAND_180 = {2{`RANDOM}};
  ram_1_52 = _RAND_180[63:0];
  _RAND_181 = {2{`RANDOM}};
  ram_1_53 = _RAND_181[63:0];
  _RAND_182 = {2{`RANDOM}};
  ram_1_54 = _RAND_182[63:0];
  _RAND_183 = {2{`RANDOM}};
  ram_1_55 = _RAND_183[63:0];
  _RAND_184 = {2{`RANDOM}};
  ram_1_56 = _RAND_184[63:0];
  _RAND_185 = {2{`RANDOM}};
  ram_1_57 = _RAND_185[63:0];
  _RAND_186 = {2{`RANDOM}};
  ram_1_58 = _RAND_186[63:0];
  _RAND_187 = {2{`RANDOM}};
  ram_1_59 = _RAND_187[63:0];
  _RAND_188 = {2{`RANDOM}};
  ram_1_60 = _RAND_188[63:0];
  _RAND_189 = {2{`RANDOM}};
  ram_1_61 = _RAND_189[63:0];
  _RAND_190 = {2{`RANDOM}};
  ram_1_62 = _RAND_190[63:0];
  _RAND_191 = {2{`RANDOM}};
  ram_1_63 = _RAND_191[63:0];
  _RAND_192 = {2{`RANDOM}};
  ram_1_64 = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  ram_1_65 = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  ram_1_66 = _RAND_194[63:0];
  _RAND_195 = {2{`RANDOM}};
  ram_1_67 = _RAND_195[63:0];
  _RAND_196 = {2{`RANDOM}};
  ram_1_68 = _RAND_196[63:0];
  _RAND_197 = {2{`RANDOM}};
  ram_1_69 = _RAND_197[63:0];
  _RAND_198 = {2{`RANDOM}};
  ram_1_70 = _RAND_198[63:0];
  _RAND_199 = {2{`RANDOM}};
  ram_1_71 = _RAND_199[63:0];
  _RAND_200 = {2{`RANDOM}};
  ram_1_72 = _RAND_200[63:0];
  _RAND_201 = {2{`RANDOM}};
  ram_1_73 = _RAND_201[63:0];
  _RAND_202 = {2{`RANDOM}};
  ram_1_74 = _RAND_202[63:0];
  _RAND_203 = {2{`RANDOM}};
  ram_1_75 = _RAND_203[63:0];
  _RAND_204 = {2{`RANDOM}};
  ram_1_76 = _RAND_204[63:0];
  _RAND_205 = {2{`RANDOM}};
  ram_1_77 = _RAND_205[63:0];
  _RAND_206 = {2{`RANDOM}};
  ram_1_78 = _RAND_206[63:0];
  _RAND_207 = {2{`RANDOM}};
  ram_1_79 = _RAND_207[63:0];
  _RAND_208 = {2{`RANDOM}};
  ram_1_80 = _RAND_208[63:0];
  _RAND_209 = {2{`RANDOM}};
  ram_1_81 = _RAND_209[63:0];
  _RAND_210 = {2{`RANDOM}};
  ram_1_82 = _RAND_210[63:0];
  _RAND_211 = {2{`RANDOM}};
  ram_1_83 = _RAND_211[63:0];
  _RAND_212 = {2{`RANDOM}};
  ram_1_84 = _RAND_212[63:0];
  _RAND_213 = {2{`RANDOM}};
  ram_1_85 = _RAND_213[63:0];
  _RAND_214 = {2{`RANDOM}};
  ram_1_86 = _RAND_214[63:0];
  _RAND_215 = {2{`RANDOM}};
  ram_1_87 = _RAND_215[63:0];
  _RAND_216 = {2{`RANDOM}};
  ram_1_88 = _RAND_216[63:0];
  _RAND_217 = {2{`RANDOM}};
  ram_1_89 = _RAND_217[63:0];
  _RAND_218 = {2{`RANDOM}};
  ram_1_90 = _RAND_218[63:0];
  _RAND_219 = {2{`RANDOM}};
  ram_1_91 = _RAND_219[63:0];
  _RAND_220 = {2{`RANDOM}};
  ram_1_92 = _RAND_220[63:0];
  _RAND_221 = {2{`RANDOM}};
  ram_1_93 = _RAND_221[63:0];
  _RAND_222 = {2{`RANDOM}};
  ram_1_94 = _RAND_222[63:0];
  _RAND_223 = {2{`RANDOM}};
  ram_1_95 = _RAND_223[63:0];
  _RAND_224 = {2{`RANDOM}};
  ram_1_96 = _RAND_224[63:0];
  _RAND_225 = {2{`RANDOM}};
  ram_1_97 = _RAND_225[63:0];
  _RAND_226 = {2{`RANDOM}};
  ram_1_98 = _RAND_226[63:0];
  _RAND_227 = {2{`RANDOM}};
  ram_1_99 = _RAND_227[63:0];
  _RAND_228 = {2{`RANDOM}};
  ram_1_100 = _RAND_228[63:0];
  _RAND_229 = {2{`RANDOM}};
  ram_1_101 = _RAND_229[63:0];
  _RAND_230 = {2{`RANDOM}};
  ram_1_102 = _RAND_230[63:0];
  _RAND_231 = {2{`RANDOM}};
  ram_1_103 = _RAND_231[63:0];
  _RAND_232 = {2{`RANDOM}};
  ram_1_104 = _RAND_232[63:0];
  _RAND_233 = {2{`RANDOM}};
  ram_1_105 = _RAND_233[63:0];
  _RAND_234 = {2{`RANDOM}};
  ram_1_106 = _RAND_234[63:0];
  _RAND_235 = {2{`RANDOM}};
  ram_1_107 = _RAND_235[63:0];
  _RAND_236 = {2{`RANDOM}};
  ram_1_108 = _RAND_236[63:0];
  _RAND_237 = {2{`RANDOM}};
  ram_1_109 = _RAND_237[63:0];
  _RAND_238 = {2{`RANDOM}};
  ram_1_110 = _RAND_238[63:0];
  _RAND_239 = {2{`RANDOM}};
  ram_1_111 = _RAND_239[63:0];
  _RAND_240 = {2{`RANDOM}};
  ram_1_112 = _RAND_240[63:0];
  _RAND_241 = {2{`RANDOM}};
  ram_1_113 = _RAND_241[63:0];
  _RAND_242 = {2{`RANDOM}};
  ram_1_114 = _RAND_242[63:0];
  _RAND_243 = {2{`RANDOM}};
  ram_1_115 = _RAND_243[63:0];
  _RAND_244 = {2{`RANDOM}};
  ram_1_116 = _RAND_244[63:0];
  _RAND_245 = {2{`RANDOM}};
  ram_1_117 = _RAND_245[63:0];
  _RAND_246 = {2{`RANDOM}};
  ram_1_118 = _RAND_246[63:0];
  _RAND_247 = {2{`RANDOM}};
  ram_1_119 = _RAND_247[63:0];
  _RAND_248 = {2{`RANDOM}};
  ram_1_120 = _RAND_248[63:0];
  _RAND_249 = {2{`RANDOM}};
  ram_1_121 = _RAND_249[63:0];
  _RAND_250 = {2{`RANDOM}};
  ram_1_122 = _RAND_250[63:0];
  _RAND_251 = {2{`RANDOM}};
  ram_1_123 = _RAND_251[63:0];
  _RAND_252 = {2{`RANDOM}};
  ram_1_124 = _RAND_252[63:0];
  _RAND_253 = {2{`RANDOM}};
  ram_1_125 = _RAND_253[63:0];
  _RAND_254 = {2{`RANDOM}};
  ram_1_126 = _RAND_254[63:0];
  _RAND_255 = {2{`RANDOM}};
  ram_1_127 = _RAND_255[63:0];
  _RAND_256 = {1{`RANDOM}};
  tag_0_0 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  tag_0_1 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  tag_0_2 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  tag_0_3 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  tag_0_4 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  tag_0_5 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  tag_0_6 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  tag_0_7 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  tag_0_8 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  tag_0_9 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  tag_0_10 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  tag_0_11 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  tag_0_12 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  tag_0_13 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  tag_0_14 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  tag_0_15 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  tag_0_16 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  tag_0_17 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  tag_0_18 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  tag_0_19 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  tag_0_20 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  tag_0_21 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  tag_0_22 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  tag_0_23 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  tag_0_24 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  tag_0_25 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  tag_0_26 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  tag_0_27 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  tag_0_28 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  tag_0_29 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  tag_0_30 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  tag_0_31 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  tag_0_32 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  tag_0_33 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  tag_0_34 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  tag_0_35 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  tag_0_36 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  tag_0_37 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  tag_0_38 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  tag_0_39 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  tag_0_40 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  tag_0_41 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  tag_0_42 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  tag_0_43 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  tag_0_44 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  tag_0_45 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  tag_0_46 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  tag_0_47 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  tag_0_48 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  tag_0_49 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  tag_0_50 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  tag_0_51 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  tag_0_52 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  tag_0_53 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  tag_0_54 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  tag_0_55 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  tag_0_56 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  tag_0_57 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  tag_0_58 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  tag_0_59 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  tag_0_60 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  tag_0_61 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  tag_0_62 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  tag_0_63 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  tag_0_64 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  tag_0_65 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  tag_0_66 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  tag_0_67 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  tag_0_68 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  tag_0_69 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  tag_0_70 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  tag_0_71 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  tag_0_72 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  tag_0_73 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  tag_0_74 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  tag_0_75 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  tag_0_76 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  tag_0_77 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  tag_0_78 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  tag_0_79 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  tag_0_80 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  tag_0_81 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  tag_0_82 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  tag_0_83 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  tag_0_84 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  tag_0_85 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  tag_0_86 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  tag_0_87 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  tag_0_88 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  tag_0_89 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  tag_0_90 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  tag_0_91 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  tag_0_92 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  tag_0_93 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  tag_0_94 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  tag_0_95 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  tag_0_96 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  tag_0_97 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  tag_0_98 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  tag_0_99 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  tag_0_100 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  tag_0_101 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  tag_0_102 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  tag_0_103 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  tag_0_104 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  tag_0_105 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  tag_0_106 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  tag_0_107 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  tag_0_108 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  tag_0_109 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  tag_0_110 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  tag_0_111 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  tag_0_112 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  tag_0_113 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  tag_0_114 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  tag_0_115 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  tag_0_116 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  tag_0_117 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  tag_0_118 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  tag_0_119 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  tag_0_120 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  tag_0_121 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  tag_0_122 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  tag_0_123 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  tag_0_124 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  tag_0_125 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  tag_0_126 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  tag_0_127 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  tag_1_0 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  tag_1_1 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  tag_1_2 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  tag_1_3 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  tag_1_4 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  tag_1_5 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  tag_1_6 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  tag_1_7 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  tag_1_8 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  tag_1_9 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  tag_1_10 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  tag_1_11 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  tag_1_12 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  tag_1_13 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  tag_1_14 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  tag_1_15 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  tag_1_16 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  tag_1_17 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  tag_1_18 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  tag_1_19 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  tag_1_20 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  tag_1_21 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  tag_1_22 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  tag_1_23 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  tag_1_24 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  tag_1_25 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  tag_1_26 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  tag_1_27 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  tag_1_28 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  tag_1_29 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  tag_1_30 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  tag_1_31 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  tag_1_32 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  tag_1_33 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  tag_1_34 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  tag_1_35 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  tag_1_36 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  tag_1_37 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  tag_1_38 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  tag_1_39 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  tag_1_40 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  tag_1_41 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  tag_1_42 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  tag_1_43 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  tag_1_44 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  tag_1_45 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  tag_1_46 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  tag_1_47 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  tag_1_48 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  tag_1_49 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  tag_1_50 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  tag_1_51 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  tag_1_52 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  tag_1_53 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  tag_1_54 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  tag_1_55 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  tag_1_56 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  tag_1_57 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  tag_1_58 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  tag_1_59 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  tag_1_60 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  tag_1_61 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  tag_1_62 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  tag_1_63 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  tag_1_64 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  tag_1_65 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  tag_1_66 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  tag_1_67 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  tag_1_68 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  tag_1_69 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  tag_1_70 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  tag_1_71 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  tag_1_72 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  tag_1_73 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  tag_1_74 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  tag_1_75 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  tag_1_76 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  tag_1_77 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  tag_1_78 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  tag_1_79 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  tag_1_80 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  tag_1_81 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  tag_1_82 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  tag_1_83 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  tag_1_84 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  tag_1_85 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  tag_1_86 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  tag_1_87 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  tag_1_88 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  tag_1_89 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  tag_1_90 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  tag_1_91 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  tag_1_92 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  tag_1_93 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  tag_1_94 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  tag_1_95 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  tag_1_96 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  tag_1_97 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  tag_1_98 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  tag_1_99 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  tag_1_100 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  tag_1_101 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  tag_1_102 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  tag_1_103 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  tag_1_104 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  tag_1_105 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  tag_1_106 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  tag_1_107 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  tag_1_108 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  tag_1_109 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  tag_1_110 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  tag_1_111 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  tag_1_112 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  tag_1_113 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  tag_1_114 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  tag_1_115 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  tag_1_116 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  tag_1_117 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  tag_1_118 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  tag_1_119 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  tag_1_120 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  tag_1_121 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  tag_1_122 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  tag_1_123 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  tag_1_124 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  tag_1_125 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  tag_1_126 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  tag_1_127 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  valid_0_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid_0_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  valid_0_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  valid_0_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  valid_0_4 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  valid_0_5 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  valid_0_6 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  valid_0_7 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  valid_0_8 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  valid_0_9 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  valid_0_10 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  valid_0_11 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  valid_0_12 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  valid_0_13 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  valid_0_14 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  valid_0_15 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  valid_0_16 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  valid_0_17 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  valid_0_18 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  valid_0_19 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  valid_0_20 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  valid_0_21 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  valid_0_22 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  valid_0_23 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  valid_0_24 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  valid_0_25 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  valid_0_26 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  valid_0_27 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  valid_0_28 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  valid_0_29 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  valid_0_30 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  valid_0_31 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  valid_0_32 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  valid_0_33 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  valid_0_34 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  valid_0_35 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  valid_0_36 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  valid_0_37 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  valid_0_38 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  valid_0_39 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  valid_0_40 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  valid_0_41 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  valid_0_42 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  valid_0_43 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  valid_0_44 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  valid_0_45 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  valid_0_46 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  valid_0_47 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  valid_0_48 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  valid_0_49 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  valid_0_50 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  valid_0_51 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  valid_0_52 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  valid_0_53 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  valid_0_54 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  valid_0_55 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  valid_0_56 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  valid_0_57 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  valid_0_58 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  valid_0_59 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  valid_0_60 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  valid_0_61 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  valid_0_62 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  valid_0_63 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  valid_0_64 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  valid_0_65 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  valid_0_66 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  valid_0_67 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  valid_0_68 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  valid_0_69 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  valid_0_70 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  valid_0_71 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  valid_0_72 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  valid_0_73 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  valid_0_74 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  valid_0_75 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  valid_0_76 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  valid_0_77 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  valid_0_78 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  valid_0_79 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  valid_0_80 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  valid_0_81 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  valid_0_82 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  valid_0_83 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  valid_0_84 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  valid_0_85 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  valid_0_86 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  valid_0_87 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  valid_0_88 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  valid_0_89 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  valid_0_90 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  valid_0_91 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  valid_0_92 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  valid_0_93 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  valid_0_94 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  valid_0_95 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  valid_0_96 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  valid_0_97 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  valid_0_98 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  valid_0_99 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  valid_0_100 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  valid_0_101 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  valid_0_102 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  valid_0_103 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  valid_0_104 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  valid_0_105 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  valid_0_106 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  valid_0_107 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  valid_0_108 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  valid_0_109 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  valid_0_110 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  valid_0_111 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  valid_0_112 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  valid_0_113 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  valid_0_114 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  valid_0_115 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  valid_0_116 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  valid_0_117 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  valid_0_118 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  valid_0_119 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  valid_0_120 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  valid_0_121 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  valid_0_122 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  valid_0_123 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  valid_0_124 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  valid_0_125 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  valid_0_126 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  valid_0_127 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  valid_1_0 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  valid_1_1 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  valid_1_2 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  valid_1_3 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  valid_1_4 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  valid_1_5 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  valid_1_6 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  valid_1_7 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  valid_1_8 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  valid_1_9 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  valid_1_10 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  valid_1_11 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  valid_1_12 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  valid_1_13 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  valid_1_14 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  valid_1_15 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  valid_1_16 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  valid_1_17 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  valid_1_18 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  valid_1_19 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  valid_1_20 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  valid_1_21 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  valid_1_22 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  valid_1_23 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  valid_1_24 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  valid_1_25 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  valid_1_26 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  valid_1_27 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  valid_1_28 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  valid_1_29 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  valid_1_30 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  valid_1_31 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  valid_1_32 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  valid_1_33 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  valid_1_34 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  valid_1_35 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  valid_1_36 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  valid_1_37 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  valid_1_38 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  valid_1_39 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  valid_1_40 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  valid_1_41 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  valid_1_42 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  valid_1_43 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  valid_1_44 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  valid_1_45 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  valid_1_46 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  valid_1_47 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  valid_1_48 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  valid_1_49 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  valid_1_50 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  valid_1_51 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  valid_1_52 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  valid_1_53 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  valid_1_54 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  valid_1_55 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  valid_1_56 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  valid_1_57 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  valid_1_58 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  valid_1_59 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  valid_1_60 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  valid_1_61 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  valid_1_62 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  valid_1_63 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  valid_1_64 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  valid_1_65 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  valid_1_66 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  valid_1_67 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  valid_1_68 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  valid_1_69 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  valid_1_70 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  valid_1_71 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  valid_1_72 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  valid_1_73 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  valid_1_74 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  valid_1_75 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  valid_1_76 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  valid_1_77 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  valid_1_78 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  valid_1_79 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  valid_1_80 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  valid_1_81 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  valid_1_82 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  valid_1_83 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  valid_1_84 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  valid_1_85 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  valid_1_86 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  valid_1_87 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  valid_1_88 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  valid_1_89 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  valid_1_90 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  valid_1_91 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  valid_1_92 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  valid_1_93 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  valid_1_94 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  valid_1_95 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  valid_1_96 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  valid_1_97 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  valid_1_98 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  valid_1_99 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  valid_1_100 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  valid_1_101 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  valid_1_102 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  valid_1_103 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  valid_1_104 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  valid_1_105 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  valid_1_106 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  valid_1_107 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  valid_1_108 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  valid_1_109 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  valid_1_110 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  valid_1_111 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  valid_1_112 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  valid_1_113 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  valid_1_114 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  valid_1_115 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  valid_1_116 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  valid_1_117 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  valid_1_118 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  valid_1_119 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  valid_1_120 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  valid_1_121 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  valid_1_122 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  valid_1_123 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  valid_1_124 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  valid_1_125 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  valid_1_126 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  valid_1_127 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  way0_hit = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  way1_hit = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  unuse_way = _RAND_770[1:0];
  _RAND_771 = {2{`RANDOM}};
  receive_data = _RAND_771[63:0];
  _RAND_772 = {1{`RANDOM}};
  quene = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  state = _RAND_773[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module D_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_lsu_araddr,
  input         io_from_lsu_arvalid,
  input         io_from_lsu_rready,
  input  [31:0] io_from_lsu_awaddr,
  input         io_from_lsu_awvalid,
  input  [31:0] io_from_lsu_wdata,
  input  [7:0]  io_from_lsu_wstrb,
  input         io_from_lsu_wvalid,
  input         io_from_lsu_bready,
  output        io_to_lsu_arready,
  output [63:0] io_to_lsu_rdata,
  output        io_to_lsu_rvalid,
  output        io_to_lsu_awready,
  output        io_to_lsu_wready,
  output        io_to_lsu_bvalid,
  output [31:0] io_to_axi_araddr,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  output [31:0] io_to_axi_awaddr,
  output        io_to_axi_awvalid,
  output [31:0] io_to_axi_wdata,
  output [7:0]  io_to_axi_wstrb,
  output        io_to_axi_wvalid,
  output        io_to_axi_bready,
  input         io_from_axi_arready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rvalid,
  input         io_from_axi_awready,
  input         io_from_axi_wready,
  input         io_from_axi_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [63:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [63:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = ~reset; // @[d_cache.scala 15:11]
  reg [63:0] ram_0_0; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_1; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_2; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_3; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_4; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_5; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_6; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_7; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_8; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_9; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_10; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_11; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_12; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_13; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_14; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_15; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_16; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_17; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_18; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_19; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_20; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_21; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_22; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_23; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_24; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_25; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_26; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_27; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_28; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_29; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_30; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_31; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_32; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_33; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_34; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_35; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_36; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_37; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_38; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_39; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_40; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_41; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_42; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_43; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_44; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_45; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_46; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_47; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_48; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_49; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_50; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_51; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_52; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_53; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_54; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_55; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_56; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_57; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_58; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_59; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_60; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_61; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_62; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_63; // @[d_cache.scala 18:24]
  reg [63:0] ram_1_0; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_1; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_2; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_3; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_4; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_5; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_6; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_7; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_8; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_9; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_10; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_11; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_12; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_13; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_14; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_15; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_16; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_17; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_18; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_19; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_20; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_21; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_22; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_23; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_24; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_25; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_26; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_27; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_28; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_29; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_30; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_31; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_32; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_33; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_34; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_35; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_36; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_37; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_38; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_39; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_40; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_41; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_42; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_43; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_44; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_45; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_46; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_47; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_48; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_49; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_50; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_51; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_52; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_53; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_54; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_55; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_56; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_57; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_58; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_59; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_60; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_61; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_62; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_63; // @[d_cache.scala 19:24]
  reg [31:0] tag_0_0; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_1; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_2; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_3; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_4; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_5; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_6; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_7; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_8; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_9; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_10; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_11; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_12; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_13; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_14; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_15; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_16; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_17; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_18; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_19; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_20; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_21; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_22; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_23; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_24; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_25; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_26; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_27; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_28; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_29; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_30; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_31; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_32; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_33; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_34; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_35; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_36; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_37; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_38; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_39; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_40; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_41; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_42; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_43; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_44; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_45; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_46; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_47; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_48; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_49; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_50; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_51; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_52; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_53; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_54; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_55; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_56; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_57; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_58; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_59; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_60; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_61; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_62; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_63; // @[d_cache.scala 22:24]
  reg [31:0] tag_1_0; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_1; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_2; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_3; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_4; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_5; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_6; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_7; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_8; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_9; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_10; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_11; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_12; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_13; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_14; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_15; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_16; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_17; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_18; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_19; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_20; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_21; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_22; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_23; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_24; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_25; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_26; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_27; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_28; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_29; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_30; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_31; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_32; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_33; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_34; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_35; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_36; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_37; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_38; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_39; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_40; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_41; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_42; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_43; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_44; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_45; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_46; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_47; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_48; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_49; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_50; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_51; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_52; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_53; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_54; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_55; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_56; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_57; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_58; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_59; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_60; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_61; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_62; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_63; // @[d_cache.scala 23:24]
  reg  valid_0_0; // @[d_cache.scala 24:26]
  reg  valid_0_1; // @[d_cache.scala 24:26]
  reg  valid_0_2; // @[d_cache.scala 24:26]
  reg  valid_0_3; // @[d_cache.scala 24:26]
  reg  valid_0_4; // @[d_cache.scala 24:26]
  reg  valid_0_5; // @[d_cache.scala 24:26]
  reg  valid_0_6; // @[d_cache.scala 24:26]
  reg  valid_0_7; // @[d_cache.scala 24:26]
  reg  valid_0_8; // @[d_cache.scala 24:26]
  reg  valid_0_9; // @[d_cache.scala 24:26]
  reg  valid_0_10; // @[d_cache.scala 24:26]
  reg  valid_0_11; // @[d_cache.scala 24:26]
  reg  valid_0_12; // @[d_cache.scala 24:26]
  reg  valid_0_13; // @[d_cache.scala 24:26]
  reg  valid_0_14; // @[d_cache.scala 24:26]
  reg  valid_0_15; // @[d_cache.scala 24:26]
  reg  valid_0_16; // @[d_cache.scala 24:26]
  reg  valid_0_17; // @[d_cache.scala 24:26]
  reg  valid_0_18; // @[d_cache.scala 24:26]
  reg  valid_0_19; // @[d_cache.scala 24:26]
  reg  valid_0_20; // @[d_cache.scala 24:26]
  reg  valid_0_21; // @[d_cache.scala 24:26]
  reg  valid_0_22; // @[d_cache.scala 24:26]
  reg  valid_0_23; // @[d_cache.scala 24:26]
  reg  valid_0_24; // @[d_cache.scala 24:26]
  reg  valid_0_25; // @[d_cache.scala 24:26]
  reg  valid_0_26; // @[d_cache.scala 24:26]
  reg  valid_0_27; // @[d_cache.scala 24:26]
  reg  valid_0_28; // @[d_cache.scala 24:26]
  reg  valid_0_29; // @[d_cache.scala 24:26]
  reg  valid_0_30; // @[d_cache.scala 24:26]
  reg  valid_0_31; // @[d_cache.scala 24:26]
  reg  valid_0_32; // @[d_cache.scala 24:26]
  reg  valid_0_33; // @[d_cache.scala 24:26]
  reg  valid_0_34; // @[d_cache.scala 24:26]
  reg  valid_0_35; // @[d_cache.scala 24:26]
  reg  valid_0_36; // @[d_cache.scala 24:26]
  reg  valid_0_37; // @[d_cache.scala 24:26]
  reg  valid_0_38; // @[d_cache.scala 24:26]
  reg  valid_0_39; // @[d_cache.scala 24:26]
  reg  valid_0_40; // @[d_cache.scala 24:26]
  reg  valid_0_41; // @[d_cache.scala 24:26]
  reg  valid_0_42; // @[d_cache.scala 24:26]
  reg  valid_0_43; // @[d_cache.scala 24:26]
  reg  valid_0_44; // @[d_cache.scala 24:26]
  reg  valid_0_45; // @[d_cache.scala 24:26]
  reg  valid_0_46; // @[d_cache.scala 24:26]
  reg  valid_0_47; // @[d_cache.scala 24:26]
  reg  valid_0_48; // @[d_cache.scala 24:26]
  reg  valid_0_49; // @[d_cache.scala 24:26]
  reg  valid_0_50; // @[d_cache.scala 24:26]
  reg  valid_0_51; // @[d_cache.scala 24:26]
  reg  valid_0_52; // @[d_cache.scala 24:26]
  reg  valid_0_53; // @[d_cache.scala 24:26]
  reg  valid_0_54; // @[d_cache.scala 24:26]
  reg  valid_0_55; // @[d_cache.scala 24:26]
  reg  valid_0_56; // @[d_cache.scala 24:26]
  reg  valid_0_57; // @[d_cache.scala 24:26]
  reg  valid_0_58; // @[d_cache.scala 24:26]
  reg  valid_0_59; // @[d_cache.scala 24:26]
  reg  valid_0_60; // @[d_cache.scala 24:26]
  reg  valid_0_61; // @[d_cache.scala 24:26]
  reg  valid_0_62; // @[d_cache.scala 24:26]
  reg  valid_0_63; // @[d_cache.scala 24:26]
  reg  valid_1_0; // @[d_cache.scala 25:26]
  reg  valid_1_1; // @[d_cache.scala 25:26]
  reg  valid_1_2; // @[d_cache.scala 25:26]
  reg  valid_1_3; // @[d_cache.scala 25:26]
  reg  valid_1_4; // @[d_cache.scala 25:26]
  reg  valid_1_5; // @[d_cache.scala 25:26]
  reg  valid_1_6; // @[d_cache.scala 25:26]
  reg  valid_1_7; // @[d_cache.scala 25:26]
  reg  valid_1_8; // @[d_cache.scala 25:26]
  reg  valid_1_9; // @[d_cache.scala 25:26]
  reg  valid_1_10; // @[d_cache.scala 25:26]
  reg  valid_1_11; // @[d_cache.scala 25:26]
  reg  valid_1_12; // @[d_cache.scala 25:26]
  reg  valid_1_13; // @[d_cache.scala 25:26]
  reg  valid_1_14; // @[d_cache.scala 25:26]
  reg  valid_1_15; // @[d_cache.scala 25:26]
  reg  valid_1_16; // @[d_cache.scala 25:26]
  reg  valid_1_17; // @[d_cache.scala 25:26]
  reg  valid_1_18; // @[d_cache.scala 25:26]
  reg  valid_1_19; // @[d_cache.scala 25:26]
  reg  valid_1_20; // @[d_cache.scala 25:26]
  reg  valid_1_21; // @[d_cache.scala 25:26]
  reg  valid_1_22; // @[d_cache.scala 25:26]
  reg  valid_1_23; // @[d_cache.scala 25:26]
  reg  valid_1_24; // @[d_cache.scala 25:26]
  reg  valid_1_25; // @[d_cache.scala 25:26]
  reg  valid_1_26; // @[d_cache.scala 25:26]
  reg  valid_1_27; // @[d_cache.scala 25:26]
  reg  valid_1_28; // @[d_cache.scala 25:26]
  reg  valid_1_29; // @[d_cache.scala 25:26]
  reg  valid_1_30; // @[d_cache.scala 25:26]
  reg  valid_1_31; // @[d_cache.scala 25:26]
  reg  valid_1_32; // @[d_cache.scala 25:26]
  reg  valid_1_33; // @[d_cache.scala 25:26]
  reg  valid_1_34; // @[d_cache.scala 25:26]
  reg  valid_1_35; // @[d_cache.scala 25:26]
  reg  valid_1_36; // @[d_cache.scala 25:26]
  reg  valid_1_37; // @[d_cache.scala 25:26]
  reg  valid_1_38; // @[d_cache.scala 25:26]
  reg  valid_1_39; // @[d_cache.scala 25:26]
  reg  valid_1_40; // @[d_cache.scala 25:26]
  reg  valid_1_41; // @[d_cache.scala 25:26]
  reg  valid_1_42; // @[d_cache.scala 25:26]
  reg  valid_1_43; // @[d_cache.scala 25:26]
  reg  valid_1_44; // @[d_cache.scala 25:26]
  reg  valid_1_45; // @[d_cache.scala 25:26]
  reg  valid_1_46; // @[d_cache.scala 25:26]
  reg  valid_1_47; // @[d_cache.scala 25:26]
  reg  valid_1_48; // @[d_cache.scala 25:26]
  reg  valid_1_49; // @[d_cache.scala 25:26]
  reg  valid_1_50; // @[d_cache.scala 25:26]
  reg  valid_1_51; // @[d_cache.scala 25:26]
  reg  valid_1_52; // @[d_cache.scala 25:26]
  reg  valid_1_53; // @[d_cache.scala 25:26]
  reg  valid_1_54; // @[d_cache.scala 25:26]
  reg  valid_1_55; // @[d_cache.scala 25:26]
  reg  valid_1_56; // @[d_cache.scala 25:26]
  reg  valid_1_57; // @[d_cache.scala 25:26]
  reg  valid_1_58; // @[d_cache.scala 25:26]
  reg  valid_1_59; // @[d_cache.scala 25:26]
  reg  valid_1_60; // @[d_cache.scala 25:26]
  reg  valid_1_61; // @[d_cache.scala 25:26]
  reg  valid_1_62; // @[d_cache.scala 25:26]
  reg  valid_1_63; // @[d_cache.scala 25:26]
  reg  dirty_0_0; // @[d_cache.scala 26:26]
  reg  dirty_0_1; // @[d_cache.scala 26:26]
  reg  dirty_0_2; // @[d_cache.scala 26:26]
  reg  dirty_0_3; // @[d_cache.scala 26:26]
  reg  dirty_0_4; // @[d_cache.scala 26:26]
  reg  dirty_0_5; // @[d_cache.scala 26:26]
  reg  dirty_0_6; // @[d_cache.scala 26:26]
  reg  dirty_0_7; // @[d_cache.scala 26:26]
  reg  dirty_0_8; // @[d_cache.scala 26:26]
  reg  dirty_0_9; // @[d_cache.scala 26:26]
  reg  dirty_0_10; // @[d_cache.scala 26:26]
  reg  dirty_0_11; // @[d_cache.scala 26:26]
  reg  dirty_0_12; // @[d_cache.scala 26:26]
  reg  dirty_0_13; // @[d_cache.scala 26:26]
  reg  dirty_0_14; // @[d_cache.scala 26:26]
  reg  dirty_0_15; // @[d_cache.scala 26:26]
  reg  dirty_0_16; // @[d_cache.scala 26:26]
  reg  dirty_0_17; // @[d_cache.scala 26:26]
  reg  dirty_0_18; // @[d_cache.scala 26:26]
  reg  dirty_0_19; // @[d_cache.scala 26:26]
  reg  dirty_0_20; // @[d_cache.scala 26:26]
  reg  dirty_0_21; // @[d_cache.scala 26:26]
  reg  dirty_0_22; // @[d_cache.scala 26:26]
  reg  dirty_0_23; // @[d_cache.scala 26:26]
  reg  dirty_0_24; // @[d_cache.scala 26:26]
  reg  dirty_0_25; // @[d_cache.scala 26:26]
  reg  dirty_0_26; // @[d_cache.scala 26:26]
  reg  dirty_0_27; // @[d_cache.scala 26:26]
  reg  dirty_0_28; // @[d_cache.scala 26:26]
  reg  dirty_0_29; // @[d_cache.scala 26:26]
  reg  dirty_0_30; // @[d_cache.scala 26:26]
  reg  dirty_0_31; // @[d_cache.scala 26:26]
  reg  dirty_0_32; // @[d_cache.scala 26:26]
  reg  dirty_0_33; // @[d_cache.scala 26:26]
  reg  dirty_0_34; // @[d_cache.scala 26:26]
  reg  dirty_0_35; // @[d_cache.scala 26:26]
  reg  dirty_0_36; // @[d_cache.scala 26:26]
  reg  dirty_0_37; // @[d_cache.scala 26:26]
  reg  dirty_0_38; // @[d_cache.scala 26:26]
  reg  dirty_0_39; // @[d_cache.scala 26:26]
  reg  dirty_0_40; // @[d_cache.scala 26:26]
  reg  dirty_0_41; // @[d_cache.scala 26:26]
  reg  dirty_0_42; // @[d_cache.scala 26:26]
  reg  dirty_0_43; // @[d_cache.scala 26:26]
  reg  dirty_0_44; // @[d_cache.scala 26:26]
  reg  dirty_0_45; // @[d_cache.scala 26:26]
  reg  dirty_0_46; // @[d_cache.scala 26:26]
  reg  dirty_0_47; // @[d_cache.scala 26:26]
  reg  dirty_0_48; // @[d_cache.scala 26:26]
  reg  dirty_0_49; // @[d_cache.scala 26:26]
  reg  dirty_0_50; // @[d_cache.scala 26:26]
  reg  dirty_0_51; // @[d_cache.scala 26:26]
  reg  dirty_0_52; // @[d_cache.scala 26:26]
  reg  dirty_0_53; // @[d_cache.scala 26:26]
  reg  dirty_0_54; // @[d_cache.scala 26:26]
  reg  dirty_0_55; // @[d_cache.scala 26:26]
  reg  dirty_0_56; // @[d_cache.scala 26:26]
  reg  dirty_0_57; // @[d_cache.scala 26:26]
  reg  dirty_0_58; // @[d_cache.scala 26:26]
  reg  dirty_0_59; // @[d_cache.scala 26:26]
  reg  dirty_0_60; // @[d_cache.scala 26:26]
  reg  dirty_0_61; // @[d_cache.scala 26:26]
  reg  dirty_0_62; // @[d_cache.scala 26:26]
  reg  dirty_0_63; // @[d_cache.scala 26:26]
  reg  dirty_1_0; // @[d_cache.scala 27:26]
  reg  dirty_1_1; // @[d_cache.scala 27:26]
  reg  dirty_1_2; // @[d_cache.scala 27:26]
  reg  dirty_1_3; // @[d_cache.scala 27:26]
  reg  dirty_1_4; // @[d_cache.scala 27:26]
  reg  dirty_1_5; // @[d_cache.scala 27:26]
  reg  dirty_1_6; // @[d_cache.scala 27:26]
  reg  dirty_1_7; // @[d_cache.scala 27:26]
  reg  dirty_1_8; // @[d_cache.scala 27:26]
  reg  dirty_1_9; // @[d_cache.scala 27:26]
  reg  dirty_1_10; // @[d_cache.scala 27:26]
  reg  dirty_1_11; // @[d_cache.scala 27:26]
  reg  dirty_1_12; // @[d_cache.scala 27:26]
  reg  dirty_1_13; // @[d_cache.scala 27:26]
  reg  dirty_1_14; // @[d_cache.scala 27:26]
  reg  dirty_1_15; // @[d_cache.scala 27:26]
  reg  dirty_1_16; // @[d_cache.scala 27:26]
  reg  dirty_1_17; // @[d_cache.scala 27:26]
  reg  dirty_1_18; // @[d_cache.scala 27:26]
  reg  dirty_1_19; // @[d_cache.scala 27:26]
  reg  dirty_1_20; // @[d_cache.scala 27:26]
  reg  dirty_1_21; // @[d_cache.scala 27:26]
  reg  dirty_1_22; // @[d_cache.scala 27:26]
  reg  dirty_1_23; // @[d_cache.scala 27:26]
  reg  dirty_1_24; // @[d_cache.scala 27:26]
  reg  dirty_1_25; // @[d_cache.scala 27:26]
  reg  dirty_1_26; // @[d_cache.scala 27:26]
  reg  dirty_1_27; // @[d_cache.scala 27:26]
  reg  dirty_1_28; // @[d_cache.scala 27:26]
  reg  dirty_1_29; // @[d_cache.scala 27:26]
  reg  dirty_1_30; // @[d_cache.scala 27:26]
  reg  dirty_1_31; // @[d_cache.scala 27:26]
  reg  dirty_1_32; // @[d_cache.scala 27:26]
  reg  dirty_1_33; // @[d_cache.scala 27:26]
  reg  dirty_1_34; // @[d_cache.scala 27:26]
  reg  dirty_1_35; // @[d_cache.scala 27:26]
  reg  dirty_1_36; // @[d_cache.scala 27:26]
  reg  dirty_1_37; // @[d_cache.scala 27:26]
  reg  dirty_1_38; // @[d_cache.scala 27:26]
  reg  dirty_1_39; // @[d_cache.scala 27:26]
  reg  dirty_1_40; // @[d_cache.scala 27:26]
  reg  dirty_1_41; // @[d_cache.scala 27:26]
  reg  dirty_1_42; // @[d_cache.scala 27:26]
  reg  dirty_1_43; // @[d_cache.scala 27:26]
  reg  dirty_1_44; // @[d_cache.scala 27:26]
  reg  dirty_1_45; // @[d_cache.scala 27:26]
  reg  dirty_1_46; // @[d_cache.scala 27:26]
  reg  dirty_1_47; // @[d_cache.scala 27:26]
  reg  dirty_1_48; // @[d_cache.scala 27:26]
  reg  dirty_1_49; // @[d_cache.scala 27:26]
  reg  dirty_1_50; // @[d_cache.scala 27:26]
  reg  dirty_1_51; // @[d_cache.scala 27:26]
  reg  dirty_1_52; // @[d_cache.scala 27:26]
  reg  dirty_1_53; // @[d_cache.scala 27:26]
  reg  dirty_1_54; // @[d_cache.scala 27:26]
  reg  dirty_1_55; // @[d_cache.scala 27:26]
  reg  dirty_1_56; // @[d_cache.scala 27:26]
  reg  dirty_1_57; // @[d_cache.scala 27:26]
  reg  dirty_1_58; // @[d_cache.scala 27:26]
  reg  dirty_1_59; // @[d_cache.scala 27:26]
  reg  dirty_1_60; // @[d_cache.scala 27:26]
  reg  dirty_1_61; // @[d_cache.scala 27:26]
  reg  dirty_1_62; // @[d_cache.scala 27:26]
  reg  dirty_1_63; // @[d_cache.scala 27:26]
  reg  way0_hit; // @[d_cache.scala 28:27]
  reg  way1_hit; // @[d_cache.scala 29:27]
  reg [63:0] write_back_data; // @[d_cache.scala 31:34]
  reg [31:0] write_back_addr; // @[d_cache.scala 32:34]
  reg [1:0] unuse_way; // @[d_cache.scala 35:28]
  reg [63:0] receive_data; // @[d_cache.scala 36:31]
  reg  quene; // @[d_cache.scala 37:24]
  wire [2:0] offset = io_from_lsu_araddr[2:0]; // @[d_cache.scala 39:36]
  wire [5:0] index = io_from_lsu_araddr[8:3]; // @[d_cache.scala 40:35]
  wire [22:0] tag = io_from_lsu_araddr[31:9]; // @[d_cache.scala 41:33]
  wire [5:0] _shift_bit_T_8 = offset == 3'h7 ? 6'h38 : 6'h0; // @[d_cache.scala 50:24]
  wire [5:0] _shift_bit_T_9 = offset == 3'h6 ? 6'h30 : _shift_bit_T_8; // @[d_cache.scala 49:24]
  wire [5:0] _shift_bit_T_10 = offset == 3'h5 ? 6'h28 : _shift_bit_T_9; // @[d_cache.scala 48:24]
  wire [5:0] _shift_bit_T_11 = offset == 3'h4 ? 6'h20 : _shift_bit_T_10; // @[d_cache.scala 47:24]
  wire [5:0] _shift_bit_T_12 = offset == 3'h3 ? 6'h18 : _shift_bit_T_11; // @[d_cache.scala 46:24]
  wire [5:0] _shift_bit_T_13 = offset == 3'h2 ? 6'h10 : _shift_bit_T_12; // @[d_cache.scala 45:24]
  wire [5:0] _shift_bit_T_14 = offset == 3'h1 ? 6'h8 : _shift_bit_T_13; // @[d_cache.scala 44:24]
  wire [5:0] shift_bit = offset == 3'h0 ? 6'h0 : _shift_bit_T_14; // @[d_cache.scala 43:24]
  wire [63:0] _wmask_T_4 = io_from_lsu_wstrb == 8'hff ? 64'hffffffffffffffff : 64'h0; // @[d_cache.scala 55:20]
  wire [63:0] _wmask_T_5 = io_from_lsu_wstrb == 8'hf ? 64'hffffffff : _wmask_T_4; // @[d_cache.scala 54:20]
  wire [63:0] _wmask_T_6 = io_from_lsu_wstrb == 8'h3 ? 64'hffff : _wmask_T_5; // @[d_cache.scala 53:20]
  wire [63:0] wmask = io_from_lsu_wstrb == 8'h1 ? 64'hff : _wmask_T_6; // @[d_cache.scala 52:20]
  wire [31:0] _GEN_1 = 6'h1 == index ? tag_0_1 : tag_0_0; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_2 = 6'h2 == index ? tag_0_2 : _GEN_1; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_3 = 6'h3 == index ? tag_0_3 : _GEN_2; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_4 = 6'h4 == index ? tag_0_4 : _GEN_3; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_5 = 6'h5 == index ? tag_0_5 : _GEN_4; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_6 = 6'h6 == index ? tag_0_6 : _GEN_5; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_7 = 6'h7 == index ? tag_0_7 : _GEN_6; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_8 = 6'h8 == index ? tag_0_8 : _GEN_7; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_9 = 6'h9 == index ? tag_0_9 : _GEN_8; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_10 = 6'ha == index ? tag_0_10 : _GEN_9; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_11 = 6'hb == index ? tag_0_11 : _GEN_10; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_12 = 6'hc == index ? tag_0_12 : _GEN_11; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_13 = 6'hd == index ? tag_0_13 : _GEN_12; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_14 = 6'he == index ? tag_0_14 : _GEN_13; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_15 = 6'hf == index ? tag_0_15 : _GEN_14; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_16 = 6'h10 == index ? tag_0_16 : _GEN_15; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_17 = 6'h11 == index ? tag_0_17 : _GEN_16; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_18 = 6'h12 == index ? tag_0_18 : _GEN_17; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_19 = 6'h13 == index ? tag_0_19 : _GEN_18; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_20 = 6'h14 == index ? tag_0_20 : _GEN_19; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_21 = 6'h15 == index ? tag_0_21 : _GEN_20; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_22 = 6'h16 == index ? tag_0_22 : _GEN_21; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_23 = 6'h17 == index ? tag_0_23 : _GEN_22; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_24 = 6'h18 == index ? tag_0_24 : _GEN_23; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_25 = 6'h19 == index ? tag_0_25 : _GEN_24; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_26 = 6'h1a == index ? tag_0_26 : _GEN_25; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_27 = 6'h1b == index ? tag_0_27 : _GEN_26; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_28 = 6'h1c == index ? tag_0_28 : _GEN_27; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_29 = 6'h1d == index ? tag_0_29 : _GEN_28; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_30 = 6'h1e == index ? tag_0_30 : _GEN_29; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_31 = 6'h1f == index ? tag_0_31 : _GEN_30; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_32 = 6'h20 == index ? tag_0_32 : _GEN_31; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_33 = 6'h21 == index ? tag_0_33 : _GEN_32; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_34 = 6'h22 == index ? tag_0_34 : _GEN_33; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_35 = 6'h23 == index ? tag_0_35 : _GEN_34; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_36 = 6'h24 == index ? tag_0_36 : _GEN_35; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_37 = 6'h25 == index ? tag_0_37 : _GEN_36; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_38 = 6'h26 == index ? tag_0_38 : _GEN_37; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_39 = 6'h27 == index ? tag_0_39 : _GEN_38; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_40 = 6'h28 == index ? tag_0_40 : _GEN_39; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_41 = 6'h29 == index ? tag_0_41 : _GEN_40; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_42 = 6'h2a == index ? tag_0_42 : _GEN_41; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_43 = 6'h2b == index ? tag_0_43 : _GEN_42; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_44 = 6'h2c == index ? tag_0_44 : _GEN_43; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_45 = 6'h2d == index ? tag_0_45 : _GEN_44; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_46 = 6'h2e == index ? tag_0_46 : _GEN_45; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_47 = 6'h2f == index ? tag_0_47 : _GEN_46; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_48 = 6'h30 == index ? tag_0_48 : _GEN_47; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_49 = 6'h31 == index ? tag_0_49 : _GEN_48; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_50 = 6'h32 == index ? tag_0_50 : _GEN_49; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_51 = 6'h33 == index ? tag_0_51 : _GEN_50; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_52 = 6'h34 == index ? tag_0_52 : _GEN_51; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_53 = 6'h35 == index ? tag_0_53 : _GEN_52; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_54 = 6'h36 == index ? tag_0_54 : _GEN_53; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_55 = 6'h37 == index ? tag_0_55 : _GEN_54; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_56 = 6'h38 == index ? tag_0_56 : _GEN_55; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_57 = 6'h39 == index ? tag_0_57 : _GEN_56; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_58 = 6'h3a == index ? tag_0_58 : _GEN_57; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_59 = 6'h3b == index ? tag_0_59 : _GEN_58; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_60 = 6'h3c == index ? tag_0_60 : _GEN_59; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_61 = 6'h3d == index ? tag_0_61 : _GEN_60; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_62 = 6'h3e == index ? tag_0_62 : _GEN_61; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_63 = 6'h3f == index ? tag_0_63 : _GEN_62; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_8027 = {{9'd0}, tag}; // @[d_cache.scala 57:24]
  wire  _GEN_65 = 6'h1 == index ? valid_0_1 : valid_0_0; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_66 = 6'h2 == index ? valid_0_2 : _GEN_65; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_67 = 6'h3 == index ? valid_0_3 : _GEN_66; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_68 = 6'h4 == index ? valid_0_4 : _GEN_67; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_69 = 6'h5 == index ? valid_0_5 : _GEN_68; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_70 = 6'h6 == index ? valid_0_6 : _GEN_69; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_71 = 6'h7 == index ? valid_0_7 : _GEN_70; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_72 = 6'h8 == index ? valid_0_8 : _GEN_71; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_73 = 6'h9 == index ? valid_0_9 : _GEN_72; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_74 = 6'ha == index ? valid_0_10 : _GEN_73; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_75 = 6'hb == index ? valid_0_11 : _GEN_74; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_76 = 6'hc == index ? valid_0_12 : _GEN_75; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_77 = 6'hd == index ? valid_0_13 : _GEN_76; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_78 = 6'he == index ? valid_0_14 : _GEN_77; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_79 = 6'hf == index ? valid_0_15 : _GEN_78; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_80 = 6'h10 == index ? valid_0_16 : _GEN_79; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_81 = 6'h11 == index ? valid_0_17 : _GEN_80; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_82 = 6'h12 == index ? valid_0_18 : _GEN_81; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_83 = 6'h13 == index ? valid_0_19 : _GEN_82; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_84 = 6'h14 == index ? valid_0_20 : _GEN_83; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_85 = 6'h15 == index ? valid_0_21 : _GEN_84; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_86 = 6'h16 == index ? valid_0_22 : _GEN_85; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_87 = 6'h17 == index ? valid_0_23 : _GEN_86; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_88 = 6'h18 == index ? valid_0_24 : _GEN_87; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_89 = 6'h19 == index ? valid_0_25 : _GEN_88; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_90 = 6'h1a == index ? valid_0_26 : _GEN_89; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_91 = 6'h1b == index ? valid_0_27 : _GEN_90; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_92 = 6'h1c == index ? valid_0_28 : _GEN_91; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_93 = 6'h1d == index ? valid_0_29 : _GEN_92; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_94 = 6'h1e == index ? valid_0_30 : _GEN_93; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_95 = 6'h1f == index ? valid_0_31 : _GEN_94; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_96 = 6'h20 == index ? valid_0_32 : _GEN_95; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_97 = 6'h21 == index ? valid_0_33 : _GEN_96; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_98 = 6'h22 == index ? valid_0_34 : _GEN_97; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_99 = 6'h23 == index ? valid_0_35 : _GEN_98; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_100 = 6'h24 == index ? valid_0_36 : _GEN_99; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_101 = 6'h25 == index ? valid_0_37 : _GEN_100; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_102 = 6'h26 == index ? valid_0_38 : _GEN_101; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_103 = 6'h27 == index ? valid_0_39 : _GEN_102; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_104 = 6'h28 == index ? valid_0_40 : _GEN_103; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_105 = 6'h29 == index ? valid_0_41 : _GEN_104; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_106 = 6'h2a == index ? valid_0_42 : _GEN_105; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_107 = 6'h2b == index ? valid_0_43 : _GEN_106; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_108 = 6'h2c == index ? valid_0_44 : _GEN_107; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_109 = 6'h2d == index ? valid_0_45 : _GEN_108; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_110 = 6'h2e == index ? valid_0_46 : _GEN_109; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_111 = 6'h2f == index ? valid_0_47 : _GEN_110; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_112 = 6'h30 == index ? valid_0_48 : _GEN_111; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_113 = 6'h31 == index ? valid_0_49 : _GEN_112; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_114 = 6'h32 == index ? valid_0_50 : _GEN_113; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_115 = 6'h33 == index ? valid_0_51 : _GEN_114; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_116 = 6'h34 == index ? valid_0_52 : _GEN_115; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_117 = 6'h35 == index ? valid_0_53 : _GEN_116; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_118 = 6'h36 == index ? valid_0_54 : _GEN_117; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_119 = 6'h37 == index ? valid_0_55 : _GEN_118; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_120 = 6'h38 == index ? valid_0_56 : _GEN_119; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_121 = 6'h39 == index ? valid_0_57 : _GEN_120; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_122 = 6'h3a == index ? valid_0_58 : _GEN_121; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_123 = 6'h3b == index ? valid_0_59 : _GEN_122; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_124 = 6'h3c == index ? valid_0_60 : _GEN_123; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_125 = 6'h3d == index ? valid_0_61 : _GEN_124; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_126 = 6'h3e == index ? valid_0_62 : _GEN_125; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_127 = 6'h3f == index ? valid_0_63 : _GEN_126; // @[d_cache.scala 57:{50,50}]
  wire  _T_4 = _GEN_63 == _GEN_8027 & _GEN_127; // @[d_cache.scala 57:33]
  wire [31:0] _GEN_130 = 6'h1 == index ? tag_1_1 : tag_1_0; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_131 = 6'h2 == index ? tag_1_2 : _GEN_130; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_132 = 6'h3 == index ? tag_1_3 : _GEN_131; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_133 = 6'h4 == index ? tag_1_4 : _GEN_132; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_134 = 6'h5 == index ? tag_1_5 : _GEN_133; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_135 = 6'h6 == index ? tag_1_6 : _GEN_134; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_136 = 6'h7 == index ? tag_1_7 : _GEN_135; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_137 = 6'h8 == index ? tag_1_8 : _GEN_136; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_138 = 6'h9 == index ? tag_1_9 : _GEN_137; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_139 = 6'ha == index ? tag_1_10 : _GEN_138; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_140 = 6'hb == index ? tag_1_11 : _GEN_139; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_141 = 6'hc == index ? tag_1_12 : _GEN_140; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_142 = 6'hd == index ? tag_1_13 : _GEN_141; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_143 = 6'he == index ? tag_1_14 : _GEN_142; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_144 = 6'hf == index ? tag_1_15 : _GEN_143; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_145 = 6'h10 == index ? tag_1_16 : _GEN_144; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_146 = 6'h11 == index ? tag_1_17 : _GEN_145; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_147 = 6'h12 == index ? tag_1_18 : _GEN_146; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_148 = 6'h13 == index ? tag_1_19 : _GEN_147; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_149 = 6'h14 == index ? tag_1_20 : _GEN_148; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_150 = 6'h15 == index ? tag_1_21 : _GEN_149; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_151 = 6'h16 == index ? tag_1_22 : _GEN_150; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_152 = 6'h17 == index ? tag_1_23 : _GEN_151; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_153 = 6'h18 == index ? tag_1_24 : _GEN_152; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_154 = 6'h19 == index ? tag_1_25 : _GEN_153; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_155 = 6'h1a == index ? tag_1_26 : _GEN_154; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_156 = 6'h1b == index ? tag_1_27 : _GEN_155; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_157 = 6'h1c == index ? tag_1_28 : _GEN_156; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_158 = 6'h1d == index ? tag_1_29 : _GEN_157; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_159 = 6'h1e == index ? tag_1_30 : _GEN_158; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_160 = 6'h1f == index ? tag_1_31 : _GEN_159; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_161 = 6'h20 == index ? tag_1_32 : _GEN_160; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_162 = 6'h21 == index ? tag_1_33 : _GEN_161; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_163 = 6'h22 == index ? tag_1_34 : _GEN_162; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_164 = 6'h23 == index ? tag_1_35 : _GEN_163; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_165 = 6'h24 == index ? tag_1_36 : _GEN_164; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_166 = 6'h25 == index ? tag_1_37 : _GEN_165; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_167 = 6'h26 == index ? tag_1_38 : _GEN_166; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_168 = 6'h27 == index ? tag_1_39 : _GEN_167; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_169 = 6'h28 == index ? tag_1_40 : _GEN_168; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_170 = 6'h29 == index ? tag_1_41 : _GEN_169; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_171 = 6'h2a == index ? tag_1_42 : _GEN_170; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_172 = 6'h2b == index ? tag_1_43 : _GEN_171; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_173 = 6'h2c == index ? tag_1_44 : _GEN_172; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_174 = 6'h2d == index ? tag_1_45 : _GEN_173; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_175 = 6'h2e == index ? tag_1_46 : _GEN_174; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_176 = 6'h2f == index ? tag_1_47 : _GEN_175; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_177 = 6'h30 == index ? tag_1_48 : _GEN_176; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_178 = 6'h31 == index ? tag_1_49 : _GEN_177; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_179 = 6'h32 == index ? tag_1_50 : _GEN_178; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_180 = 6'h33 == index ? tag_1_51 : _GEN_179; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_181 = 6'h34 == index ? tag_1_52 : _GEN_180; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_182 = 6'h35 == index ? tag_1_53 : _GEN_181; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_183 = 6'h36 == index ? tag_1_54 : _GEN_182; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_184 = 6'h37 == index ? tag_1_55 : _GEN_183; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_185 = 6'h38 == index ? tag_1_56 : _GEN_184; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_186 = 6'h39 == index ? tag_1_57 : _GEN_185; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_187 = 6'h3a == index ? tag_1_58 : _GEN_186; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_188 = 6'h3b == index ? tag_1_59 : _GEN_187; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_189 = 6'h3c == index ? tag_1_60 : _GEN_188; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_190 = 6'h3d == index ? tag_1_61 : _GEN_189; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_191 = 6'h3e == index ? tag_1_62 : _GEN_190; // @[d_cache.scala 62:{24,24}]
  wire [31:0] _GEN_192 = 6'h3f == index ? tag_1_63 : _GEN_191; // @[d_cache.scala 62:{24,24}]
  wire  _GEN_194 = 6'h1 == index ? valid_1_1 : valid_1_0; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_195 = 6'h2 == index ? valid_1_2 : _GEN_194; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_196 = 6'h3 == index ? valid_1_3 : _GEN_195; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_197 = 6'h4 == index ? valid_1_4 : _GEN_196; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_198 = 6'h5 == index ? valid_1_5 : _GEN_197; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_199 = 6'h6 == index ? valid_1_6 : _GEN_198; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_200 = 6'h7 == index ? valid_1_7 : _GEN_199; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_201 = 6'h8 == index ? valid_1_8 : _GEN_200; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_202 = 6'h9 == index ? valid_1_9 : _GEN_201; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_203 = 6'ha == index ? valid_1_10 : _GEN_202; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_204 = 6'hb == index ? valid_1_11 : _GEN_203; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_205 = 6'hc == index ? valid_1_12 : _GEN_204; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_206 = 6'hd == index ? valid_1_13 : _GEN_205; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_207 = 6'he == index ? valid_1_14 : _GEN_206; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_208 = 6'hf == index ? valid_1_15 : _GEN_207; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_209 = 6'h10 == index ? valid_1_16 : _GEN_208; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_210 = 6'h11 == index ? valid_1_17 : _GEN_209; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_211 = 6'h12 == index ? valid_1_18 : _GEN_210; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_212 = 6'h13 == index ? valid_1_19 : _GEN_211; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_213 = 6'h14 == index ? valid_1_20 : _GEN_212; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_214 = 6'h15 == index ? valid_1_21 : _GEN_213; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_215 = 6'h16 == index ? valid_1_22 : _GEN_214; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_216 = 6'h17 == index ? valid_1_23 : _GEN_215; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_217 = 6'h18 == index ? valid_1_24 : _GEN_216; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_218 = 6'h19 == index ? valid_1_25 : _GEN_217; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_219 = 6'h1a == index ? valid_1_26 : _GEN_218; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_220 = 6'h1b == index ? valid_1_27 : _GEN_219; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_221 = 6'h1c == index ? valid_1_28 : _GEN_220; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_222 = 6'h1d == index ? valid_1_29 : _GEN_221; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_223 = 6'h1e == index ? valid_1_30 : _GEN_222; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_224 = 6'h1f == index ? valid_1_31 : _GEN_223; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_225 = 6'h20 == index ? valid_1_32 : _GEN_224; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_226 = 6'h21 == index ? valid_1_33 : _GEN_225; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_227 = 6'h22 == index ? valid_1_34 : _GEN_226; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_228 = 6'h23 == index ? valid_1_35 : _GEN_227; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_229 = 6'h24 == index ? valid_1_36 : _GEN_228; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_230 = 6'h25 == index ? valid_1_37 : _GEN_229; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_231 = 6'h26 == index ? valid_1_38 : _GEN_230; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_232 = 6'h27 == index ? valid_1_39 : _GEN_231; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_233 = 6'h28 == index ? valid_1_40 : _GEN_232; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_234 = 6'h29 == index ? valid_1_41 : _GEN_233; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_235 = 6'h2a == index ? valid_1_42 : _GEN_234; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_236 = 6'h2b == index ? valid_1_43 : _GEN_235; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_237 = 6'h2c == index ? valid_1_44 : _GEN_236; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_238 = 6'h2d == index ? valid_1_45 : _GEN_237; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_239 = 6'h2e == index ? valid_1_46 : _GEN_238; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_240 = 6'h2f == index ? valid_1_47 : _GEN_239; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_241 = 6'h30 == index ? valid_1_48 : _GEN_240; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_242 = 6'h31 == index ? valid_1_49 : _GEN_241; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_243 = 6'h32 == index ? valid_1_50 : _GEN_242; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_244 = 6'h33 == index ? valid_1_51 : _GEN_243; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_245 = 6'h34 == index ? valid_1_52 : _GEN_244; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_246 = 6'h35 == index ? valid_1_53 : _GEN_245; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_247 = 6'h36 == index ? valid_1_54 : _GEN_246; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_248 = 6'h37 == index ? valid_1_55 : _GEN_247; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_249 = 6'h38 == index ? valid_1_56 : _GEN_248; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_250 = 6'h39 == index ? valid_1_57 : _GEN_249; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_251 = 6'h3a == index ? valid_1_58 : _GEN_250; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_252 = 6'h3b == index ? valid_1_59 : _GEN_251; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_253 = 6'h3c == index ? valid_1_60 : _GEN_252; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_254 = 6'h3d == index ? valid_1_61 : _GEN_253; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_255 = 6'h3e == index ? valid_1_62 : _GEN_254; // @[d_cache.scala 62:{50,50}]
  wire  _GEN_256 = 6'h3f == index ? valid_1_63 : _GEN_255; // @[d_cache.scala 62:{50,50}]
  wire  _T_7 = _GEN_192 == _GEN_8027 & _GEN_256; // @[d_cache.scala 62:33]
  reg [2:0] state; // @[d_cache.scala 76:24]
  wire  _T_14 = 3'h0 == state; // @[d_cache.scala 81:18]
  wire  _T_15 = 3'h1 == state; // @[d_cache.scala 81:18]
  wire  _GEN_263 = 6'h1 == index ? dirty_0_1 : dirty_0_0; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_264 = 6'h2 == index ? dirty_0_2 : _GEN_263; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_265 = 6'h3 == index ? dirty_0_3 : _GEN_264; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_266 = 6'h4 == index ? dirty_0_4 : _GEN_265; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_267 = 6'h5 == index ? dirty_0_5 : _GEN_266; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_268 = 6'h6 == index ? dirty_0_6 : _GEN_267; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_269 = 6'h7 == index ? dirty_0_7 : _GEN_268; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_270 = 6'h8 == index ? dirty_0_8 : _GEN_269; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_271 = 6'h9 == index ? dirty_0_9 : _GEN_270; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_272 = 6'ha == index ? dirty_0_10 : _GEN_271; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_273 = 6'hb == index ? dirty_0_11 : _GEN_272; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_274 = 6'hc == index ? dirty_0_12 : _GEN_273; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_275 = 6'hd == index ? dirty_0_13 : _GEN_274; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_276 = 6'he == index ? dirty_0_14 : _GEN_275; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_277 = 6'hf == index ? dirty_0_15 : _GEN_276; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_278 = 6'h10 == index ? dirty_0_16 : _GEN_277; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_279 = 6'h11 == index ? dirty_0_17 : _GEN_278; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_280 = 6'h12 == index ? dirty_0_18 : _GEN_279; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_281 = 6'h13 == index ? dirty_0_19 : _GEN_280; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_282 = 6'h14 == index ? dirty_0_20 : _GEN_281; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_283 = 6'h15 == index ? dirty_0_21 : _GEN_282; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_284 = 6'h16 == index ? dirty_0_22 : _GEN_283; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_285 = 6'h17 == index ? dirty_0_23 : _GEN_284; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_286 = 6'h18 == index ? dirty_0_24 : _GEN_285; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_287 = 6'h19 == index ? dirty_0_25 : _GEN_286; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_288 = 6'h1a == index ? dirty_0_26 : _GEN_287; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_289 = 6'h1b == index ? dirty_0_27 : _GEN_288; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_290 = 6'h1c == index ? dirty_0_28 : _GEN_289; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_291 = 6'h1d == index ? dirty_0_29 : _GEN_290; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_292 = 6'h1e == index ? dirty_0_30 : _GEN_291; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_293 = 6'h1f == index ? dirty_0_31 : _GEN_292; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_294 = 6'h20 == index ? dirty_0_32 : _GEN_293; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_295 = 6'h21 == index ? dirty_0_33 : _GEN_294; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_296 = 6'h22 == index ? dirty_0_34 : _GEN_295; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_297 = 6'h23 == index ? dirty_0_35 : _GEN_296; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_298 = 6'h24 == index ? dirty_0_36 : _GEN_297; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_299 = 6'h25 == index ? dirty_0_37 : _GEN_298; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_300 = 6'h26 == index ? dirty_0_38 : _GEN_299; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_301 = 6'h27 == index ? dirty_0_39 : _GEN_300; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_302 = 6'h28 == index ? dirty_0_40 : _GEN_301; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_303 = 6'h29 == index ? dirty_0_41 : _GEN_302; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_304 = 6'h2a == index ? dirty_0_42 : _GEN_303; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_305 = 6'h2b == index ? dirty_0_43 : _GEN_304; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_306 = 6'h2c == index ? dirty_0_44 : _GEN_305; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_307 = 6'h2d == index ? dirty_0_45 : _GEN_306; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_308 = 6'h2e == index ? dirty_0_46 : _GEN_307; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_309 = 6'h2f == index ? dirty_0_47 : _GEN_308; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_310 = 6'h30 == index ? dirty_0_48 : _GEN_309; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_311 = 6'h31 == index ? dirty_0_49 : _GEN_310; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_312 = 6'h32 == index ? dirty_0_50 : _GEN_311; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_313 = 6'h33 == index ? dirty_0_51 : _GEN_312; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_314 = 6'h34 == index ? dirty_0_52 : _GEN_313; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_315 = 6'h35 == index ? dirty_0_53 : _GEN_314; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_316 = 6'h36 == index ? dirty_0_54 : _GEN_315; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_317 = 6'h37 == index ? dirty_0_55 : _GEN_316; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_318 = 6'h38 == index ? dirty_0_56 : _GEN_317; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_319 = 6'h39 == index ? dirty_0_57 : _GEN_318; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_320 = 6'h3a == index ? dirty_0_58 : _GEN_319; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_321 = 6'h3b == index ? dirty_0_59 : _GEN_320; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_322 = 6'h3c == index ? dirty_0_60 : _GEN_321; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_323 = 6'h3d == index ? dirty_0_61 : _GEN_322; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_324 = 6'h3e == index ? dirty_0_62 : _GEN_323; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_325 = 6'h3f == index ? dirty_0_63 : _GEN_324; // @[d_cache.scala 93:{27,27}]
  wire [2:0] _GEN_326 = io_from_lsu_rready ? 3'h0 : state; // @[d_cache.scala 76:24 92:41 94:27]
  wire  _GEN_328 = 6'h1 == index ? dirty_1_1 : dirty_1_0; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_329 = 6'h2 == index ? dirty_1_2 : _GEN_328; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_330 = 6'h3 == index ? dirty_1_3 : _GEN_329; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_331 = 6'h4 == index ? dirty_1_4 : _GEN_330; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_332 = 6'h5 == index ? dirty_1_5 : _GEN_331; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_333 = 6'h6 == index ? dirty_1_6 : _GEN_332; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_334 = 6'h7 == index ? dirty_1_7 : _GEN_333; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_335 = 6'h8 == index ? dirty_1_8 : _GEN_334; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_336 = 6'h9 == index ? dirty_1_9 : _GEN_335; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_337 = 6'ha == index ? dirty_1_10 : _GEN_336; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_338 = 6'hb == index ? dirty_1_11 : _GEN_337; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_339 = 6'hc == index ? dirty_1_12 : _GEN_338; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_340 = 6'hd == index ? dirty_1_13 : _GEN_339; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_341 = 6'he == index ? dirty_1_14 : _GEN_340; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_342 = 6'hf == index ? dirty_1_15 : _GEN_341; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_343 = 6'h10 == index ? dirty_1_16 : _GEN_342; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_344 = 6'h11 == index ? dirty_1_17 : _GEN_343; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_345 = 6'h12 == index ? dirty_1_18 : _GEN_344; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_346 = 6'h13 == index ? dirty_1_19 : _GEN_345; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_347 = 6'h14 == index ? dirty_1_20 : _GEN_346; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_348 = 6'h15 == index ? dirty_1_21 : _GEN_347; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_349 = 6'h16 == index ? dirty_1_22 : _GEN_348; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_350 = 6'h17 == index ? dirty_1_23 : _GEN_349; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_351 = 6'h18 == index ? dirty_1_24 : _GEN_350; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_352 = 6'h19 == index ? dirty_1_25 : _GEN_351; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_353 = 6'h1a == index ? dirty_1_26 : _GEN_352; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_354 = 6'h1b == index ? dirty_1_27 : _GEN_353; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_355 = 6'h1c == index ? dirty_1_28 : _GEN_354; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_356 = 6'h1d == index ? dirty_1_29 : _GEN_355; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_357 = 6'h1e == index ? dirty_1_30 : _GEN_356; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_358 = 6'h1f == index ? dirty_1_31 : _GEN_357; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_359 = 6'h20 == index ? dirty_1_32 : _GEN_358; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_360 = 6'h21 == index ? dirty_1_33 : _GEN_359; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_361 = 6'h22 == index ? dirty_1_34 : _GEN_360; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_362 = 6'h23 == index ? dirty_1_35 : _GEN_361; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_363 = 6'h24 == index ? dirty_1_36 : _GEN_362; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_364 = 6'h25 == index ? dirty_1_37 : _GEN_363; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_365 = 6'h26 == index ? dirty_1_38 : _GEN_364; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_366 = 6'h27 == index ? dirty_1_39 : _GEN_365; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_367 = 6'h28 == index ? dirty_1_40 : _GEN_366; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_368 = 6'h29 == index ? dirty_1_41 : _GEN_367; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_369 = 6'h2a == index ? dirty_1_42 : _GEN_368; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_370 = 6'h2b == index ? dirty_1_43 : _GEN_369; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_371 = 6'h2c == index ? dirty_1_44 : _GEN_370; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_372 = 6'h2d == index ? dirty_1_45 : _GEN_371; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_373 = 6'h2e == index ? dirty_1_46 : _GEN_372; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_374 = 6'h2f == index ? dirty_1_47 : _GEN_373; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_375 = 6'h30 == index ? dirty_1_48 : _GEN_374; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_376 = 6'h31 == index ? dirty_1_49 : _GEN_375; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_377 = 6'h32 == index ? dirty_1_50 : _GEN_376; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_378 = 6'h33 == index ? dirty_1_51 : _GEN_377; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_379 = 6'h34 == index ? dirty_1_52 : _GEN_378; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_380 = 6'h35 == index ? dirty_1_53 : _GEN_379; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_381 = 6'h36 == index ? dirty_1_54 : _GEN_380; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_382 = 6'h37 == index ? dirty_1_55 : _GEN_381; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_383 = 6'h38 == index ? dirty_1_56 : _GEN_382; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_384 = 6'h39 == index ? dirty_1_57 : _GEN_383; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_385 = 6'h3a == index ? dirty_1_58 : _GEN_384; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_386 = 6'h3b == index ? dirty_1_59 : _GEN_385; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_387 = 6'h3c == index ? dirty_1_60 : _GEN_386; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_388 = 6'h3d == index ? dirty_1_61 : _GEN_387; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_389 = 6'h3e == index ? dirty_1_62 : _GEN_388; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_390 = 6'h3f == index ? dirty_1_63 : _GEN_389; // @[d_cache.scala 99:{27,27}]
  wire [2:0] _GEN_391 = way1_hit ? _GEN_326 : 3'h3; // @[d_cache.scala 103:23 97:33]
  wire [63:0] _GEN_8029 = {{32'd0}, io_from_lsu_wdata}; // @[d_cache.scala 109:53]
  wire [63:0] _ram_0_T = _GEN_8029 & wmask; // @[d_cache.scala 109:53]
  wire [126:0] _GEN_8685 = {{63'd0}, _ram_0_T}; // @[d_cache.scala 109:62]
  wire [126:0] _ram_0_T_1 = _GEN_8685 << shift_bit; // @[d_cache.scala 109:62]
  wire [126:0] _GEN_8686 = {{63'd0}, wmask}; // @[d_cache.scala 109:102]
  wire [126:0] _ram_0_T_2 = _GEN_8686 << shift_bit; // @[d_cache.scala 109:102]
  wire [126:0] _ram_0_T_3 = ~_ram_0_T_2; // @[d_cache.scala 109:94]
  wire [63:0] _GEN_394 = 6'h1 == index ? ram_0_1 : ram_0_0; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_395 = 6'h2 == index ? ram_0_2 : _GEN_394; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_396 = 6'h3 == index ? ram_0_3 : _GEN_395; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_397 = 6'h4 == index ? ram_0_4 : _GEN_396; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_398 = 6'h5 == index ? ram_0_5 : _GEN_397; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_399 = 6'h6 == index ? ram_0_6 : _GEN_398; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_400 = 6'h7 == index ? ram_0_7 : _GEN_399; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_401 = 6'h8 == index ? ram_0_8 : _GEN_400; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_402 = 6'h9 == index ? ram_0_9 : _GEN_401; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_403 = 6'ha == index ? ram_0_10 : _GEN_402; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_404 = 6'hb == index ? ram_0_11 : _GEN_403; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_405 = 6'hc == index ? ram_0_12 : _GEN_404; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_406 = 6'hd == index ? ram_0_13 : _GEN_405; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_407 = 6'he == index ? ram_0_14 : _GEN_406; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_408 = 6'hf == index ? ram_0_15 : _GEN_407; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_409 = 6'h10 == index ? ram_0_16 : _GEN_408; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_410 = 6'h11 == index ? ram_0_17 : _GEN_409; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_411 = 6'h12 == index ? ram_0_18 : _GEN_410; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_412 = 6'h13 == index ? ram_0_19 : _GEN_411; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_413 = 6'h14 == index ? ram_0_20 : _GEN_412; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_414 = 6'h15 == index ? ram_0_21 : _GEN_413; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_415 = 6'h16 == index ? ram_0_22 : _GEN_414; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_416 = 6'h17 == index ? ram_0_23 : _GEN_415; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_417 = 6'h18 == index ? ram_0_24 : _GEN_416; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_418 = 6'h19 == index ? ram_0_25 : _GEN_417; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_419 = 6'h1a == index ? ram_0_26 : _GEN_418; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_420 = 6'h1b == index ? ram_0_27 : _GEN_419; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_421 = 6'h1c == index ? ram_0_28 : _GEN_420; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_422 = 6'h1d == index ? ram_0_29 : _GEN_421; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_423 = 6'h1e == index ? ram_0_30 : _GEN_422; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_424 = 6'h1f == index ? ram_0_31 : _GEN_423; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_425 = 6'h20 == index ? ram_0_32 : _GEN_424; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_426 = 6'h21 == index ? ram_0_33 : _GEN_425; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_427 = 6'h22 == index ? ram_0_34 : _GEN_426; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_428 = 6'h23 == index ? ram_0_35 : _GEN_427; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_429 = 6'h24 == index ? ram_0_36 : _GEN_428; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_430 = 6'h25 == index ? ram_0_37 : _GEN_429; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_431 = 6'h26 == index ? ram_0_38 : _GEN_430; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_432 = 6'h27 == index ? ram_0_39 : _GEN_431; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_433 = 6'h28 == index ? ram_0_40 : _GEN_432; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_434 = 6'h29 == index ? ram_0_41 : _GEN_433; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_435 = 6'h2a == index ? ram_0_42 : _GEN_434; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_436 = 6'h2b == index ? ram_0_43 : _GEN_435; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_437 = 6'h2c == index ? ram_0_44 : _GEN_436; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_438 = 6'h2d == index ? ram_0_45 : _GEN_437; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_439 = 6'h2e == index ? ram_0_46 : _GEN_438; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_440 = 6'h2f == index ? ram_0_47 : _GEN_439; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_441 = 6'h30 == index ? ram_0_48 : _GEN_440; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_442 = 6'h31 == index ? ram_0_49 : _GEN_441; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_443 = 6'h32 == index ? ram_0_50 : _GEN_442; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_444 = 6'h33 == index ? ram_0_51 : _GEN_443; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_445 = 6'h34 == index ? ram_0_52 : _GEN_444; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_446 = 6'h35 == index ? ram_0_53 : _GEN_445; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_447 = 6'h36 == index ? ram_0_54 : _GEN_446; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_448 = 6'h37 == index ? ram_0_55 : _GEN_447; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_449 = 6'h38 == index ? ram_0_56 : _GEN_448; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_450 = 6'h39 == index ? ram_0_57 : _GEN_449; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_451 = 6'h3a == index ? ram_0_58 : _GEN_450; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_452 = 6'h3b == index ? ram_0_59 : _GEN_451; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_453 = 6'h3c == index ? ram_0_60 : _GEN_452; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_454 = 6'h3d == index ? ram_0_61 : _GEN_453; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_455 = 6'h3e == index ? ram_0_62 : _GEN_454; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_456 = 6'h3f == index ? ram_0_63 : _GEN_455; // @[d_cache.scala 109:{92,92}]
  wire [126:0] _GEN_8030 = {{63'd0}, _GEN_456}; // @[d_cache.scala 109:92]
  wire [126:0] _ram_0_T_4 = _GEN_8030 & _ram_0_T_3; // @[d_cache.scala 109:92]
  wire [126:0] _ram_0_T_5 = _ram_0_T_1 | _ram_0_T_4; // @[d_cache.scala 109:76]
  wire [63:0] _GEN_457 = 6'h0 == index ? _ram_0_T_5[63:0] : ram_0_0; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_458 = 6'h1 == index ? _ram_0_T_5[63:0] : ram_0_1; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_459 = 6'h2 == index ? _ram_0_T_5[63:0] : ram_0_2; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_460 = 6'h3 == index ? _ram_0_T_5[63:0] : ram_0_3; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_461 = 6'h4 == index ? _ram_0_T_5[63:0] : ram_0_4; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_462 = 6'h5 == index ? _ram_0_T_5[63:0] : ram_0_5; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_463 = 6'h6 == index ? _ram_0_T_5[63:0] : ram_0_6; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_464 = 6'h7 == index ? _ram_0_T_5[63:0] : ram_0_7; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_465 = 6'h8 == index ? _ram_0_T_5[63:0] : ram_0_8; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_466 = 6'h9 == index ? _ram_0_T_5[63:0] : ram_0_9; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_467 = 6'ha == index ? _ram_0_T_5[63:0] : ram_0_10; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_468 = 6'hb == index ? _ram_0_T_5[63:0] : ram_0_11; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_469 = 6'hc == index ? _ram_0_T_5[63:0] : ram_0_12; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_470 = 6'hd == index ? _ram_0_T_5[63:0] : ram_0_13; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_471 = 6'he == index ? _ram_0_T_5[63:0] : ram_0_14; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_472 = 6'hf == index ? _ram_0_T_5[63:0] : ram_0_15; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_473 = 6'h10 == index ? _ram_0_T_5[63:0] : ram_0_16; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_474 = 6'h11 == index ? _ram_0_T_5[63:0] : ram_0_17; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_475 = 6'h12 == index ? _ram_0_T_5[63:0] : ram_0_18; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_476 = 6'h13 == index ? _ram_0_T_5[63:0] : ram_0_19; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_477 = 6'h14 == index ? _ram_0_T_5[63:0] : ram_0_20; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_478 = 6'h15 == index ? _ram_0_T_5[63:0] : ram_0_21; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_479 = 6'h16 == index ? _ram_0_T_5[63:0] : ram_0_22; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_480 = 6'h17 == index ? _ram_0_T_5[63:0] : ram_0_23; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_481 = 6'h18 == index ? _ram_0_T_5[63:0] : ram_0_24; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_482 = 6'h19 == index ? _ram_0_T_5[63:0] : ram_0_25; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_483 = 6'h1a == index ? _ram_0_T_5[63:0] : ram_0_26; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_484 = 6'h1b == index ? _ram_0_T_5[63:0] : ram_0_27; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_485 = 6'h1c == index ? _ram_0_T_5[63:0] : ram_0_28; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_486 = 6'h1d == index ? _ram_0_T_5[63:0] : ram_0_29; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_487 = 6'h1e == index ? _ram_0_T_5[63:0] : ram_0_30; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_488 = 6'h1f == index ? _ram_0_T_5[63:0] : ram_0_31; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_489 = 6'h20 == index ? _ram_0_T_5[63:0] : ram_0_32; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_490 = 6'h21 == index ? _ram_0_T_5[63:0] : ram_0_33; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_491 = 6'h22 == index ? _ram_0_T_5[63:0] : ram_0_34; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_492 = 6'h23 == index ? _ram_0_T_5[63:0] : ram_0_35; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_493 = 6'h24 == index ? _ram_0_T_5[63:0] : ram_0_36; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_494 = 6'h25 == index ? _ram_0_T_5[63:0] : ram_0_37; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_495 = 6'h26 == index ? _ram_0_T_5[63:0] : ram_0_38; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_496 = 6'h27 == index ? _ram_0_T_5[63:0] : ram_0_39; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_497 = 6'h28 == index ? _ram_0_T_5[63:0] : ram_0_40; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_498 = 6'h29 == index ? _ram_0_T_5[63:0] : ram_0_41; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_499 = 6'h2a == index ? _ram_0_T_5[63:0] : ram_0_42; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_500 = 6'h2b == index ? _ram_0_T_5[63:0] : ram_0_43; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_501 = 6'h2c == index ? _ram_0_T_5[63:0] : ram_0_44; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_502 = 6'h2d == index ? _ram_0_T_5[63:0] : ram_0_45; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_503 = 6'h2e == index ? _ram_0_T_5[63:0] : ram_0_46; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_504 = 6'h2f == index ? _ram_0_T_5[63:0] : ram_0_47; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_505 = 6'h30 == index ? _ram_0_T_5[63:0] : ram_0_48; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_506 = 6'h31 == index ? _ram_0_T_5[63:0] : ram_0_49; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_507 = 6'h32 == index ? _ram_0_T_5[63:0] : ram_0_50; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_508 = 6'h33 == index ? _ram_0_T_5[63:0] : ram_0_51; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_509 = 6'h34 == index ? _ram_0_T_5[63:0] : ram_0_52; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_510 = 6'h35 == index ? _ram_0_T_5[63:0] : ram_0_53; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_511 = 6'h36 == index ? _ram_0_T_5[63:0] : ram_0_54; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_512 = 6'h37 == index ? _ram_0_T_5[63:0] : ram_0_55; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_513 = 6'h38 == index ? _ram_0_T_5[63:0] : ram_0_56; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_514 = 6'h39 == index ? _ram_0_T_5[63:0] : ram_0_57; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_515 = 6'h3a == index ? _ram_0_T_5[63:0] : ram_0_58; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_516 = 6'h3b == index ? _ram_0_T_5[63:0] : ram_0_59; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_517 = 6'h3c == index ? _ram_0_T_5[63:0] : ram_0_60; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_518 = 6'h3d == index ? _ram_0_T_5[63:0] : ram_0_61; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_519 = 6'h3e == index ? _ram_0_T_5[63:0] : ram_0_62; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_520 = 6'h3f == index ? _ram_0_T_5[63:0] : ram_0_63; // @[d_cache.scala 109:{30,30} 18:24]
  wire  _GEN_8031 = 6'h0 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_521 = 6'h0 == index | valid_0_0; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8032 = 6'h1 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_522 = 6'h1 == index | valid_0_1; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8033 = 6'h2 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_523 = 6'h2 == index | valid_0_2; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8034 = 6'h3 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_524 = 6'h3 == index | valid_0_3; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8035 = 6'h4 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_525 = 6'h4 == index | valid_0_4; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8036 = 6'h5 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_526 = 6'h5 == index | valid_0_5; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8037 = 6'h6 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_527 = 6'h6 == index | valid_0_6; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8038 = 6'h7 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_528 = 6'h7 == index | valid_0_7; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8039 = 6'h8 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_529 = 6'h8 == index | valid_0_8; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8040 = 6'h9 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_530 = 6'h9 == index | valid_0_9; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8041 = 6'ha == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_531 = 6'ha == index | valid_0_10; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8042 = 6'hb == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_532 = 6'hb == index | valid_0_11; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8043 = 6'hc == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_533 = 6'hc == index | valid_0_12; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8044 = 6'hd == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_534 = 6'hd == index | valid_0_13; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8045 = 6'he == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_535 = 6'he == index | valid_0_14; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8046 = 6'hf == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_536 = 6'hf == index | valid_0_15; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8047 = 6'h10 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_537 = 6'h10 == index | valid_0_16; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8048 = 6'h11 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_538 = 6'h11 == index | valid_0_17; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8049 = 6'h12 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_539 = 6'h12 == index | valid_0_18; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8050 = 6'h13 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_540 = 6'h13 == index | valid_0_19; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8051 = 6'h14 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_541 = 6'h14 == index | valid_0_20; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8052 = 6'h15 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_542 = 6'h15 == index | valid_0_21; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8053 = 6'h16 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_543 = 6'h16 == index | valid_0_22; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8054 = 6'h17 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_544 = 6'h17 == index | valid_0_23; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8055 = 6'h18 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_545 = 6'h18 == index | valid_0_24; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8056 = 6'h19 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_546 = 6'h19 == index | valid_0_25; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8057 = 6'h1a == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_547 = 6'h1a == index | valid_0_26; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8058 = 6'h1b == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_548 = 6'h1b == index | valid_0_27; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8059 = 6'h1c == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_549 = 6'h1c == index | valid_0_28; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8060 = 6'h1d == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_550 = 6'h1d == index | valid_0_29; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8061 = 6'h1e == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_551 = 6'h1e == index | valid_0_30; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8062 = 6'h1f == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_552 = 6'h1f == index | valid_0_31; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8063 = 6'h20 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_553 = 6'h20 == index | valid_0_32; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8064 = 6'h21 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_554 = 6'h21 == index | valid_0_33; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8065 = 6'h22 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_555 = 6'h22 == index | valid_0_34; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8066 = 6'h23 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_556 = 6'h23 == index | valid_0_35; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8067 = 6'h24 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_557 = 6'h24 == index | valid_0_36; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8068 = 6'h25 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_558 = 6'h25 == index | valid_0_37; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8069 = 6'h26 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_559 = 6'h26 == index | valid_0_38; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8070 = 6'h27 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_560 = 6'h27 == index | valid_0_39; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8071 = 6'h28 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_561 = 6'h28 == index | valid_0_40; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8072 = 6'h29 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_562 = 6'h29 == index | valid_0_41; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8073 = 6'h2a == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_563 = 6'h2a == index | valid_0_42; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8074 = 6'h2b == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_564 = 6'h2b == index | valid_0_43; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8075 = 6'h2c == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_565 = 6'h2c == index | valid_0_44; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8076 = 6'h2d == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_566 = 6'h2d == index | valid_0_45; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8077 = 6'h2e == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_567 = 6'h2e == index | valid_0_46; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8078 = 6'h2f == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_568 = 6'h2f == index | valid_0_47; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8079 = 6'h30 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_569 = 6'h30 == index | valid_0_48; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8080 = 6'h31 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_570 = 6'h31 == index | valid_0_49; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8081 = 6'h32 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_571 = 6'h32 == index | valid_0_50; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8082 = 6'h33 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_572 = 6'h33 == index | valid_0_51; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8083 = 6'h34 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_573 = 6'h34 == index | valid_0_52; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8084 = 6'h35 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_574 = 6'h35 == index | valid_0_53; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8085 = 6'h36 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_575 = 6'h36 == index | valid_0_54; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8086 = 6'h37 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_576 = 6'h37 == index | valid_0_55; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8087 = 6'h38 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_577 = 6'h38 == index | valid_0_56; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8088 = 6'h39 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_578 = 6'h39 == index | valid_0_57; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8089 = 6'h3a == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_579 = 6'h3a == index | valid_0_58; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8090 = 6'h3b == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_580 = 6'h3b == index | valid_0_59; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8091 = 6'h3c == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_581 = 6'h3c == index | valid_0_60; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8092 = 6'h3d == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_582 = 6'h3d == index | valid_0_61; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8093 = 6'h3e == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_583 = 6'h3e == index | valid_0_62; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_8094 = 6'h3f == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_584 = 6'h3f == index | valid_0_63; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_585 = _GEN_8031 | dirty_0_0; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_586 = _GEN_8032 | dirty_0_1; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_587 = _GEN_8033 | dirty_0_2; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_588 = _GEN_8034 | dirty_0_3; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_589 = _GEN_8035 | dirty_0_4; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_590 = _GEN_8036 | dirty_0_5; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_591 = _GEN_8037 | dirty_0_6; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_592 = _GEN_8038 | dirty_0_7; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_593 = _GEN_8039 | dirty_0_8; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_594 = _GEN_8040 | dirty_0_9; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_595 = _GEN_8041 | dirty_0_10; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_596 = _GEN_8042 | dirty_0_11; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_597 = _GEN_8043 | dirty_0_12; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_598 = _GEN_8044 | dirty_0_13; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_599 = _GEN_8045 | dirty_0_14; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_600 = _GEN_8046 | dirty_0_15; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_601 = _GEN_8047 | dirty_0_16; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_602 = _GEN_8048 | dirty_0_17; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_603 = _GEN_8049 | dirty_0_18; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_604 = _GEN_8050 | dirty_0_19; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_605 = _GEN_8051 | dirty_0_20; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_606 = _GEN_8052 | dirty_0_21; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_607 = _GEN_8053 | dirty_0_22; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_608 = _GEN_8054 | dirty_0_23; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_609 = _GEN_8055 | dirty_0_24; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_610 = _GEN_8056 | dirty_0_25; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_611 = _GEN_8057 | dirty_0_26; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_612 = _GEN_8058 | dirty_0_27; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_613 = _GEN_8059 | dirty_0_28; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_614 = _GEN_8060 | dirty_0_29; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_615 = _GEN_8061 | dirty_0_30; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_616 = _GEN_8062 | dirty_0_31; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_617 = _GEN_8063 | dirty_0_32; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_618 = _GEN_8064 | dirty_0_33; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_619 = _GEN_8065 | dirty_0_34; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_620 = _GEN_8066 | dirty_0_35; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_621 = _GEN_8067 | dirty_0_36; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_622 = _GEN_8068 | dirty_0_37; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_623 = _GEN_8069 | dirty_0_38; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_624 = _GEN_8070 | dirty_0_39; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_625 = _GEN_8071 | dirty_0_40; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_626 = _GEN_8072 | dirty_0_41; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_627 = _GEN_8073 | dirty_0_42; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_628 = _GEN_8074 | dirty_0_43; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_629 = _GEN_8075 | dirty_0_44; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_630 = _GEN_8076 | dirty_0_45; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_631 = _GEN_8077 | dirty_0_46; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_632 = _GEN_8078 | dirty_0_47; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_633 = _GEN_8079 | dirty_0_48; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_634 = _GEN_8080 | dirty_0_49; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_635 = _GEN_8081 | dirty_0_50; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_636 = _GEN_8082 | dirty_0_51; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_637 = _GEN_8083 | dirty_0_52; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_638 = _GEN_8084 | dirty_0_53; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_639 = _GEN_8085 | dirty_0_54; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_640 = _GEN_8086 | dirty_0_55; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_641 = _GEN_8087 | dirty_0_56; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_642 = _GEN_8088 | dirty_0_57; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_643 = _GEN_8089 | dirty_0_58; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_644 = _GEN_8090 | dirty_0_59; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_645 = _GEN_8091 | dirty_0_60; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_646 = _GEN_8092 | dirty_0_61; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_647 = _GEN_8093 | dirty_0_62; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_648 = _GEN_8094 | dirty_0_63; // @[d_cache.scala 113:{32,32} 26:26]
  wire [63:0] _GEN_650 = 6'h1 == index ? ram_1_1 : ram_1_0; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_651 = 6'h2 == index ? ram_1_2 : _GEN_650; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_652 = 6'h3 == index ? ram_1_3 : _GEN_651; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_653 = 6'h4 == index ? ram_1_4 : _GEN_652; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_654 = 6'h5 == index ? ram_1_5 : _GEN_653; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_655 = 6'h6 == index ? ram_1_6 : _GEN_654; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_656 = 6'h7 == index ? ram_1_7 : _GEN_655; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_657 = 6'h8 == index ? ram_1_8 : _GEN_656; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_658 = 6'h9 == index ? ram_1_9 : _GEN_657; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_659 = 6'ha == index ? ram_1_10 : _GEN_658; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_660 = 6'hb == index ? ram_1_11 : _GEN_659; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_661 = 6'hc == index ? ram_1_12 : _GEN_660; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_662 = 6'hd == index ? ram_1_13 : _GEN_661; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_663 = 6'he == index ? ram_1_14 : _GEN_662; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_664 = 6'hf == index ? ram_1_15 : _GEN_663; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_665 = 6'h10 == index ? ram_1_16 : _GEN_664; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_666 = 6'h11 == index ? ram_1_17 : _GEN_665; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_667 = 6'h12 == index ? ram_1_18 : _GEN_666; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_668 = 6'h13 == index ? ram_1_19 : _GEN_667; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_669 = 6'h14 == index ? ram_1_20 : _GEN_668; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_670 = 6'h15 == index ? ram_1_21 : _GEN_669; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_671 = 6'h16 == index ? ram_1_22 : _GEN_670; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_672 = 6'h17 == index ? ram_1_23 : _GEN_671; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_673 = 6'h18 == index ? ram_1_24 : _GEN_672; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_674 = 6'h19 == index ? ram_1_25 : _GEN_673; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_675 = 6'h1a == index ? ram_1_26 : _GEN_674; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_676 = 6'h1b == index ? ram_1_27 : _GEN_675; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_677 = 6'h1c == index ? ram_1_28 : _GEN_676; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_678 = 6'h1d == index ? ram_1_29 : _GEN_677; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_679 = 6'h1e == index ? ram_1_30 : _GEN_678; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_680 = 6'h1f == index ? ram_1_31 : _GEN_679; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_681 = 6'h20 == index ? ram_1_32 : _GEN_680; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_682 = 6'h21 == index ? ram_1_33 : _GEN_681; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_683 = 6'h22 == index ? ram_1_34 : _GEN_682; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_684 = 6'h23 == index ? ram_1_35 : _GEN_683; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_685 = 6'h24 == index ? ram_1_36 : _GEN_684; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_686 = 6'h25 == index ? ram_1_37 : _GEN_685; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_687 = 6'h26 == index ? ram_1_38 : _GEN_686; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_688 = 6'h27 == index ? ram_1_39 : _GEN_687; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_689 = 6'h28 == index ? ram_1_40 : _GEN_688; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_690 = 6'h29 == index ? ram_1_41 : _GEN_689; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_691 = 6'h2a == index ? ram_1_42 : _GEN_690; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_692 = 6'h2b == index ? ram_1_43 : _GEN_691; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_693 = 6'h2c == index ? ram_1_44 : _GEN_692; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_694 = 6'h2d == index ? ram_1_45 : _GEN_693; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_695 = 6'h2e == index ? ram_1_46 : _GEN_694; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_696 = 6'h2f == index ? ram_1_47 : _GEN_695; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_697 = 6'h30 == index ? ram_1_48 : _GEN_696; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_698 = 6'h31 == index ? ram_1_49 : _GEN_697; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_699 = 6'h32 == index ? ram_1_50 : _GEN_698; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_700 = 6'h33 == index ? ram_1_51 : _GEN_699; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_701 = 6'h34 == index ? ram_1_52 : _GEN_700; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_702 = 6'h35 == index ? ram_1_53 : _GEN_701; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_703 = 6'h36 == index ? ram_1_54 : _GEN_702; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_704 = 6'h37 == index ? ram_1_55 : _GEN_703; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_705 = 6'h38 == index ? ram_1_56 : _GEN_704; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_706 = 6'h39 == index ? ram_1_57 : _GEN_705; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_707 = 6'h3a == index ? ram_1_58 : _GEN_706; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_708 = 6'h3b == index ? ram_1_59 : _GEN_707; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_709 = 6'h3c == index ? ram_1_60 : _GEN_708; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_710 = 6'h3d == index ? ram_1_61 : _GEN_709; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_711 = 6'h3e == index ? ram_1_62 : _GEN_710; // @[d_cache.scala 118:{92,92}]
  wire [63:0] _GEN_712 = 6'h3f == index ? ram_1_63 : _GEN_711; // @[d_cache.scala 118:{92,92}]
  wire [126:0] _GEN_8160 = {{63'd0}, _GEN_712}; // @[d_cache.scala 118:92]
  wire [126:0] _ram_1_T_4 = _GEN_8160 & _ram_0_T_3; // @[d_cache.scala 118:92]
  wire [126:0] _ram_1_T_5 = _ram_0_T_1 | _ram_1_T_4; // @[d_cache.scala 118:76]
  wire [63:0] _GEN_713 = 6'h0 == index ? _ram_1_T_5[63:0] : ram_1_0; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_714 = 6'h1 == index ? _ram_1_T_5[63:0] : ram_1_1; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_715 = 6'h2 == index ? _ram_1_T_5[63:0] : ram_1_2; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_716 = 6'h3 == index ? _ram_1_T_5[63:0] : ram_1_3; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_717 = 6'h4 == index ? _ram_1_T_5[63:0] : ram_1_4; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_718 = 6'h5 == index ? _ram_1_T_5[63:0] : ram_1_5; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_719 = 6'h6 == index ? _ram_1_T_5[63:0] : ram_1_6; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_720 = 6'h7 == index ? _ram_1_T_5[63:0] : ram_1_7; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_721 = 6'h8 == index ? _ram_1_T_5[63:0] : ram_1_8; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_722 = 6'h9 == index ? _ram_1_T_5[63:0] : ram_1_9; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_723 = 6'ha == index ? _ram_1_T_5[63:0] : ram_1_10; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_724 = 6'hb == index ? _ram_1_T_5[63:0] : ram_1_11; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_725 = 6'hc == index ? _ram_1_T_5[63:0] : ram_1_12; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_726 = 6'hd == index ? _ram_1_T_5[63:0] : ram_1_13; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_727 = 6'he == index ? _ram_1_T_5[63:0] : ram_1_14; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_728 = 6'hf == index ? _ram_1_T_5[63:0] : ram_1_15; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_729 = 6'h10 == index ? _ram_1_T_5[63:0] : ram_1_16; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_730 = 6'h11 == index ? _ram_1_T_5[63:0] : ram_1_17; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_731 = 6'h12 == index ? _ram_1_T_5[63:0] : ram_1_18; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_732 = 6'h13 == index ? _ram_1_T_5[63:0] : ram_1_19; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_733 = 6'h14 == index ? _ram_1_T_5[63:0] : ram_1_20; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_734 = 6'h15 == index ? _ram_1_T_5[63:0] : ram_1_21; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_735 = 6'h16 == index ? _ram_1_T_5[63:0] : ram_1_22; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_736 = 6'h17 == index ? _ram_1_T_5[63:0] : ram_1_23; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_737 = 6'h18 == index ? _ram_1_T_5[63:0] : ram_1_24; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_738 = 6'h19 == index ? _ram_1_T_5[63:0] : ram_1_25; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_739 = 6'h1a == index ? _ram_1_T_5[63:0] : ram_1_26; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_740 = 6'h1b == index ? _ram_1_T_5[63:0] : ram_1_27; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_741 = 6'h1c == index ? _ram_1_T_5[63:0] : ram_1_28; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_742 = 6'h1d == index ? _ram_1_T_5[63:0] : ram_1_29; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_743 = 6'h1e == index ? _ram_1_T_5[63:0] : ram_1_30; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_744 = 6'h1f == index ? _ram_1_T_5[63:0] : ram_1_31; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_745 = 6'h20 == index ? _ram_1_T_5[63:0] : ram_1_32; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_746 = 6'h21 == index ? _ram_1_T_5[63:0] : ram_1_33; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_747 = 6'h22 == index ? _ram_1_T_5[63:0] : ram_1_34; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_748 = 6'h23 == index ? _ram_1_T_5[63:0] : ram_1_35; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_749 = 6'h24 == index ? _ram_1_T_5[63:0] : ram_1_36; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_750 = 6'h25 == index ? _ram_1_T_5[63:0] : ram_1_37; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_751 = 6'h26 == index ? _ram_1_T_5[63:0] : ram_1_38; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_752 = 6'h27 == index ? _ram_1_T_5[63:0] : ram_1_39; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_753 = 6'h28 == index ? _ram_1_T_5[63:0] : ram_1_40; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_754 = 6'h29 == index ? _ram_1_T_5[63:0] : ram_1_41; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_755 = 6'h2a == index ? _ram_1_T_5[63:0] : ram_1_42; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_756 = 6'h2b == index ? _ram_1_T_5[63:0] : ram_1_43; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_757 = 6'h2c == index ? _ram_1_T_5[63:0] : ram_1_44; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_758 = 6'h2d == index ? _ram_1_T_5[63:0] : ram_1_45; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_759 = 6'h2e == index ? _ram_1_T_5[63:0] : ram_1_46; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_760 = 6'h2f == index ? _ram_1_T_5[63:0] : ram_1_47; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_761 = 6'h30 == index ? _ram_1_T_5[63:0] : ram_1_48; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_762 = 6'h31 == index ? _ram_1_T_5[63:0] : ram_1_49; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_763 = 6'h32 == index ? _ram_1_T_5[63:0] : ram_1_50; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_764 = 6'h33 == index ? _ram_1_T_5[63:0] : ram_1_51; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_765 = 6'h34 == index ? _ram_1_T_5[63:0] : ram_1_52; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_766 = 6'h35 == index ? _ram_1_T_5[63:0] : ram_1_53; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_767 = 6'h36 == index ? _ram_1_T_5[63:0] : ram_1_54; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_768 = 6'h37 == index ? _ram_1_T_5[63:0] : ram_1_55; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_769 = 6'h38 == index ? _ram_1_T_5[63:0] : ram_1_56; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_770 = 6'h39 == index ? _ram_1_T_5[63:0] : ram_1_57; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_771 = 6'h3a == index ? _ram_1_T_5[63:0] : ram_1_58; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_772 = 6'h3b == index ? _ram_1_T_5[63:0] : ram_1_59; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_773 = 6'h3c == index ? _ram_1_T_5[63:0] : ram_1_60; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_774 = 6'h3d == index ? _ram_1_T_5[63:0] : ram_1_61; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_775 = 6'h3e == index ? _ram_1_T_5[63:0] : ram_1_62; // @[d_cache.scala 118:{30,30} 19:24]
  wire [63:0] _GEN_776 = 6'h3f == index ? _ram_1_T_5[63:0] : ram_1_63; // @[d_cache.scala 118:{30,30} 19:24]
  wire  _GEN_777 = _GEN_8031 | valid_1_0; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_778 = _GEN_8032 | valid_1_1; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_779 = _GEN_8033 | valid_1_2; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_780 = _GEN_8034 | valid_1_3; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_781 = _GEN_8035 | valid_1_4; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_782 = _GEN_8036 | valid_1_5; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_783 = _GEN_8037 | valid_1_6; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_784 = _GEN_8038 | valid_1_7; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_785 = _GEN_8039 | valid_1_8; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_786 = _GEN_8040 | valid_1_9; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_787 = _GEN_8041 | valid_1_10; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_788 = _GEN_8042 | valid_1_11; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_789 = _GEN_8043 | valid_1_12; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_790 = _GEN_8044 | valid_1_13; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_791 = _GEN_8045 | valid_1_14; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_792 = _GEN_8046 | valid_1_15; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_793 = _GEN_8047 | valid_1_16; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_794 = _GEN_8048 | valid_1_17; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_795 = _GEN_8049 | valid_1_18; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_796 = _GEN_8050 | valid_1_19; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_797 = _GEN_8051 | valid_1_20; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_798 = _GEN_8052 | valid_1_21; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_799 = _GEN_8053 | valid_1_22; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_800 = _GEN_8054 | valid_1_23; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_801 = _GEN_8055 | valid_1_24; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_802 = _GEN_8056 | valid_1_25; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_803 = _GEN_8057 | valid_1_26; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_804 = _GEN_8058 | valid_1_27; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_805 = _GEN_8059 | valid_1_28; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_806 = _GEN_8060 | valid_1_29; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_807 = _GEN_8061 | valid_1_30; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_808 = _GEN_8062 | valid_1_31; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_809 = _GEN_8063 | valid_1_32; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_810 = _GEN_8064 | valid_1_33; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_811 = _GEN_8065 | valid_1_34; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_812 = _GEN_8066 | valid_1_35; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_813 = _GEN_8067 | valid_1_36; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_814 = _GEN_8068 | valid_1_37; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_815 = _GEN_8069 | valid_1_38; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_816 = _GEN_8070 | valid_1_39; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_817 = _GEN_8071 | valid_1_40; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_818 = _GEN_8072 | valid_1_41; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_819 = _GEN_8073 | valid_1_42; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_820 = _GEN_8074 | valid_1_43; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_821 = _GEN_8075 | valid_1_44; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_822 = _GEN_8076 | valid_1_45; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_823 = _GEN_8077 | valid_1_46; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_824 = _GEN_8078 | valid_1_47; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_825 = _GEN_8079 | valid_1_48; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_826 = _GEN_8080 | valid_1_49; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_827 = _GEN_8081 | valid_1_50; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_828 = _GEN_8082 | valid_1_51; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_829 = _GEN_8083 | valid_1_52; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_830 = _GEN_8084 | valid_1_53; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_831 = _GEN_8085 | valid_1_54; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_832 = _GEN_8086 | valid_1_55; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_833 = _GEN_8087 | valid_1_56; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_834 = _GEN_8088 | valid_1_57; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_835 = _GEN_8089 | valid_1_58; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_836 = _GEN_8090 | valid_1_59; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_837 = _GEN_8091 | valid_1_60; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_838 = _GEN_8092 | valid_1_61; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_839 = _GEN_8093 | valid_1_62; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_840 = _GEN_8094 | valid_1_63; // @[d_cache.scala 119:{32,32} 25:26]
  wire  _GEN_841 = _GEN_8031 | dirty_1_0; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_842 = _GEN_8032 | dirty_1_1; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_843 = _GEN_8033 | dirty_1_2; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_844 = _GEN_8034 | dirty_1_3; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_845 = _GEN_8035 | dirty_1_4; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_846 = _GEN_8036 | dirty_1_5; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_847 = _GEN_8037 | dirty_1_6; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_848 = _GEN_8038 | dirty_1_7; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_849 = _GEN_8039 | dirty_1_8; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_850 = _GEN_8040 | dirty_1_9; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_851 = _GEN_8041 | dirty_1_10; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_852 = _GEN_8042 | dirty_1_11; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_853 = _GEN_8043 | dirty_1_12; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_854 = _GEN_8044 | dirty_1_13; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_855 = _GEN_8045 | dirty_1_14; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_856 = _GEN_8046 | dirty_1_15; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_857 = _GEN_8047 | dirty_1_16; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_858 = _GEN_8048 | dirty_1_17; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_859 = _GEN_8049 | dirty_1_18; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_860 = _GEN_8050 | dirty_1_19; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_861 = _GEN_8051 | dirty_1_20; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_862 = _GEN_8052 | dirty_1_21; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_863 = _GEN_8053 | dirty_1_22; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_864 = _GEN_8054 | dirty_1_23; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_865 = _GEN_8055 | dirty_1_24; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_866 = _GEN_8056 | dirty_1_25; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_867 = _GEN_8057 | dirty_1_26; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_868 = _GEN_8058 | dirty_1_27; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_869 = _GEN_8059 | dirty_1_28; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_870 = _GEN_8060 | dirty_1_29; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_871 = _GEN_8061 | dirty_1_30; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_872 = _GEN_8062 | dirty_1_31; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_873 = _GEN_8063 | dirty_1_32; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_874 = _GEN_8064 | dirty_1_33; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_875 = _GEN_8065 | dirty_1_34; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_876 = _GEN_8066 | dirty_1_35; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_877 = _GEN_8067 | dirty_1_36; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_878 = _GEN_8068 | dirty_1_37; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_879 = _GEN_8069 | dirty_1_38; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_880 = _GEN_8070 | dirty_1_39; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_881 = _GEN_8071 | dirty_1_40; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_882 = _GEN_8072 | dirty_1_41; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_883 = _GEN_8073 | dirty_1_42; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_884 = _GEN_8074 | dirty_1_43; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_885 = _GEN_8075 | dirty_1_44; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_886 = _GEN_8076 | dirty_1_45; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_887 = _GEN_8077 | dirty_1_46; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_888 = _GEN_8078 | dirty_1_47; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_889 = _GEN_8079 | dirty_1_48; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_890 = _GEN_8080 | dirty_1_49; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_891 = _GEN_8081 | dirty_1_50; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_892 = _GEN_8082 | dirty_1_51; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_893 = _GEN_8083 | dirty_1_52; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_894 = _GEN_8084 | dirty_1_53; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_895 = _GEN_8085 | dirty_1_54; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_896 = _GEN_8086 | dirty_1_55; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_897 = _GEN_8087 | dirty_1_56; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_898 = _GEN_8088 | dirty_1_57; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_899 = _GEN_8089 | dirty_1_58; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_900 = _GEN_8090 | dirty_1_59; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_901 = _GEN_8091 | dirty_1_60; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_902 = _GEN_8092 | dirty_1_61; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_903 = _GEN_8093 | dirty_1_62; // @[d_cache.scala 121:{32,32} 27:26]
  wire  _GEN_904 = _GEN_8094 | dirty_1_63; // @[d_cache.scala 121:{32,32} 27:26]
  wire [2:0] _GEN_905 = way1_hit ? 3'h0 : 3'h4; // @[d_cache.scala 116:33 117:23 124:23]
  wire [63:0] _GEN_906 = way1_hit ? _GEN_713 : ram_1_0; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_907 = way1_hit ? _GEN_714 : ram_1_1; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_908 = way1_hit ? _GEN_715 : ram_1_2; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_909 = way1_hit ? _GEN_716 : ram_1_3; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_910 = way1_hit ? _GEN_717 : ram_1_4; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_911 = way1_hit ? _GEN_718 : ram_1_5; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_912 = way1_hit ? _GEN_719 : ram_1_6; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_913 = way1_hit ? _GEN_720 : ram_1_7; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_914 = way1_hit ? _GEN_721 : ram_1_8; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_915 = way1_hit ? _GEN_722 : ram_1_9; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_916 = way1_hit ? _GEN_723 : ram_1_10; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_917 = way1_hit ? _GEN_724 : ram_1_11; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_918 = way1_hit ? _GEN_725 : ram_1_12; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_919 = way1_hit ? _GEN_726 : ram_1_13; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_920 = way1_hit ? _GEN_727 : ram_1_14; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_921 = way1_hit ? _GEN_728 : ram_1_15; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_922 = way1_hit ? _GEN_729 : ram_1_16; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_923 = way1_hit ? _GEN_730 : ram_1_17; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_924 = way1_hit ? _GEN_731 : ram_1_18; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_925 = way1_hit ? _GEN_732 : ram_1_19; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_926 = way1_hit ? _GEN_733 : ram_1_20; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_927 = way1_hit ? _GEN_734 : ram_1_21; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_928 = way1_hit ? _GEN_735 : ram_1_22; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_929 = way1_hit ? _GEN_736 : ram_1_23; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_930 = way1_hit ? _GEN_737 : ram_1_24; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_931 = way1_hit ? _GEN_738 : ram_1_25; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_932 = way1_hit ? _GEN_739 : ram_1_26; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_933 = way1_hit ? _GEN_740 : ram_1_27; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_934 = way1_hit ? _GEN_741 : ram_1_28; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_935 = way1_hit ? _GEN_742 : ram_1_29; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_936 = way1_hit ? _GEN_743 : ram_1_30; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_937 = way1_hit ? _GEN_744 : ram_1_31; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_938 = way1_hit ? _GEN_745 : ram_1_32; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_939 = way1_hit ? _GEN_746 : ram_1_33; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_940 = way1_hit ? _GEN_747 : ram_1_34; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_941 = way1_hit ? _GEN_748 : ram_1_35; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_942 = way1_hit ? _GEN_749 : ram_1_36; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_943 = way1_hit ? _GEN_750 : ram_1_37; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_944 = way1_hit ? _GEN_751 : ram_1_38; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_945 = way1_hit ? _GEN_752 : ram_1_39; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_946 = way1_hit ? _GEN_753 : ram_1_40; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_947 = way1_hit ? _GEN_754 : ram_1_41; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_948 = way1_hit ? _GEN_755 : ram_1_42; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_949 = way1_hit ? _GEN_756 : ram_1_43; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_950 = way1_hit ? _GEN_757 : ram_1_44; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_951 = way1_hit ? _GEN_758 : ram_1_45; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_952 = way1_hit ? _GEN_759 : ram_1_46; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_953 = way1_hit ? _GEN_760 : ram_1_47; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_954 = way1_hit ? _GEN_761 : ram_1_48; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_955 = way1_hit ? _GEN_762 : ram_1_49; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_956 = way1_hit ? _GEN_763 : ram_1_50; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_957 = way1_hit ? _GEN_764 : ram_1_51; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_958 = way1_hit ? _GEN_765 : ram_1_52; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_959 = way1_hit ? _GEN_766 : ram_1_53; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_960 = way1_hit ? _GEN_767 : ram_1_54; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_961 = way1_hit ? _GEN_768 : ram_1_55; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_962 = way1_hit ? _GEN_769 : ram_1_56; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_963 = way1_hit ? _GEN_770 : ram_1_57; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_964 = way1_hit ? _GEN_771 : ram_1_58; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_965 = way1_hit ? _GEN_772 : ram_1_59; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_966 = way1_hit ? _GEN_773 : ram_1_60; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_967 = way1_hit ? _GEN_774 : ram_1_61; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_968 = way1_hit ? _GEN_775 : ram_1_62; // @[d_cache.scala 116:33 19:24]
  wire [63:0] _GEN_969 = way1_hit ? _GEN_776 : ram_1_63; // @[d_cache.scala 116:33 19:24]
  wire  _GEN_970 = way1_hit ? _GEN_777 : valid_1_0; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_971 = way1_hit ? _GEN_778 : valid_1_1; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_972 = way1_hit ? _GEN_779 : valid_1_2; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_973 = way1_hit ? _GEN_780 : valid_1_3; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_974 = way1_hit ? _GEN_781 : valid_1_4; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_975 = way1_hit ? _GEN_782 : valid_1_5; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_976 = way1_hit ? _GEN_783 : valid_1_6; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_977 = way1_hit ? _GEN_784 : valid_1_7; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_978 = way1_hit ? _GEN_785 : valid_1_8; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_979 = way1_hit ? _GEN_786 : valid_1_9; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_980 = way1_hit ? _GEN_787 : valid_1_10; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_981 = way1_hit ? _GEN_788 : valid_1_11; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_982 = way1_hit ? _GEN_789 : valid_1_12; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_983 = way1_hit ? _GEN_790 : valid_1_13; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_984 = way1_hit ? _GEN_791 : valid_1_14; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_985 = way1_hit ? _GEN_792 : valid_1_15; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_986 = way1_hit ? _GEN_793 : valid_1_16; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_987 = way1_hit ? _GEN_794 : valid_1_17; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_988 = way1_hit ? _GEN_795 : valid_1_18; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_989 = way1_hit ? _GEN_796 : valid_1_19; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_990 = way1_hit ? _GEN_797 : valid_1_20; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_991 = way1_hit ? _GEN_798 : valid_1_21; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_992 = way1_hit ? _GEN_799 : valid_1_22; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_993 = way1_hit ? _GEN_800 : valid_1_23; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_994 = way1_hit ? _GEN_801 : valid_1_24; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_995 = way1_hit ? _GEN_802 : valid_1_25; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_996 = way1_hit ? _GEN_803 : valid_1_26; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_997 = way1_hit ? _GEN_804 : valid_1_27; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_998 = way1_hit ? _GEN_805 : valid_1_28; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_999 = way1_hit ? _GEN_806 : valid_1_29; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1000 = way1_hit ? _GEN_807 : valid_1_30; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1001 = way1_hit ? _GEN_808 : valid_1_31; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1002 = way1_hit ? _GEN_809 : valid_1_32; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1003 = way1_hit ? _GEN_810 : valid_1_33; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1004 = way1_hit ? _GEN_811 : valid_1_34; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1005 = way1_hit ? _GEN_812 : valid_1_35; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1006 = way1_hit ? _GEN_813 : valid_1_36; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1007 = way1_hit ? _GEN_814 : valid_1_37; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1008 = way1_hit ? _GEN_815 : valid_1_38; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1009 = way1_hit ? _GEN_816 : valid_1_39; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1010 = way1_hit ? _GEN_817 : valid_1_40; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1011 = way1_hit ? _GEN_818 : valid_1_41; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1012 = way1_hit ? _GEN_819 : valid_1_42; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1013 = way1_hit ? _GEN_820 : valid_1_43; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1014 = way1_hit ? _GEN_821 : valid_1_44; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1015 = way1_hit ? _GEN_822 : valid_1_45; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1016 = way1_hit ? _GEN_823 : valid_1_46; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1017 = way1_hit ? _GEN_824 : valid_1_47; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1018 = way1_hit ? _GEN_825 : valid_1_48; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1019 = way1_hit ? _GEN_826 : valid_1_49; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1020 = way1_hit ? _GEN_827 : valid_1_50; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1021 = way1_hit ? _GEN_828 : valid_1_51; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1022 = way1_hit ? _GEN_829 : valid_1_52; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1023 = way1_hit ? _GEN_830 : valid_1_53; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1024 = way1_hit ? _GEN_831 : valid_1_54; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1025 = way1_hit ? _GEN_832 : valid_1_55; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1026 = way1_hit ? _GEN_833 : valid_1_56; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1027 = way1_hit ? _GEN_834 : valid_1_57; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1028 = way1_hit ? _GEN_835 : valid_1_58; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1029 = way1_hit ? _GEN_836 : valid_1_59; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1030 = way1_hit ? _GEN_837 : valid_1_60; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1031 = way1_hit ? _GEN_838 : valid_1_61; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1032 = way1_hit ? _GEN_839 : valid_1_62; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1033 = way1_hit ? _GEN_840 : valid_1_63; // @[d_cache.scala 116:33 25:26]
  wire  _GEN_1034 = way1_hit ? _GEN_841 : dirty_1_0; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1035 = way1_hit ? _GEN_842 : dirty_1_1; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1036 = way1_hit ? _GEN_843 : dirty_1_2; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1037 = way1_hit ? _GEN_844 : dirty_1_3; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1038 = way1_hit ? _GEN_845 : dirty_1_4; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1039 = way1_hit ? _GEN_846 : dirty_1_5; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1040 = way1_hit ? _GEN_847 : dirty_1_6; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1041 = way1_hit ? _GEN_848 : dirty_1_7; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1042 = way1_hit ? _GEN_849 : dirty_1_8; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1043 = way1_hit ? _GEN_850 : dirty_1_9; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1044 = way1_hit ? _GEN_851 : dirty_1_10; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1045 = way1_hit ? _GEN_852 : dirty_1_11; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1046 = way1_hit ? _GEN_853 : dirty_1_12; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1047 = way1_hit ? _GEN_854 : dirty_1_13; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1048 = way1_hit ? _GEN_855 : dirty_1_14; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1049 = way1_hit ? _GEN_856 : dirty_1_15; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1050 = way1_hit ? _GEN_857 : dirty_1_16; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1051 = way1_hit ? _GEN_858 : dirty_1_17; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1052 = way1_hit ? _GEN_859 : dirty_1_18; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1053 = way1_hit ? _GEN_860 : dirty_1_19; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1054 = way1_hit ? _GEN_861 : dirty_1_20; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1055 = way1_hit ? _GEN_862 : dirty_1_21; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1056 = way1_hit ? _GEN_863 : dirty_1_22; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1057 = way1_hit ? _GEN_864 : dirty_1_23; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1058 = way1_hit ? _GEN_865 : dirty_1_24; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1059 = way1_hit ? _GEN_866 : dirty_1_25; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1060 = way1_hit ? _GEN_867 : dirty_1_26; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1061 = way1_hit ? _GEN_868 : dirty_1_27; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1062 = way1_hit ? _GEN_869 : dirty_1_28; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1063 = way1_hit ? _GEN_870 : dirty_1_29; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1064 = way1_hit ? _GEN_871 : dirty_1_30; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1065 = way1_hit ? _GEN_872 : dirty_1_31; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1066 = way1_hit ? _GEN_873 : dirty_1_32; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1067 = way1_hit ? _GEN_874 : dirty_1_33; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1068 = way1_hit ? _GEN_875 : dirty_1_34; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1069 = way1_hit ? _GEN_876 : dirty_1_35; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1070 = way1_hit ? _GEN_877 : dirty_1_36; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1071 = way1_hit ? _GEN_878 : dirty_1_37; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1072 = way1_hit ? _GEN_879 : dirty_1_38; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1073 = way1_hit ? _GEN_880 : dirty_1_39; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1074 = way1_hit ? _GEN_881 : dirty_1_40; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1075 = way1_hit ? _GEN_882 : dirty_1_41; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1076 = way1_hit ? _GEN_883 : dirty_1_42; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1077 = way1_hit ? _GEN_884 : dirty_1_43; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1078 = way1_hit ? _GEN_885 : dirty_1_44; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1079 = way1_hit ? _GEN_886 : dirty_1_45; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1080 = way1_hit ? _GEN_887 : dirty_1_46; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1081 = way1_hit ? _GEN_888 : dirty_1_47; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1082 = way1_hit ? _GEN_889 : dirty_1_48; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1083 = way1_hit ? _GEN_890 : dirty_1_49; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1084 = way1_hit ? _GEN_891 : dirty_1_50; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1085 = way1_hit ? _GEN_892 : dirty_1_51; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1086 = way1_hit ? _GEN_893 : dirty_1_52; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1087 = way1_hit ? _GEN_894 : dirty_1_53; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1088 = way1_hit ? _GEN_895 : dirty_1_54; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1089 = way1_hit ? _GEN_896 : dirty_1_55; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1090 = way1_hit ? _GEN_897 : dirty_1_56; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1091 = way1_hit ? _GEN_898 : dirty_1_57; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1092 = way1_hit ? _GEN_899 : dirty_1_58; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1093 = way1_hit ? _GEN_900 : dirty_1_59; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1094 = way1_hit ? _GEN_901 : dirty_1_60; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1095 = way1_hit ? _GEN_902 : dirty_1_61; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1096 = way1_hit ? _GEN_903 : dirty_1_62; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1097 = way1_hit ? _GEN_904 : dirty_1_63; // @[d_cache.scala 116:33 27:26]
  wire  _GEN_1098 = way1_hit ? 1'h0 : quene; // @[d_cache.scala 116:33 122:23 37:24]
  wire [2:0] _GEN_1099 = way0_hit ? 3'h0 : _GEN_905; // @[d_cache.scala 107:27 108:23]
  wire [63:0] _GEN_1100 = way0_hit ? _GEN_457 : ram_0_0; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1101 = way0_hit ? _GEN_458 : ram_0_1; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1102 = way0_hit ? _GEN_459 : ram_0_2; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1103 = way0_hit ? _GEN_460 : ram_0_3; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1104 = way0_hit ? _GEN_461 : ram_0_4; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1105 = way0_hit ? _GEN_462 : ram_0_5; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1106 = way0_hit ? _GEN_463 : ram_0_6; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1107 = way0_hit ? _GEN_464 : ram_0_7; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1108 = way0_hit ? _GEN_465 : ram_0_8; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1109 = way0_hit ? _GEN_466 : ram_0_9; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1110 = way0_hit ? _GEN_467 : ram_0_10; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1111 = way0_hit ? _GEN_468 : ram_0_11; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1112 = way0_hit ? _GEN_469 : ram_0_12; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1113 = way0_hit ? _GEN_470 : ram_0_13; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1114 = way0_hit ? _GEN_471 : ram_0_14; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1115 = way0_hit ? _GEN_472 : ram_0_15; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1116 = way0_hit ? _GEN_473 : ram_0_16; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1117 = way0_hit ? _GEN_474 : ram_0_17; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1118 = way0_hit ? _GEN_475 : ram_0_18; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1119 = way0_hit ? _GEN_476 : ram_0_19; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1120 = way0_hit ? _GEN_477 : ram_0_20; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1121 = way0_hit ? _GEN_478 : ram_0_21; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1122 = way0_hit ? _GEN_479 : ram_0_22; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1123 = way0_hit ? _GEN_480 : ram_0_23; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1124 = way0_hit ? _GEN_481 : ram_0_24; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1125 = way0_hit ? _GEN_482 : ram_0_25; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1126 = way0_hit ? _GEN_483 : ram_0_26; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1127 = way0_hit ? _GEN_484 : ram_0_27; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1128 = way0_hit ? _GEN_485 : ram_0_28; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1129 = way0_hit ? _GEN_486 : ram_0_29; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1130 = way0_hit ? _GEN_487 : ram_0_30; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1131 = way0_hit ? _GEN_488 : ram_0_31; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1132 = way0_hit ? _GEN_489 : ram_0_32; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1133 = way0_hit ? _GEN_490 : ram_0_33; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1134 = way0_hit ? _GEN_491 : ram_0_34; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1135 = way0_hit ? _GEN_492 : ram_0_35; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1136 = way0_hit ? _GEN_493 : ram_0_36; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1137 = way0_hit ? _GEN_494 : ram_0_37; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1138 = way0_hit ? _GEN_495 : ram_0_38; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1139 = way0_hit ? _GEN_496 : ram_0_39; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1140 = way0_hit ? _GEN_497 : ram_0_40; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1141 = way0_hit ? _GEN_498 : ram_0_41; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1142 = way0_hit ? _GEN_499 : ram_0_42; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1143 = way0_hit ? _GEN_500 : ram_0_43; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1144 = way0_hit ? _GEN_501 : ram_0_44; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1145 = way0_hit ? _GEN_502 : ram_0_45; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1146 = way0_hit ? _GEN_503 : ram_0_46; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1147 = way0_hit ? _GEN_504 : ram_0_47; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1148 = way0_hit ? _GEN_505 : ram_0_48; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1149 = way0_hit ? _GEN_506 : ram_0_49; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1150 = way0_hit ? _GEN_507 : ram_0_50; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1151 = way0_hit ? _GEN_508 : ram_0_51; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1152 = way0_hit ? _GEN_509 : ram_0_52; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1153 = way0_hit ? _GEN_510 : ram_0_53; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1154 = way0_hit ? _GEN_511 : ram_0_54; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1155 = way0_hit ? _GEN_512 : ram_0_55; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1156 = way0_hit ? _GEN_513 : ram_0_56; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1157 = way0_hit ? _GEN_514 : ram_0_57; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1158 = way0_hit ? _GEN_515 : ram_0_58; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1159 = way0_hit ? _GEN_516 : ram_0_59; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1160 = way0_hit ? _GEN_517 : ram_0_60; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1161 = way0_hit ? _GEN_518 : ram_0_61; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1162 = way0_hit ? _GEN_519 : ram_0_62; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_1163 = way0_hit ? _GEN_520 : ram_0_63; // @[d_cache.scala 107:27 18:24]
  wire  _GEN_1164 = way0_hit ? _GEN_521 : valid_0_0; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1165 = way0_hit ? _GEN_522 : valid_0_1; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1166 = way0_hit ? _GEN_523 : valid_0_2; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1167 = way0_hit ? _GEN_524 : valid_0_3; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1168 = way0_hit ? _GEN_525 : valid_0_4; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1169 = way0_hit ? _GEN_526 : valid_0_5; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1170 = way0_hit ? _GEN_527 : valid_0_6; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1171 = way0_hit ? _GEN_528 : valid_0_7; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1172 = way0_hit ? _GEN_529 : valid_0_8; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1173 = way0_hit ? _GEN_530 : valid_0_9; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1174 = way0_hit ? _GEN_531 : valid_0_10; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1175 = way0_hit ? _GEN_532 : valid_0_11; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1176 = way0_hit ? _GEN_533 : valid_0_12; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1177 = way0_hit ? _GEN_534 : valid_0_13; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1178 = way0_hit ? _GEN_535 : valid_0_14; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1179 = way0_hit ? _GEN_536 : valid_0_15; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1180 = way0_hit ? _GEN_537 : valid_0_16; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1181 = way0_hit ? _GEN_538 : valid_0_17; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1182 = way0_hit ? _GEN_539 : valid_0_18; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1183 = way0_hit ? _GEN_540 : valid_0_19; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1184 = way0_hit ? _GEN_541 : valid_0_20; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1185 = way0_hit ? _GEN_542 : valid_0_21; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1186 = way0_hit ? _GEN_543 : valid_0_22; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1187 = way0_hit ? _GEN_544 : valid_0_23; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1188 = way0_hit ? _GEN_545 : valid_0_24; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1189 = way0_hit ? _GEN_546 : valid_0_25; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1190 = way0_hit ? _GEN_547 : valid_0_26; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1191 = way0_hit ? _GEN_548 : valid_0_27; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1192 = way0_hit ? _GEN_549 : valid_0_28; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1193 = way0_hit ? _GEN_550 : valid_0_29; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1194 = way0_hit ? _GEN_551 : valid_0_30; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1195 = way0_hit ? _GEN_552 : valid_0_31; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1196 = way0_hit ? _GEN_553 : valid_0_32; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1197 = way0_hit ? _GEN_554 : valid_0_33; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1198 = way0_hit ? _GEN_555 : valid_0_34; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1199 = way0_hit ? _GEN_556 : valid_0_35; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1200 = way0_hit ? _GEN_557 : valid_0_36; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1201 = way0_hit ? _GEN_558 : valid_0_37; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1202 = way0_hit ? _GEN_559 : valid_0_38; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1203 = way0_hit ? _GEN_560 : valid_0_39; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1204 = way0_hit ? _GEN_561 : valid_0_40; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1205 = way0_hit ? _GEN_562 : valid_0_41; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1206 = way0_hit ? _GEN_563 : valid_0_42; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1207 = way0_hit ? _GEN_564 : valid_0_43; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1208 = way0_hit ? _GEN_565 : valid_0_44; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1209 = way0_hit ? _GEN_566 : valid_0_45; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1210 = way0_hit ? _GEN_567 : valid_0_46; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1211 = way0_hit ? _GEN_568 : valid_0_47; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1212 = way0_hit ? _GEN_569 : valid_0_48; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1213 = way0_hit ? _GEN_570 : valid_0_49; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1214 = way0_hit ? _GEN_571 : valid_0_50; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1215 = way0_hit ? _GEN_572 : valid_0_51; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1216 = way0_hit ? _GEN_573 : valid_0_52; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1217 = way0_hit ? _GEN_574 : valid_0_53; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1218 = way0_hit ? _GEN_575 : valid_0_54; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1219 = way0_hit ? _GEN_576 : valid_0_55; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1220 = way0_hit ? _GEN_577 : valid_0_56; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1221 = way0_hit ? _GEN_578 : valid_0_57; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1222 = way0_hit ? _GEN_579 : valid_0_58; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1223 = way0_hit ? _GEN_580 : valid_0_59; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1224 = way0_hit ? _GEN_581 : valid_0_60; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1225 = way0_hit ? _GEN_582 : valid_0_61; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1226 = way0_hit ? _GEN_583 : valid_0_62; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1227 = way0_hit ? _GEN_584 : valid_0_63; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_1228 = way0_hit ? _GEN_585 : dirty_0_0; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1229 = way0_hit ? _GEN_586 : dirty_0_1; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1230 = way0_hit ? _GEN_587 : dirty_0_2; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1231 = way0_hit ? _GEN_588 : dirty_0_3; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1232 = way0_hit ? _GEN_589 : dirty_0_4; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1233 = way0_hit ? _GEN_590 : dirty_0_5; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1234 = way0_hit ? _GEN_591 : dirty_0_6; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1235 = way0_hit ? _GEN_592 : dirty_0_7; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1236 = way0_hit ? _GEN_593 : dirty_0_8; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1237 = way0_hit ? _GEN_594 : dirty_0_9; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1238 = way0_hit ? _GEN_595 : dirty_0_10; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1239 = way0_hit ? _GEN_596 : dirty_0_11; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1240 = way0_hit ? _GEN_597 : dirty_0_12; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1241 = way0_hit ? _GEN_598 : dirty_0_13; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1242 = way0_hit ? _GEN_599 : dirty_0_14; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1243 = way0_hit ? _GEN_600 : dirty_0_15; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1244 = way0_hit ? _GEN_601 : dirty_0_16; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1245 = way0_hit ? _GEN_602 : dirty_0_17; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1246 = way0_hit ? _GEN_603 : dirty_0_18; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1247 = way0_hit ? _GEN_604 : dirty_0_19; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1248 = way0_hit ? _GEN_605 : dirty_0_20; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1249 = way0_hit ? _GEN_606 : dirty_0_21; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1250 = way0_hit ? _GEN_607 : dirty_0_22; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1251 = way0_hit ? _GEN_608 : dirty_0_23; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1252 = way0_hit ? _GEN_609 : dirty_0_24; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1253 = way0_hit ? _GEN_610 : dirty_0_25; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1254 = way0_hit ? _GEN_611 : dirty_0_26; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1255 = way0_hit ? _GEN_612 : dirty_0_27; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1256 = way0_hit ? _GEN_613 : dirty_0_28; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1257 = way0_hit ? _GEN_614 : dirty_0_29; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1258 = way0_hit ? _GEN_615 : dirty_0_30; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1259 = way0_hit ? _GEN_616 : dirty_0_31; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1260 = way0_hit ? _GEN_617 : dirty_0_32; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1261 = way0_hit ? _GEN_618 : dirty_0_33; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1262 = way0_hit ? _GEN_619 : dirty_0_34; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1263 = way0_hit ? _GEN_620 : dirty_0_35; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1264 = way0_hit ? _GEN_621 : dirty_0_36; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1265 = way0_hit ? _GEN_622 : dirty_0_37; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1266 = way0_hit ? _GEN_623 : dirty_0_38; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1267 = way0_hit ? _GEN_624 : dirty_0_39; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1268 = way0_hit ? _GEN_625 : dirty_0_40; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1269 = way0_hit ? _GEN_626 : dirty_0_41; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1270 = way0_hit ? _GEN_627 : dirty_0_42; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1271 = way0_hit ? _GEN_628 : dirty_0_43; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1272 = way0_hit ? _GEN_629 : dirty_0_44; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1273 = way0_hit ? _GEN_630 : dirty_0_45; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1274 = way0_hit ? _GEN_631 : dirty_0_46; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1275 = way0_hit ? _GEN_632 : dirty_0_47; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1276 = way0_hit ? _GEN_633 : dirty_0_48; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1277 = way0_hit ? _GEN_634 : dirty_0_49; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1278 = way0_hit ? _GEN_635 : dirty_0_50; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1279 = way0_hit ? _GEN_636 : dirty_0_51; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1280 = way0_hit ? _GEN_637 : dirty_0_52; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1281 = way0_hit ? _GEN_638 : dirty_0_53; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1282 = way0_hit ? _GEN_639 : dirty_0_54; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1283 = way0_hit ? _GEN_640 : dirty_0_55; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1284 = way0_hit ? _GEN_641 : dirty_0_56; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1285 = way0_hit ? _GEN_642 : dirty_0_57; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1286 = way0_hit ? _GEN_643 : dirty_0_58; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1287 = way0_hit ? _GEN_644 : dirty_0_59; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1288 = way0_hit ? _GEN_645 : dirty_0_60; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1289 = way0_hit ? _GEN_646 : dirty_0_61; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1290 = way0_hit ? _GEN_647 : dirty_0_62; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1291 = way0_hit ? _GEN_648 : dirty_0_63; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_1292 = way0_hit | _GEN_1098; // @[d_cache.scala 107:27 115:23]
  wire [63:0] _GEN_1293 = way0_hit ? ram_1_0 : _GEN_906; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1294 = way0_hit ? ram_1_1 : _GEN_907; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1295 = way0_hit ? ram_1_2 : _GEN_908; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1296 = way0_hit ? ram_1_3 : _GEN_909; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1297 = way0_hit ? ram_1_4 : _GEN_910; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1298 = way0_hit ? ram_1_5 : _GEN_911; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1299 = way0_hit ? ram_1_6 : _GEN_912; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1300 = way0_hit ? ram_1_7 : _GEN_913; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1301 = way0_hit ? ram_1_8 : _GEN_914; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1302 = way0_hit ? ram_1_9 : _GEN_915; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1303 = way0_hit ? ram_1_10 : _GEN_916; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1304 = way0_hit ? ram_1_11 : _GEN_917; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1305 = way0_hit ? ram_1_12 : _GEN_918; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1306 = way0_hit ? ram_1_13 : _GEN_919; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1307 = way0_hit ? ram_1_14 : _GEN_920; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1308 = way0_hit ? ram_1_15 : _GEN_921; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1309 = way0_hit ? ram_1_16 : _GEN_922; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1310 = way0_hit ? ram_1_17 : _GEN_923; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1311 = way0_hit ? ram_1_18 : _GEN_924; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1312 = way0_hit ? ram_1_19 : _GEN_925; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1313 = way0_hit ? ram_1_20 : _GEN_926; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1314 = way0_hit ? ram_1_21 : _GEN_927; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1315 = way0_hit ? ram_1_22 : _GEN_928; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1316 = way0_hit ? ram_1_23 : _GEN_929; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1317 = way0_hit ? ram_1_24 : _GEN_930; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1318 = way0_hit ? ram_1_25 : _GEN_931; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1319 = way0_hit ? ram_1_26 : _GEN_932; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1320 = way0_hit ? ram_1_27 : _GEN_933; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1321 = way0_hit ? ram_1_28 : _GEN_934; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1322 = way0_hit ? ram_1_29 : _GEN_935; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1323 = way0_hit ? ram_1_30 : _GEN_936; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1324 = way0_hit ? ram_1_31 : _GEN_937; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1325 = way0_hit ? ram_1_32 : _GEN_938; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1326 = way0_hit ? ram_1_33 : _GEN_939; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1327 = way0_hit ? ram_1_34 : _GEN_940; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1328 = way0_hit ? ram_1_35 : _GEN_941; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1329 = way0_hit ? ram_1_36 : _GEN_942; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1330 = way0_hit ? ram_1_37 : _GEN_943; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1331 = way0_hit ? ram_1_38 : _GEN_944; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1332 = way0_hit ? ram_1_39 : _GEN_945; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1333 = way0_hit ? ram_1_40 : _GEN_946; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1334 = way0_hit ? ram_1_41 : _GEN_947; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1335 = way0_hit ? ram_1_42 : _GEN_948; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1336 = way0_hit ? ram_1_43 : _GEN_949; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1337 = way0_hit ? ram_1_44 : _GEN_950; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1338 = way0_hit ? ram_1_45 : _GEN_951; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1339 = way0_hit ? ram_1_46 : _GEN_952; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1340 = way0_hit ? ram_1_47 : _GEN_953; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1341 = way0_hit ? ram_1_48 : _GEN_954; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1342 = way0_hit ? ram_1_49 : _GEN_955; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1343 = way0_hit ? ram_1_50 : _GEN_956; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1344 = way0_hit ? ram_1_51 : _GEN_957; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1345 = way0_hit ? ram_1_52 : _GEN_958; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1346 = way0_hit ? ram_1_53 : _GEN_959; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1347 = way0_hit ? ram_1_54 : _GEN_960; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1348 = way0_hit ? ram_1_55 : _GEN_961; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1349 = way0_hit ? ram_1_56 : _GEN_962; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1350 = way0_hit ? ram_1_57 : _GEN_963; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1351 = way0_hit ? ram_1_58 : _GEN_964; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1352 = way0_hit ? ram_1_59 : _GEN_965; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1353 = way0_hit ? ram_1_60 : _GEN_966; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1354 = way0_hit ? ram_1_61 : _GEN_967; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1355 = way0_hit ? ram_1_62 : _GEN_968; // @[d_cache.scala 107:27 19:24]
  wire [63:0] _GEN_1356 = way0_hit ? ram_1_63 : _GEN_969; // @[d_cache.scala 107:27 19:24]
  wire  _GEN_1357 = way0_hit ? valid_1_0 : _GEN_970; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1358 = way0_hit ? valid_1_1 : _GEN_971; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1359 = way0_hit ? valid_1_2 : _GEN_972; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1360 = way0_hit ? valid_1_3 : _GEN_973; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1361 = way0_hit ? valid_1_4 : _GEN_974; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1362 = way0_hit ? valid_1_5 : _GEN_975; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1363 = way0_hit ? valid_1_6 : _GEN_976; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1364 = way0_hit ? valid_1_7 : _GEN_977; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1365 = way0_hit ? valid_1_8 : _GEN_978; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1366 = way0_hit ? valid_1_9 : _GEN_979; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1367 = way0_hit ? valid_1_10 : _GEN_980; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1368 = way0_hit ? valid_1_11 : _GEN_981; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1369 = way0_hit ? valid_1_12 : _GEN_982; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1370 = way0_hit ? valid_1_13 : _GEN_983; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1371 = way0_hit ? valid_1_14 : _GEN_984; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1372 = way0_hit ? valid_1_15 : _GEN_985; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1373 = way0_hit ? valid_1_16 : _GEN_986; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1374 = way0_hit ? valid_1_17 : _GEN_987; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1375 = way0_hit ? valid_1_18 : _GEN_988; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1376 = way0_hit ? valid_1_19 : _GEN_989; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1377 = way0_hit ? valid_1_20 : _GEN_990; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1378 = way0_hit ? valid_1_21 : _GEN_991; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1379 = way0_hit ? valid_1_22 : _GEN_992; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1380 = way0_hit ? valid_1_23 : _GEN_993; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1381 = way0_hit ? valid_1_24 : _GEN_994; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1382 = way0_hit ? valid_1_25 : _GEN_995; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1383 = way0_hit ? valid_1_26 : _GEN_996; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1384 = way0_hit ? valid_1_27 : _GEN_997; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1385 = way0_hit ? valid_1_28 : _GEN_998; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1386 = way0_hit ? valid_1_29 : _GEN_999; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1387 = way0_hit ? valid_1_30 : _GEN_1000; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1388 = way0_hit ? valid_1_31 : _GEN_1001; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1389 = way0_hit ? valid_1_32 : _GEN_1002; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1390 = way0_hit ? valid_1_33 : _GEN_1003; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1391 = way0_hit ? valid_1_34 : _GEN_1004; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1392 = way0_hit ? valid_1_35 : _GEN_1005; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1393 = way0_hit ? valid_1_36 : _GEN_1006; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1394 = way0_hit ? valid_1_37 : _GEN_1007; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1395 = way0_hit ? valid_1_38 : _GEN_1008; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1396 = way0_hit ? valid_1_39 : _GEN_1009; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1397 = way0_hit ? valid_1_40 : _GEN_1010; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1398 = way0_hit ? valid_1_41 : _GEN_1011; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1399 = way0_hit ? valid_1_42 : _GEN_1012; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1400 = way0_hit ? valid_1_43 : _GEN_1013; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1401 = way0_hit ? valid_1_44 : _GEN_1014; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1402 = way0_hit ? valid_1_45 : _GEN_1015; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1403 = way0_hit ? valid_1_46 : _GEN_1016; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1404 = way0_hit ? valid_1_47 : _GEN_1017; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1405 = way0_hit ? valid_1_48 : _GEN_1018; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1406 = way0_hit ? valid_1_49 : _GEN_1019; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1407 = way0_hit ? valid_1_50 : _GEN_1020; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1408 = way0_hit ? valid_1_51 : _GEN_1021; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1409 = way0_hit ? valid_1_52 : _GEN_1022; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1410 = way0_hit ? valid_1_53 : _GEN_1023; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1411 = way0_hit ? valid_1_54 : _GEN_1024; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1412 = way0_hit ? valid_1_55 : _GEN_1025; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1413 = way0_hit ? valid_1_56 : _GEN_1026; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1414 = way0_hit ? valid_1_57 : _GEN_1027; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1415 = way0_hit ? valid_1_58 : _GEN_1028; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1416 = way0_hit ? valid_1_59 : _GEN_1029; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1417 = way0_hit ? valid_1_60 : _GEN_1030; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1418 = way0_hit ? valid_1_61 : _GEN_1031; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1419 = way0_hit ? valid_1_62 : _GEN_1032; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1420 = way0_hit ? valid_1_63 : _GEN_1033; // @[d_cache.scala 107:27 25:26]
  wire  _GEN_1421 = way0_hit ? dirty_1_0 : _GEN_1034; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1422 = way0_hit ? dirty_1_1 : _GEN_1035; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1423 = way0_hit ? dirty_1_2 : _GEN_1036; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1424 = way0_hit ? dirty_1_3 : _GEN_1037; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1425 = way0_hit ? dirty_1_4 : _GEN_1038; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1426 = way0_hit ? dirty_1_5 : _GEN_1039; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1427 = way0_hit ? dirty_1_6 : _GEN_1040; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1428 = way0_hit ? dirty_1_7 : _GEN_1041; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1429 = way0_hit ? dirty_1_8 : _GEN_1042; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1430 = way0_hit ? dirty_1_9 : _GEN_1043; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1431 = way0_hit ? dirty_1_10 : _GEN_1044; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1432 = way0_hit ? dirty_1_11 : _GEN_1045; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1433 = way0_hit ? dirty_1_12 : _GEN_1046; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1434 = way0_hit ? dirty_1_13 : _GEN_1047; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1435 = way0_hit ? dirty_1_14 : _GEN_1048; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1436 = way0_hit ? dirty_1_15 : _GEN_1049; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1437 = way0_hit ? dirty_1_16 : _GEN_1050; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1438 = way0_hit ? dirty_1_17 : _GEN_1051; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1439 = way0_hit ? dirty_1_18 : _GEN_1052; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1440 = way0_hit ? dirty_1_19 : _GEN_1053; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1441 = way0_hit ? dirty_1_20 : _GEN_1054; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1442 = way0_hit ? dirty_1_21 : _GEN_1055; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1443 = way0_hit ? dirty_1_22 : _GEN_1056; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1444 = way0_hit ? dirty_1_23 : _GEN_1057; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1445 = way0_hit ? dirty_1_24 : _GEN_1058; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1446 = way0_hit ? dirty_1_25 : _GEN_1059; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1447 = way0_hit ? dirty_1_26 : _GEN_1060; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1448 = way0_hit ? dirty_1_27 : _GEN_1061; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1449 = way0_hit ? dirty_1_28 : _GEN_1062; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1450 = way0_hit ? dirty_1_29 : _GEN_1063; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1451 = way0_hit ? dirty_1_30 : _GEN_1064; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1452 = way0_hit ? dirty_1_31 : _GEN_1065; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1453 = way0_hit ? dirty_1_32 : _GEN_1066; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1454 = way0_hit ? dirty_1_33 : _GEN_1067; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1455 = way0_hit ? dirty_1_34 : _GEN_1068; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1456 = way0_hit ? dirty_1_35 : _GEN_1069; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1457 = way0_hit ? dirty_1_36 : _GEN_1070; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1458 = way0_hit ? dirty_1_37 : _GEN_1071; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1459 = way0_hit ? dirty_1_38 : _GEN_1072; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1460 = way0_hit ? dirty_1_39 : _GEN_1073; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1461 = way0_hit ? dirty_1_40 : _GEN_1074; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1462 = way0_hit ? dirty_1_41 : _GEN_1075; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1463 = way0_hit ? dirty_1_42 : _GEN_1076; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1464 = way0_hit ? dirty_1_43 : _GEN_1077; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1465 = way0_hit ? dirty_1_44 : _GEN_1078; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1466 = way0_hit ? dirty_1_45 : _GEN_1079; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1467 = way0_hit ? dirty_1_46 : _GEN_1080; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1468 = way0_hit ? dirty_1_47 : _GEN_1081; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1469 = way0_hit ? dirty_1_48 : _GEN_1082; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1470 = way0_hit ? dirty_1_49 : _GEN_1083; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1471 = way0_hit ? dirty_1_50 : _GEN_1084; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1472 = way0_hit ? dirty_1_51 : _GEN_1085; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1473 = way0_hit ? dirty_1_52 : _GEN_1086; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1474 = way0_hit ? dirty_1_53 : _GEN_1087; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1475 = way0_hit ? dirty_1_54 : _GEN_1088; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1476 = way0_hit ? dirty_1_55 : _GEN_1089; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1477 = way0_hit ? dirty_1_56 : _GEN_1090; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1478 = way0_hit ? dirty_1_57 : _GEN_1091; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1479 = way0_hit ? dirty_1_58 : _GEN_1092; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1480 = way0_hit ? dirty_1_59 : _GEN_1093; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1481 = way0_hit ? dirty_1_60 : _GEN_1094; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1482 = way0_hit ? dirty_1_61 : _GEN_1095; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1483 = way0_hit ? dirty_1_62 : _GEN_1096; // @[d_cache.scala 107:27 27:26]
  wire  _GEN_1484 = way0_hit ? dirty_1_63 : _GEN_1097; // @[d_cache.scala 107:27 27:26]
  wire [2:0] _GEN_1485 = io_from_axi_rvalid ? 3'h5 : state; // @[d_cache.scala 128:37 129:23 76:24]
  wire [63:0] _GEN_1486 = io_from_axi_rvalid ? io_from_axi_rdata : receive_data; // @[d_cache.scala 131:37 132:30 36:31]
  wire [2:0] _GEN_1487 = io_from_axi_bvalid ? 3'h0 : state; // @[d_cache.scala 136:37 137:23 76:24]
  wire [63:0] _GEN_1488 = 6'h0 == index ? receive_data : ram_0_0; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1489 = 6'h1 == index ? receive_data : ram_0_1; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1490 = 6'h2 == index ? receive_data : ram_0_2; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1491 = 6'h3 == index ? receive_data : ram_0_3; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1492 = 6'h4 == index ? receive_data : ram_0_4; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1493 = 6'h5 == index ? receive_data : ram_0_5; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1494 = 6'h6 == index ? receive_data : ram_0_6; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1495 = 6'h7 == index ? receive_data : ram_0_7; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1496 = 6'h8 == index ? receive_data : ram_0_8; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1497 = 6'h9 == index ? receive_data : ram_0_9; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1498 = 6'ha == index ? receive_data : ram_0_10; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1499 = 6'hb == index ? receive_data : ram_0_11; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1500 = 6'hc == index ? receive_data : ram_0_12; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1501 = 6'hd == index ? receive_data : ram_0_13; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1502 = 6'he == index ? receive_data : ram_0_14; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1503 = 6'hf == index ? receive_data : ram_0_15; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1504 = 6'h10 == index ? receive_data : ram_0_16; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1505 = 6'h11 == index ? receive_data : ram_0_17; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1506 = 6'h12 == index ? receive_data : ram_0_18; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1507 = 6'h13 == index ? receive_data : ram_0_19; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1508 = 6'h14 == index ? receive_data : ram_0_20; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1509 = 6'h15 == index ? receive_data : ram_0_21; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1510 = 6'h16 == index ? receive_data : ram_0_22; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1511 = 6'h17 == index ? receive_data : ram_0_23; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1512 = 6'h18 == index ? receive_data : ram_0_24; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1513 = 6'h19 == index ? receive_data : ram_0_25; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1514 = 6'h1a == index ? receive_data : ram_0_26; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1515 = 6'h1b == index ? receive_data : ram_0_27; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1516 = 6'h1c == index ? receive_data : ram_0_28; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1517 = 6'h1d == index ? receive_data : ram_0_29; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1518 = 6'h1e == index ? receive_data : ram_0_30; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1519 = 6'h1f == index ? receive_data : ram_0_31; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1520 = 6'h20 == index ? receive_data : ram_0_32; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1521 = 6'h21 == index ? receive_data : ram_0_33; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1522 = 6'h22 == index ? receive_data : ram_0_34; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1523 = 6'h23 == index ? receive_data : ram_0_35; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1524 = 6'h24 == index ? receive_data : ram_0_36; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1525 = 6'h25 == index ? receive_data : ram_0_37; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1526 = 6'h26 == index ? receive_data : ram_0_38; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1527 = 6'h27 == index ? receive_data : ram_0_39; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1528 = 6'h28 == index ? receive_data : ram_0_40; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1529 = 6'h29 == index ? receive_data : ram_0_41; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1530 = 6'h2a == index ? receive_data : ram_0_42; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1531 = 6'h2b == index ? receive_data : ram_0_43; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1532 = 6'h2c == index ? receive_data : ram_0_44; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1533 = 6'h2d == index ? receive_data : ram_0_45; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1534 = 6'h2e == index ? receive_data : ram_0_46; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1535 = 6'h2f == index ? receive_data : ram_0_47; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1536 = 6'h30 == index ? receive_data : ram_0_48; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1537 = 6'h31 == index ? receive_data : ram_0_49; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1538 = 6'h32 == index ? receive_data : ram_0_50; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1539 = 6'h33 == index ? receive_data : ram_0_51; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1540 = 6'h34 == index ? receive_data : ram_0_52; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1541 = 6'h35 == index ? receive_data : ram_0_53; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1542 = 6'h36 == index ? receive_data : ram_0_54; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1543 = 6'h37 == index ? receive_data : ram_0_55; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1544 = 6'h38 == index ? receive_data : ram_0_56; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1545 = 6'h39 == index ? receive_data : ram_0_57; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1546 = 6'h3a == index ? receive_data : ram_0_58; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1547 = 6'h3b == index ? receive_data : ram_0_59; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1548 = 6'h3c == index ? receive_data : ram_0_60; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1549 = 6'h3d == index ? receive_data : ram_0_61; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1550 = 6'h3e == index ? receive_data : ram_0_62; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_1551 = 6'h3f == index ? receive_data : ram_0_63; // @[d_cache.scala 143:{30,30} 18:24]
  wire [31:0] _GEN_1552 = 6'h0 == index ? _GEN_8027 : tag_0_0; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1553 = 6'h1 == index ? _GEN_8027 : tag_0_1; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1554 = 6'h2 == index ? _GEN_8027 : tag_0_2; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1555 = 6'h3 == index ? _GEN_8027 : tag_0_3; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1556 = 6'h4 == index ? _GEN_8027 : tag_0_4; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1557 = 6'h5 == index ? _GEN_8027 : tag_0_5; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1558 = 6'h6 == index ? _GEN_8027 : tag_0_6; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1559 = 6'h7 == index ? _GEN_8027 : tag_0_7; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1560 = 6'h8 == index ? _GEN_8027 : tag_0_8; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1561 = 6'h9 == index ? _GEN_8027 : tag_0_9; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1562 = 6'ha == index ? _GEN_8027 : tag_0_10; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1563 = 6'hb == index ? _GEN_8027 : tag_0_11; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1564 = 6'hc == index ? _GEN_8027 : tag_0_12; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1565 = 6'hd == index ? _GEN_8027 : tag_0_13; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1566 = 6'he == index ? _GEN_8027 : tag_0_14; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1567 = 6'hf == index ? _GEN_8027 : tag_0_15; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1568 = 6'h10 == index ? _GEN_8027 : tag_0_16; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1569 = 6'h11 == index ? _GEN_8027 : tag_0_17; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1570 = 6'h12 == index ? _GEN_8027 : tag_0_18; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1571 = 6'h13 == index ? _GEN_8027 : tag_0_19; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1572 = 6'h14 == index ? _GEN_8027 : tag_0_20; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1573 = 6'h15 == index ? _GEN_8027 : tag_0_21; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1574 = 6'h16 == index ? _GEN_8027 : tag_0_22; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1575 = 6'h17 == index ? _GEN_8027 : tag_0_23; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1576 = 6'h18 == index ? _GEN_8027 : tag_0_24; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1577 = 6'h19 == index ? _GEN_8027 : tag_0_25; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1578 = 6'h1a == index ? _GEN_8027 : tag_0_26; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1579 = 6'h1b == index ? _GEN_8027 : tag_0_27; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1580 = 6'h1c == index ? _GEN_8027 : tag_0_28; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1581 = 6'h1d == index ? _GEN_8027 : tag_0_29; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1582 = 6'h1e == index ? _GEN_8027 : tag_0_30; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1583 = 6'h1f == index ? _GEN_8027 : tag_0_31; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1584 = 6'h20 == index ? _GEN_8027 : tag_0_32; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1585 = 6'h21 == index ? _GEN_8027 : tag_0_33; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1586 = 6'h22 == index ? _GEN_8027 : tag_0_34; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1587 = 6'h23 == index ? _GEN_8027 : tag_0_35; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1588 = 6'h24 == index ? _GEN_8027 : tag_0_36; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1589 = 6'h25 == index ? _GEN_8027 : tag_0_37; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1590 = 6'h26 == index ? _GEN_8027 : tag_0_38; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1591 = 6'h27 == index ? _GEN_8027 : tag_0_39; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1592 = 6'h28 == index ? _GEN_8027 : tag_0_40; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1593 = 6'h29 == index ? _GEN_8027 : tag_0_41; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1594 = 6'h2a == index ? _GEN_8027 : tag_0_42; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1595 = 6'h2b == index ? _GEN_8027 : tag_0_43; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1596 = 6'h2c == index ? _GEN_8027 : tag_0_44; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1597 = 6'h2d == index ? _GEN_8027 : tag_0_45; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1598 = 6'h2e == index ? _GEN_8027 : tag_0_46; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1599 = 6'h2f == index ? _GEN_8027 : tag_0_47; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1600 = 6'h30 == index ? _GEN_8027 : tag_0_48; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1601 = 6'h31 == index ? _GEN_8027 : tag_0_49; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1602 = 6'h32 == index ? _GEN_8027 : tag_0_50; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1603 = 6'h33 == index ? _GEN_8027 : tag_0_51; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1604 = 6'h34 == index ? _GEN_8027 : tag_0_52; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1605 = 6'h35 == index ? _GEN_8027 : tag_0_53; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1606 = 6'h36 == index ? _GEN_8027 : tag_0_54; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1607 = 6'h37 == index ? _GEN_8027 : tag_0_55; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1608 = 6'h38 == index ? _GEN_8027 : tag_0_56; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1609 = 6'h39 == index ? _GEN_8027 : tag_0_57; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1610 = 6'h3a == index ? _GEN_8027 : tag_0_58; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1611 = 6'h3b == index ? _GEN_8027 : tag_0_59; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1612 = 6'h3c == index ? _GEN_8027 : tag_0_60; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1613 = 6'h3d == index ? _GEN_8027 : tag_0_61; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1614 = 6'h3e == index ? _GEN_8027 : tag_0_62; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_1615 = 6'h3f == index ? _GEN_8027 : tag_0_63; // @[d_cache.scala 144:{30,30} 22:24]
  wire [63:0] _GEN_1680 = 6'h0 == index ? receive_data : ram_1_0; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1681 = 6'h1 == index ? receive_data : ram_1_1; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1682 = 6'h2 == index ? receive_data : ram_1_2; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1683 = 6'h3 == index ? receive_data : ram_1_3; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1684 = 6'h4 == index ? receive_data : ram_1_4; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1685 = 6'h5 == index ? receive_data : ram_1_5; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1686 = 6'h6 == index ? receive_data : ram_1_6; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1687 = 6'h7 == index ? receive_data : ram_1_7; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1688 = 6'h8 == index ? receive_data : ram_1_8; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1689 = 6'h9 == index ? receive_data : ram_1_9; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1690 = 6'ha == index ? receive_data : ram_1_10; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1691 = 6'hb == index ? receive_data : ram_1_11; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1692 = 6'hc == index ? receive_data : ram_1_12; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1693 = 6'hd == index ? receive_data : ram_1_13; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1694 = 6'he == index ? receive_data : ram_1_14; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1695 = 6'hf == index ? receive_data : ram_1_15; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1696 = 6'h10 == index ? receive_data : ram_1_16; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1697 = 6'h11 == index ? receive_data : ram_1_17; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1698 = 6'h12 == index ? receive_data : ram_1_18; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1699 = 6'h13 == index ? receive_data : ram_1_19; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1700 = 6'h14 == index ? receive_data : ram_1_20; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1701 = 6'h15 == index ? receive_data : ram_1_21; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1702 = 6'h16 == index ? receive_data : ram_1_22; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1703 = 6'h17 == index ? receive_data : ram_1_23; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1704 = 6'h18 == index ? receive_data : ram_1_24; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1705 = 6'h19 == index ? receive_data : ram_1_25; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1706 = 6'h1a == index ? receive_data : ram_1_26; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1707 = 6'h1b == index ? receive_data : ram_1_27; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1708 = 6'h1c == index ? receive_data : ram_1_28; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1709 = 6'h1d == index ? receive_data : ram_1_29; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1710 = 6'h1e == index ? receive_data : ram_1_30; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1711 = 6'h1f == index ? receive_data : ram_1_31; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1712 = 6'h20 == index ? receive_data : ram_1_32; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1713 = 6'h21 == index ? receive_data : ram_1_33; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1714 = 6'h22 == index ? receive_data : ram_1_34; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1715 = 6'h23 == index ? receive_data : ram_1_35; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1716 = 6'h24 == index ? receive_data : ram_1_36; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1717 = 6'h25 == index ? receive_data : ram_1_37; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1718 = 6'h26 == index ? receive_data : ram_1_38; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1719 = 6'h27 == index ? receive_data : ram_1_39; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1720 = 6'h28 == index ? receive_data : ram_1_40; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1721 = 6'h29 == index ? receive_data : ram_1_41; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1722 = 6'h2a == index ? receive_data : ram_1_42; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1723 = 6'h2b == index ? receive_data : ram_1_43; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1724 = 6'h2c == index ? receive_data : ram_1_44; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1725 = 6'h2d == index ? receive_data : ram_1_45; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1726 = 6'h2e == index ? receive_data : ram_1_46; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1727 = 6'h2f == index ? receive_data : ram_1_47; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1728 = 6'h30 == index ? receive_data : ram_1_48; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1729 = 6'h31 == index ? receive_data : ram_1_49; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1730 = 6'h32 == index ? receive_data : ram_1_50; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1731 = 6'h33 == index ? receive_data : ram_1_51; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1732 = 6'h34 == index ? receive_data : ram_1_52; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1733 = 6'h35 == index ? receive_data : ram_1_53; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1734 = 6'h36 == index ? receive_data : ram_1_54; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1735 = 6'h37 == index ? receive_data : ram_1_55; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1736 = 6'h38 == index ? receive_data : ram_1_56; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1737 = 6'h39 == index ? receive_data : ram_1_57; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1738 = 6'h3a == index ? receive_data : ram_1_58; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1739 = 6'h3b == index ? receive_data : ram_1_59; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1740 = 6'h3c == index ? receive_data : ram_1_60; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1741 = 6'h3d == index ? receive_data : ram_1_61; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1742 = 6'h3e == index ? receive_data : ram_1_62; // @[d_cache.scala 149:{30,30} 19:24]
  wire [63:0] _GEN_1743 = 6'h3f == index ? receive_data : ram_1_63; // @[d_cache.scala 149:{30,30} 19:24]
  wire [31:0] _GEN_1744 = 6'h0 == index ? _GEN_8027 : tag_1_0; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1745 = 6'h1 == index ? _GEN_8027 : tag_1_1; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1746 = 6'h2 == index ? _GEN_8027 : tag_1_2; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1747 = 6'h3 == index ? _GEN_8027 : tag_1_3; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1748 = 6'h4 == index ? _GEN_8027 : tag_1_4; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1749 = 6'h5 == index ? _GEN_8027 : tag_1_5; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1750 = 6'h6 == index ? _GEN_8027 : tag_1_6; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1751 = 6'h7 == index ? _GEN_8027 : tag_1_7; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1752 = 6'h8 == index ? _GEN_8027 : tag_1_8; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1753 = 6'h9 == index ? _GEN_8027 : tag_1_9; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1754 = 6'ha == index ? _GEN_8027 : tag_1_10; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1755 = 6'hb == index ? _GEN_8027 : tag_1_11; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1756 = 6'hc == index ? _GEN_8027 : tag_1_12; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1757 = 6'hd == index ? _GEN_8027 : tag_1_13; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1758 = 6'he == index ? _GEN_8027 : tag_1_14; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1759 = 6'hf == index ? _GEN_8027 : tag_1_15; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1760 = 6'h10 == index ? _GEN_8027 : tag_1_16; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1761 = 6'h11 == index ? _GEN_8027 : tag_1_17; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1762 = 6'h12 == index ? _GEN_8027 : tag_1_18; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1763 = 6'h13 == index ? _GEN_8027 : tag_1_19; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1764 = 6'h14 == index ? _GEN_8027 : tag_1_20; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1765 = 6'h15 == index ? _GEN_8027 : tag_1_21; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1766 = 6'h16 == index ? _GEN_8027 : tag_1_22; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1767 = 6'h17 == index ? _GEN_8027 : tag_1_23; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1768 = 6'h18 == index ? _GEN_8027 : tag_1_24; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1769 = 6'h19 == index ? _GEN_8027 : tag_1_25; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1770 = 6'h1a == index ? _GEN_8027 : tag_1_26; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1771 = 6'h1b == index ? _GEN_8027 : tag_1_27; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1772 = 6'h1c == index ? _GEN_8027 : tag_1_28; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1773 = 6'h1d == index ? _GEN_8027 : tag_1_29; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1774 = 6'h1e == index ? _GEN_8027 : tag_1_30; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1775 = 6'h1f == index ? _GEN_8027 : tag_1_31; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1776 = 6'h20 == index ? _GEN_8027 : tag_1_32; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1777 = 6'h21 == index ? _GEN_8027 : tag_1_33; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1778 = 6'h22 == index ? _GEN_8027 : tag_1_34; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1779 = 6'h23 == index ? _GEN_8027 : tag_1_35; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1780 = 6'h24 == index ? _GEN_8027 : tag_1_36; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1781 = 6'h25 == index ? _GEN_8027 : tag_1_37; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1782 = 6'h26 == index ? _GEN_8027 : tag_1_38; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1783 = 6'h27 == index ? _GEN_8027 : tag_1_39; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1784 = 6'h28 == index ? _GEN_8027 : tag_1_40; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1785 = 6'h29 == index ? _GEN_8027 : tag_1_41; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1786 = 6'h2a == index ? _GEN_8027 : tag_1_42; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1787 = 6'h2b == index ? _GEN_8027 : tag_1_43; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1788 = 6'h2c == index ? _GEN_8027 : tag_1_44; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1789 = 6'h2d == index ? _GEN_8027 : tag_1_45; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1790 = 6'h2e == index ? _GEN_8027 : tag_1_46; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1791 = 6'h2f == index ? _GEN_8027 : tag_1_47; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1792 = 6'h30 == index ? _GEN_8027 : tag_1_48; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1793 = 6'h31 == index ? _GEN_8027 : tag_1_49; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1794 = 6'h32 == index ? _GEN_8027 : tag_1_50; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1795 = 6'h33 == index ? _GEN_8027 : tag_1_51; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1796 = 6'h34 == index ? _GEN_8027 : tag_1_52; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1797 = 6'h35 == index ? _GEN_8027 : tag_1_53; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1798 = 6'h36 == index ? _GEN_8027 : tag_1_54; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1799 = 6'h37 == index ? _GEN_8027 : tag_1_55; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1800 = 6'h38 == index ? _GEN_8027 : tag_1_56; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1801 = 6'h39 == index ? _GEN_8027 : tag_1_57; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1802 = 6'h3a == index ? _GEN_8027 : tag_1_58; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1803 = 6'h3b == index ? _GEN_8027 : tag_1_59; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1804 = 6'h3c == index ? _GEN_8027 : tag_1_60; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1805 = 6'h3d == index ? _GEN_8027 : tag_1_61; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1806 = 6'h3e == index ? _GEN_8027 : tag_1_62; // @[d_cache.scala 150:{30,30} 23:24]
  wire [31:0] _GEN_1807 = 6'h3f == index ? _GEN_8027 : tag_1_63; // @[d_cache.scala 150:{30,30} 23:24]
  wire [40:0] _write_back_addr_T_1 = {_GEN_63,index,3'h0}; // @[Cat.scala 31:58]
  wire  _GEN_2000 = 6'h0 == index ? 1'h0 : dirty_0_0; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2001 = 6'h1 == index ? 1'h0 : dirty_0_1; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2002 = 6'h2 == index ? 1'h0 : dirty_0_2; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2003 = 6'h3 == index ? 1'h0 : dirty_0_3; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2004 = 6'h4 == index ? 1'h0 : dirty_0_4; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2005 = 6'h5 == index ? 1'h0 : dirty_0_5; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2006 = 6'h6 == index ? 1'h0 : dirty_0_6; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2007 = 6'h7 == index ? 1'h0 : dirty_0_7; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2008 = 6'h8 == index ? 1'h0 : dirty_0_8; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2009 = 6'h9 == index ? 1'h0 : dirty_0_9; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2010 = 6'ha == index ? 1'h0 : dirty_0_10; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2011 = 6'hb == index ? 1'h0 : dirty_0_11; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2012 = 6'hc == index ? 1'h0 : dirty_0_12; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2013 = 6'hd == index ? 1'h0 : dirty_0_13; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2014 = 6'he == index ? 1'h0 : dirty_0_14; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2015 = 6'hf == index ? 1'h0 : dirty_0_15; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2016 = 6'h10 == index ? 1'h0 : dirty_0_16; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2017 = 6'h11 == index ? 1'h0 : dirty_0_17; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2018 = 6'h12 == index ? 1'h0 : dirty_0_18; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2019 = 6'h13 == index ? 1'h0 : dirty_0_19; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2020 = 6'h14 == index ? 1'h0 : dirty_0_20; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2021 = 6'h15 == index ? 1'h0 : dirty_0_21; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2022 = 6'h16 == index ? 1'h0 : dirty_0_22; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2023 = 6'h17 == index ? 1'h0 : dirty_0_23; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2024 = 6'h18 == index ? 1'h0 : dirty_0_24; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2025 = 6'h19 == index ? 1'h0 : dirty_0_25; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2026 = 6'h1a == index ? 1'h0 : dirty_0_26; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2027 = 6'h1b == index ? 1'h0 : dirty_0_27; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2028 = 6'h1c == index ? 1'h0 : dirty_0_28; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2029 = 6'h1d == index ? 1'h0 : dirty_0_29; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2030 = 6'h1e == index ? 1'h0 : dirty_0_30; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2031 = 6'h1f == index ? 1'h0 : dirty_0_31; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2032 = 6'h20 == index ? 1'h0 : dirty_0_32; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2033 = 6'h21 == index ? 1'h0 : dirty_0_33; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2034 = 6'h22 == index ? 1'h0 : dirty_0_34; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2035 = 6'h23 == index ? 1'h0 : dirty_0_35; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2036 = 6'h24 == index ? 1'h0 : dirty_0_36; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2037 = 6'h25 == index ? 1'h0 : dirty_0_37; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2038 = 6'h26 == index ? 1'h0 : dirty_0_38; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2039 = 6'h27 == index ? 1'h0 : dirty_0_39; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2040 = 6'h28 == index ? 1'h0 : dirty_0_40; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2041 = 6'h29 == index ? 1'h0 : dirty_0_41; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2042 = 6'h2a == index ? 1'h0 : dirty_0_42; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2043 = 6'h2b == index ? 1'h0 : dirty_0_43; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2044 = 6'h2c == index ? 1'h0 : dirty_0_44; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2045 = 6'h2d == index ? 1'h0 : dirty_0_45; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2046 = 6'h2e == index ? 1'h0 : dirty_0_46; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2047 = 6'h2f == index ? 1'h0 : dirty_0_47; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2048 = 6'h30 == index ? 1'h0 : dirty_0_48; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2049 = 6'h31 == index ? 1'h0 : dirty_0_49; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2050 = 6'h32 == index ? 1'h0 : dirty_0_50; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2051 = 6'h33 == index ? 1'h0 : dirty_0_51; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2052 = 6'h34 == index ? 1'h0 : dirty_0_52; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2053 = 6'h35 == index ? 1'h0 : dirty_0_53; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2054 = 6'h36 == index ? 1'h0 : dirty_0_54; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2055 = 6'h37 == index ? 1'h0 : dirty_0_55; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2056 = 6'h38 == index ? 1'h0 : dirty_0_56; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2057 = 6'h39 == index ? 1'h0 : dirty_0_57; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2058 = 6'h3a == index ? 1'h0 : dirty_0_58; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2059 = 6'h3b == index ? 1'h0 : dirty_0_59; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2060 = 6'h3c == index ? 1'h0 : dirty_0_60; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2061 = 6'h3d == index ? 1'h0 : dirty_0_61; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2062 = 6'h3e == index ? 1'h0 : dirty_0_62; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_2063 = 6'h3f == index ? 1'h0 : dirty_0_63; // @[d_cache.scala 161:{40,40} 26:26]
  wire [63:0] _GEN_2320 = _GEN_325 ? _GEN_456 : write_back_data; // @[d_cache.scala 156:47 157:41 31:34]
  wire [40:0] _GEN_2321 = _GEN_325 ? _write_back_addr_T_1 : {{9'd0}, write_back_addr}; // @[d_cache.scala 156:47 158:41 32:34]
  wire [63:0] _GEN_2322 = _GEN_325 ? _GEN_1488 : _GEN_1488; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2323 = _GEN_325 ? _GEN_1489 : _GEN_1489; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2324 = _GEN_325 ? _GEN_1490 : _GEN_1490; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2325 = _GEN_325 ? _GEN_1491 : _GEN_1491; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2326 = _GEN_325 ? _GEN_1492 : _GEN_1492; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2327 = _GEN_325 ? _GEN_1493 : _GEN_1493; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2328 = _GEN_325 ? _GEN_1494 : _GEN_1494; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2329 = _GEN_325 ? _GEN_1495 : _GEN_1495; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2330 = _GEN_325 ? _GEN_1496 : _GEN_1496; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2331 = _GEN_325 ? _GEN_1497 : _GEN_1497; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2332 = _GEN_325 ? _GEN_1498 : _GEN_1498; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2333 = _GEN_325 ? _GEN_1499 : _GEN_1499; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2334 = _GEN_325 ? _GEN_1500 : _GEN_1500; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2335 = _GEN_325 ? _GEN_1501 : _GEN_1501; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2336 = _GEN_325 ? _GEN_1502 : _GEN_1502; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2337 = _GEN_325 ? _GEN_1503 : _GEN_1503; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2338 = _GEN_325 ? _GEN_1504 : _GEN_1504; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2339 = _GEN_325 ? _GEN_1505 : _GEN_1505; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2340 = _GEN_325 ? _GEN_1506 : _GEN_1506; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2341 = _GEN_325 ? _GEN_1507 : _GEN_1507; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2342 = _GEN_325 ? _GEN_1508 : _GEN_1508; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2343 = _GEN_325 ? _GEN_1509 : _GEN_1509; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2344 = _GEN_325 ? _GEN_1510 : _GEN_1510; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2345 = _GEN_325 ? _GEN_1511 : _GEN_1511; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2346 = _GEN_325 ? _GEN_1512 : _GEN_1512; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2347 = _GEN_325 ? _GEN_1513 : _GEN_1513; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2348 = _GEN_325 ? _GEN_1514 : _GEN_1514; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2349 = _GEN_325 ? _GEN_1515 : _GEN_1515; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2350 = _GEN_325 ? _GEN_1516 : _GEN_1516; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2351 = _GEN_325 ? _GEN_1517 : _GEN_1517; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2352 = _GEN_325 ? _GEN_1518 : _GEN_1518; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2353 = _GEN_325 ? _GEN_1519 : _GEN_1519; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2354 = _GEN_325 ? _GEN_1520 : _GEN_1520; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2355 = _GEN_325 ? _GEN_1521 : _GEN_1521; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2356 = _GEN_325 ? _GEN_1522 : _GEN_1522; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2357 = _GEN_325 ? _GEN_1523 : _GEN_1523; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2358 = _GEN_325 ? _GEN_1524 : _GEN_1524; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2359 = _GEN_325 ? _GEN_1525 : _GEN_1525; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2360 = _GEN_325 ? _GEN_1526 : _GEN_1526; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2361 = _GEN_325 ? _GEN_1527 : _GEN_1527; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2362 = _GEN_325 ? _GEN_1528 : _GEN_1528; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2363 = _GEN_325 ? _GEN_1529 : _GEN_1529; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2364 = _GEN_325 ? _GEN_1530 : _GEN_1530; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2365 = _GEN_325 ? _GEN_1531 : _GEN_1531; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2366 = _GEN_325 ? _GEN_1532 : _GEN_1532; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2367 = _GEN_325 ? _GEN_1533 : _GEN_1533; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2368 = _GEN_325 ? _GEN_1534 : _GEN_1534; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2369 = _GEN_325 ? _GEN_1535 : _GEN_1535; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2370 = _GEN_325 ? _GEN_1536 : _GEN_1536; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2371 = _GEN_325 ? _GEN_1537 : _GEN_1537; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2372 = _GEN_325 ? _GEN_1538 : _GEN_1538; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2373 = _GEN_325 ? _GEN_1539 : _GEN_1539; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2374 = _GEN_325 ? _GEN_1540 : _GEN_1540; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2375 = _GEN_325 ? _GEN_1541 : _GEN_1541; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2376 = _GEN_325 ? _GEN_1542 : _GEN_1542; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2377 = _GEN_325 ? _GEN_1543 : _GEN_1543; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2378 = _GEN_325 ? _GEN_1544 : _GEN_1544; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2379 = _GEN_325 ? _GEN_1545 : _GEN_1545; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2380 = _GEN_325 ? _GEN_1546 : _GEN_1546; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2381 = _GEN_325 ? _GEN_1547 : _GEN_1547; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2382 = _GEN_325 ? _GEN_1548 : _GEN_1548; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2383 = _GEN_325 ? _GEN_1549 : _GEN_1549; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2384 = _GEN_325 ? _GEN_1550 : _GEN_1550; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_2385 = _GEN_325 ? _GEN_1551 : _GEN_1551; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2386 = _GEN_325 ? _GEN_1552 : _GEN_1552; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2387 = _GEN_325 ? _GEN_1553 : _GEN_1553; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2388 = _GEN_325 ? _GEN_1554 : _GEN_1554; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2389 = _GEN_325 ? _GEN_1555 : _GEN_1555; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2390 = _GEN_325 ? _GEN_1556 : _GEN_1556; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2391 = _GEN_325 ? _GEN_1557 : _GEN_1557; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2392 = _GEN_325 ? _GEN_1558 : _GEN_1558; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2393 = _GEN_325 ? _GEN_1559 : _GEN_1559; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2394 = _GEN_325 ? _GEN_1560 : _GEN_1560; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2395 = _GEN_325 ? _GEN_1561 : _GEN_1561; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2396 = _GEN_325 ? _GEN_1562 : _GEN_1562; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2397 = _GEN_325 ? _GEN_1563 : _GEN_1563; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2398 = _GEN_325 ? _GEN_1564 : _GEN_1564; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2399 = _GEN_325 ? _GEN_1565 : _GEN_1565; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2400 = _GEN_325 ? _GEN_1566 : _GEN_1566; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2401 = _GEN_325 ? _GEN_1567 : _GEN_1567; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2402 = _GEN_325 ? _GEN_1568 : _GEN_1568; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2403 = _GEN_325 ? _GEN_1569 : _GEN_1569; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2404 = _GEN_325 ? _GEN_1570 : _GEN_1570; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2405 = _GEN_325 ? _GEN_1571 : _GEN_1571; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2406 = _GEN_325 ? _GEN_1572 : _GEN_1572; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2407 = _GEN_325 ? _GEN_1573 : _GEN_1573; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2408 = _GEN_325 ? _GEN_1574 : _GEN_1574; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2409 = _GEN_325 ? _GEN_1575 : _GEN_1575; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2410 = _GEN_325 ? _GEN_1576 : _GEN_1576; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2411 = _GEN_325 ? _GEN_1577 : _GEN_1577; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2412 = _GEN_325 ? _GEN_1578 : _GEN_1578; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2413 = _GEN_325 ? _GEN_1579 : _GEN_1579; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2414 = _GEN_325 ? _GEN_1580 : _GEN_1580; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2415 = _GEN_325 ? _GEN_1581 : _GEN_1581; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2416 = _GEN_325 ? _GEN_1582 : _GEN_1582; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2417 = _GEN_325 ? _GEN_1583 : _GEN_1583; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2418 = _GEN_325 ? _GEN_1584 : _GEN_1584; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2419 = _GEN_325 ? _GEN_1585 : _GEN_1585; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2420 = _GEN_325 ? _GEN_1586 : _GEN_1586; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2421 = _GEN_325 ? _GEN_1587 : _GEN_1587; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2422 = _GEN_325 ? _GEN_1588 : _GEN_1588; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2423 = _GEN_325 ? _GEN_1589 : _GEN_1589; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2424 = _GEN_325 ? _GEN_1590 : _GEN_1590; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2425 = _GEN_325 ? _GEN_1591 : _GEN_1591; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2426 = _GEN_325 ? _GEN_1592 : _GEN_1592; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2427 = _GEN_325 ? _GEN_1593 : _GEN_1593; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2428 = _GEN_325 ? _GEN_1594 : _GEN_1594; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2429 = _GEN_325 ? _GEN_1595 : _GEN_1595; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2430 = _GEN_325 ? _GEN_1596 : _GEN_1596; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2431 = _GEN_325 ? _GEN_1597 : _GEN_1597; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2432 = _GEN_325 ? _GEN_1598 : _GEN_1598; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2433 = _GEN_325 ? _GEN_1599 : _GEN_1599; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2434 = _GEN_325 ? _GEN_1600 : _GEN_1600; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2435 = _GEN_325 ? _GEN_1601 : _GEN_1601; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2436 = _GEN_325 ? _GEN_1602 : _GEN_1602; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2437 = _GEN_325 ? _GEN_1603 : _GEN_1603; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2438 = _GEN_325 ? _GEN_1604 : _GEN_1604; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2439 = _GEN_325 ? _GEN_1605 : _GEN_1605; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2440 = _GEN_325 ? _GEN_1606 : _GEN_1606; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2441 = _GEN_325 ? _GEN_1607 : _GEN_1607; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2442 = _GEN_325 ? _GEN_1608 : _GEN_1608; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2443 = _GEN_325 ? _GEN_1609 : _GEN_1609; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2444 = _GEN_325 ? _GEN_1610 : _GEN_1610; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2445 = _GEN_325 ? _GEN_1611 : _GEN_1611; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2446 = _GEN_325 ? _GEN_1612 : _GEN_1612; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2447 = _GEN_325 ? _GEN_1613 : _GEN_1613; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2448 = _GEN_325 ? _GEN_1614 : _GEN_1614; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_2449 = _GEN_325 ? _GEN_1615 : _GEN_1615; // @[d_cache.scala 156:47]
  wire  _GEN_2450 = _GEN_325 ? _GEN_2000 : dirty_0_0; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2451 = _GEN_325 ? _GEN_2001 : dirty_0_1; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2452 = _GEN_325 ? _GEN_2002 : dirty_0_2; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2453 = _GEN_325 ? _GEN_2003 : dirty_0_3; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2454 = _GEN_325 ? _GEN_2004 : dirty_0_4; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2455 = _GEN_325 ? _GEN_2005 : dirty_0_5; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2456 = _GEN_325 ? _GEN_2006 : dirty_0_6; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2457 = _GEN_325 ? _GEN_2007 : dirty_0_7; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2458 = _GEN_325 ? _GEN_2008 : dirty_0_8; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2459 = _GEN_325 ? _GEN_2009 : dirty_0_9; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2460 = _GEN_325 ? _GEN_2010 : dirty_0_10; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2461 = _GEN_325 ? _GEN_2011 : dirty_0_11; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2462 = _GEN_325 ? _GEN_2012 : dirty_0_12; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2463 = _GEN_325 ? _GEN_2013 : dirty_0_13; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2464 = _GEN_325 ? _GEN_2014 : dirty_0_14; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2465 = _GEN_325 ? _GEN_2015 : dirty_0_15; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2466 = _GEN_325 ? _GEN_2016 : dirty_0_16; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2467 = _GEN_325 ? _GEN_2017 : dirty_0_17; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2468 = _GEN_325 ? _GEN_2018 : dirty_0_18; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2469 = _GEN_325 ? _GEN_2019 : dirty_0_19; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2470 = _GEN_325 ? _GEN_2020 : dirty_0_20; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2471 = _GEN_325 ? _GEN_2021 : dirty_0_21; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2472 = _GEN_325 ? _GEN_2022 : dirty_0_22; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2473 = _GEN_325 ? _GEN_2023 : dirty_0_23; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2474 = _GEN_325 ? _GEN_2024 : dirty_0_24; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2475 = _GEN_325 ? _GEN_2025 : dirty_0_25; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2476 = _GEN_325 ? _GEN_2026 : dirty_0_26; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2477 = _GEN_325 ? _GEN_2027 : dirty_0_27; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2478 = _GEN_325 ? _GEN_2028 : dirty_0_28; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2479 = _GEN_325 ? _GEN_2029 : dirty_0_29; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2480 = _GEN_325 ? _GEN_2030 : dirty_0_30; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2481 = _GEN_325 ? _GEN_2031 : dirty_0_31; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2482 = _GEN_325 ? _GEN_2032 : dirty_0_32; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2483 = _GEN_325 ? _GEN_2033 : dirty_0_33; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2484 = _GEN_325 ? _GEN_2034 : dirty_0_34; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2485 = _GEN_325 ? _GEN_2035 : dirty_0_35; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2486 = _GEN_325 ? _GEN_2036 : dirty_0_36; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2487 = _GEN_325 ? _GEN_2037 : dirty_0_37; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2488 = _GEN_325 ? _GEN_2038 : dirty_0_38; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2489 = _GEN_325 ? _GEN_2039 : dirty_0_39; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2490 = _GEN_325 ? _GEN_2040 : dirty_0_40; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2491 = _GEN_325 ? _GEN_2041 : dirty_0_41; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2492 = _GEN_325 ? _GEN_2042 : dirty_0_42; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2493 = _GEN_325 ? _GEN_2043 : dirty_0_43; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2494 = _GEN_325 ? _GEN_2044 : dirty_0_44; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2495 = _GEN_325 ? _GEN_2045 : dirty_0_45; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2496 = _GEN_325 ? _GEN_2046 : dirty_0_46; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2497 = _GEN_325 ? _GEN_2047 : dirty_0_47; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2498 = _GEN_325 ? _GEN_2048 : dirty_0_48; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2499 = _GEN_325 ? _GEN_2049 : dirty_0_49; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2500 = _GEN_325 ? _GEN_2050 : dirty_0_50; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2501 = _GEN_325 ? _GEN_2051 : dirty_0_51; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2502 = _GEN_325 ? _GEN_2052 : dirty_0_52; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2503 = _GEN_325 ? _GEN_2053 : dirty_0_53; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2504 = _GEN_325 ? _GEN_2054 : dirty_0_54; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2505 = _GEN_325 ? _GEN_2055 : dirty_0_55; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2506 = _GEN_325 ? _GEN_2056 : dirty_0_56; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2507 = _GEN_325 ? _GEN_2057 : dirty_0_57; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2508 = _GEN_325 ? _GEN_2058 : dirty_0_58; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2509 = _GEN_325 ? _GEN_2059 : dirty_0_59; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2510 = _GEN_325 ? _GEN_2060 : dirty_0_60; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2511 = _GEN_325 ? _GEN_2061 : dirty_0_61; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2512 = _GEN_325 ? _GEN_2062 : dirty_0_62; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2513 = _GEN_325 ? _GEN_2063 : dirty_0_63; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_2514 = _GEN_325 ? _GEN_521 : _GEN_521; // @[d_cache.scala 156:47]
  wire  _GEN_2515 = _GEN_325 ? _GEN_522 : _GEN_522; // @[d_cache.scala 156:47]
  wire  _GEN_2516 = _GEN_325 ? _GEN_523 : _GEN_523; // @[d_cache.scala 156:47]
  wire  _GEN_2517 = _GEN_325 ? _GEN_524 : _GEN_524; // @[d_cache.scala 156:47]
  wire  _GEN_2518 = _GEN_325 ? _GEN_525 : _GEN_525; // @[d_cache.scala 156:47]
  wire  _GEN_2519 = _GEN_325 ? _GEN_526 : _GEN_526; // @[d_cache.scala 156:47]
  wire  _GEN_2520 = _GEN_325 ? _GEN_527 : _GEN_527; // @[d_cache.scala 156:47]
  wire  _GEN_2521 = _GEN_325 ? _GEN_528 : _GEN_528; // @[d_cache.scala 156:47]
  wire  _GEN_2522 = _GEN_325 ? _GEN_529 : _GEN_529; // @[d_cache.scala 156:47]
  wire  _GEN_2523 = _GEN_325 ? _GEN_530 : _GEN_530; // @[d_cache.scala 156:47]
  wire  _GEN_2524 = _GEN_325 ? _GEN_531 : _GEN_531; // @[d_cache.scala 156:47]
  wire  _GEN_2525 = _GEN_325 ? _GEN_532 : _GEN_532; // @[d_cache.scala 156:47]
  wire  _GEN_2526 = _GEN_325 ? _GEN_533 : _GEN_533; // @[d_cache.scala 156:47]
  wire  _GEN_2527 = _GEN_325 ? _GEN_534 : _GEN_534; // @[d_cache.scala 156:47]
  wire  _GEN_2528 = _GEN_325 ? _GEN_535 : _GEN_535; // @[d_cache.scala 156:47]
  wire  _GEN_2529 = _GEN_325 ? _GEN_536 : _GEN_536; // @[d_cache.scala 156:47]
  wire  _GEN_2530 = _GEN_325 ? _GEN_537 : _GEN_537; // @[d_cache.scala 156:47]
  wire  _GEN_2531 = _GEN_325 ? _GEN_538 : _GEN_538; // @[d_cache.scala 156:47]
  wire  _GEN_2532 = _GEN_325 ? _GEN_539 : _GEN_539; // @[d_cache.scala 156:47]
  wire  _GEN_2533 = _GEN_325 ? _GEN_540 : _GEN_540; // @[d_cache.scala 156:47]
  wire  _GEN_2534 = _GEN_325 ? _GEN_541 : _GEN_541; // @[d_cache.scala 156:47]
  wire  _GEN_2535 = _GEN_325 ? _GEN_542 : _GEN_542; // @[d_cache.scala 156:47]
  wire  _GEN_2536 = _GEN_325 ? _GEN_543 : _GEN_543; // @[d_cache.scala 156:47]
  wire  _GEN_2537 = _GEN_325 ? _GEN_544 : _GEN_544; // @[d_cache.scala 156:47]
  wire  _GEN_2538 = _GEN_325 ? _GEN_545 : _GEN_545; // @[d_cache.scala 156:47]
  wire  _GEN_2539 = _GEN_325 ? _GEN_546 : _GEN_546; // @[d_cache.scala 156:47]
  wire  _GEN_2540 = _GEN_325 ? _GEN_547 : _GEN_547; // @[d_cache.scala 156:47]
  wire  _GEN_2541 = _GEN_325 ? _GEN_548 : _GEN_548; // @[d_cache.scala 156:47]
  wire  _GEN_2542 = _GEN_325 ? _GEN_549 : _GEN_549; // @[d_cache.scala 156:47]
  wire  _GEN_2543 = _GEN_325 ? _GEN_550 : _GEN_550; // @[d_cache.scala 156:47]
  wire  _GEN_2544 = _GEN_325 ? _GEN_551 : _GEN_551; // @[d_cache.scala 156:47]
  wire  _GEN_2545 = _GEN_325 ? _GEN_552 : _GEN_552; // @[d_cache.scala 156:47]
  wire  _GEN_2546 = _GEN_325 ? _GEN_553 : _GEN_553; // @[d_cache.scala 156:47]
  wire  _GEN_2547 = _GEN_325 ? _GEN_554 : _GEN_554; // @[d_cache.scala 156:47]
  wire  _GEN_2548 = _GEN_325 ? _GEN_555 : _GEN_555; // @[d_cache.scala 156:47]
  wire  _GEN_2549 = _GEN_325 ? _GEN_556 : _GEN_556; // @[d_cache.scala 156:47]
  wire  _GEN_2550 = _GEN_325 ? _GEN_557 : _GEN_557; // @[d_cache.scala 156:47]
  wire  _GEN_2551 = _GEN_325 ? _GEN_558 : _GEN_558; // @[d_cache.scala 156:47]
  wire  _GEN_2552 = _GEN_325 ? _GEN_559 : _GEN_559; // @[d_cache.scala 156:47]
  wire  _GEN_2553 = _GEN_325 ? _GEN_560 : _GEN_560; // @[d_cache.scala 156:47]
  wire  _GEN_2554 = _GEN_325 ? _GEN_561 : _GEN_561; // @[d_cache.scala 156:47]
  wire  _GEN_2555 = _GEN_325 ? _GEN_562 : _GEN_562; // @[d_cache.scala 156:47]
  wire  _GEN_2556 = _GEN_325 ? _GEN_563 : _GEN_563; // @[d_cache.scala 156:47]
  wire  _GEN_2557 = _GEN_325 ? _GEN_564 : _GEN_564; // @[d_cache.scala 156:47]
  wire  _GEN_2558 = _GEN_325 ? _GEN_565 : _GEN_565; // @[d_cache.scala 156:47]
  wire  _GEN_2559 = _GEN_325 ? _GEN_566 : _GEN_566; // @[d_cache.scala 156:47]
  wire  _GEN_2560 = _GEN_325 ? _GEN_567 : _GEN_567; // @[d_cache.scala 156:47]
  wire  _GEN_2561 = _GEN_325 ? _GEN_568 : _GEN_568; // @[d_cache.scala 156:47]
  wire  _GEN_2562 = _GEN_325 ? _GEN_569 : _GEN_569; // @[d_cache.scala 156:47]
  wire  _GEN_2563 = _GEN_325 ? _GEN_570 : _GEN_570; // @[d_cache.scala 156:47]
  wire  _GEN_2564 = _GEN_325 ? _GEN_571 : _GEN_571; // @[d_cache.scala 156:47]
  wire  _GEN_2565 = _GEN_325 ? _GEN_572 : _GEN_572; // @[d_cache.scala 156:47]
  wire  _GEN_2566 = _GEN_325 ? _GEN_573 : _GEN_573; // @[d_cache.scala 156:47]
  wire  _GEN_2567 = _GEN_325 ? _GEN_574 : _GEN_574; // @[d_cache.scala 156:47]
  wire  _GEN_2568 = _GEN_325 ? _GEN_575 : _GEN_575; // @[d_cache.scala 156:47]
  wire  _GEN_2569 = _GEN_325 ? _GEN_576 : _GEN_576; // @[d_cache.scala 156:47]
  wire  _GEN_2570 = _GEN_325 ? _GEN_577 : _GEN_577; // @[d_cache.scala 156:47]
  wire  _GEN_2571 = _GEN_325 ? _GEN_578 : _GEN_578; // @[d_cache.scala 156:47]
  wire  _GEN_2572 = _GEN_325 ? _GEN_579 : _GEN_579; // @[d_cache.scala 156:47]
  wire  _GEN_2573 = _GEN_325 ? _GEN_580 : _GEN_580; // @[d_cache.scala 156:47]
  wire  _GEN_2574 = _GEN_325 ? _GEN_581 : _GEN_581; // @[d_cache.scala 156:47]
  wire  _GEN_2575 = _GEN_325 ? _GEN_582 : _GEN_582; // @[d_cache.scala 156:47]
  wire  _GEN_2576 = _GEN_325 ? _GEN_583 : _GEN_583; // @[d_cache.scala 156:47]
  wire  _GEN_2577 = _GEN_325 ? _GEN_584 : _GEN_584; // @[d_cache.scala 156:47]
  wire [2:0] _GEN_2578 = _GEN_325 ? 3'h6 : 3'h7; // @[d_cache.scala 156:47 163:31 166:31]
  wire [40:0] _write_back_addr_T_3 = {_GEN_192,index,3'h0}; // @[Cat.scala 31:58]
  wire  _GEN_2707 = 6'h0 == index ? 1'h0 : dirty_1_0; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2708 = 6'h1 == index ? 1'h0 : dirty_1_1; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2709 = 6'h2 == index ? 1'h0 : dirty_1_2; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2710 = 6'h3 == index ? 1'h0 : dirty_1_3; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2711 = 6'h4 == index ? 1'h0 : dirty_1_4; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2712 = 6'h5 == index ? 1'h0 : dirty_1_5; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2713 = 6'h6 == index ? 1'h0 : dirty_1_6; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2714 = 6'h7 == index ? 1'h0 : dirty_1_7; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2715 = 6'h8 == index ? 1'h0 : dirty_1_8; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2716 = 6'h9 == index ? 1'h0 : dirty_1_9; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2717 = 6'ha == index ? 1'h0 : dirty_1_10; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2718 = 6'hb == index ? 1'h0 : dirty_1_11; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2719 = 6'hc == index ? 1'h0 : dirty_1_12; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2720 = 6'hd == index ? 1'h0 : dirty_1_13; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2721 = 6'he == index ? 1'h0 : dirty_1_14; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2722 = 6'hf == index ? 1'h0 : dirty_1_15; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2723 = 6'h10 == index ? 1'h0 : dirty_1_16; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2724 = 6'h11 == index ? 1'h0 : dirty_1_17; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2725 = 6'h12 == index ? 1'h0 : dirty_1_18; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2726 = 6'h13 == index ? 1'h0 : dirty_1_19; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2727 = 6'h14 == index ? 1'h0 : dirty_1_20; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2728 = 6'h15 == index ? 1'h0 : dirty_1_21; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2729 = 6'h16 == index ? 1'h0 : dirty_1_22; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2730 = 6'h17 == index ? 1'h0 : dirty_1_23; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2731 = 6'h18 == index ? 1'h0 : dirty_1_24; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2732 = 6'h19 == index ? 1'h0 : dirty_1_25; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2733 = 6'h1a == index ? 1'h0 : dirty_1_26; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2734 = 6'h1b == index ? 1'h0 : dirty_1_27; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2735 = 6'h1c == index ? 1'h0 : dirty_1_28; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2736 = 6'h1d == index ? 1'h0 : dirty_1_29; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2737 = 6'h1e == index ? 1'h0 : dirty_1_30; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2738 = 6'h1f == index ? 1'h0 : dirty_1_31; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2739 = 6'h20 == index ? 1'h0 : dirty_1_32; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2740 = 6'h21 == index ? 1'h0 : dirty_1_33; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2741 = 6'h22 == index ? 1'h0 : dirty_1_34; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2742 = 6'h23 == index ? 1'h0 : dirty_1_35; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2743 = 6'h24 == index ? 1'h0 : dirty_1_36; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2744 = 6'h25 == index ? 1'h0 : dirty_1_37; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2745 = 6'h26 == index ? 1'h0 : dirty_1_38; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2746 = 6'h27 == index ? 1'h0 : dirty_1_39; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2747 = 6'h28 == index ? 1'h0 : dirty_1_40; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2748 = 6'h29 == index ? 1'h0 : dirty_1_41; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2749 = 6'h2a == index ? 1'h0 : dirty_1_42; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2750 = 6'h2b == index ? 1'h0 : dirty_1_43; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2751 = 6'h2c == index ? 1'h0 : dirty_1_44; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2752 = 6'h2d == index ? 1'h0 : dirty_1_45; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2753 = 6'h2e == index ? 1'h0 : dirty_1_46; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2754 = 6'h2f == index ? 1'h0 : dirty_1_47; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2755 = 6'h30 == index ? 1'h0 : dirty_1_48; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2756 = 6'h31 == index ? 1'h0 : dirty_1_49; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2757 = 6'h32 == index ? 1'h0 : dirty_1_50; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2758 = 6'h33 == index ? 1'h0 : dirty_1_51; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2759 = 6'h34 == index ? 1'h0 : dirty_1_52; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2760 = 6'h35 == index ? 1'h0 : dirty_1_53; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2761 = 6'h36 == index ? 1'h0 : dirty_1_54; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2762 = 6'h37 == index ? 1'h0 : dirty_1_55; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2763 = 6'h38 == index ? 1'h0 : dirty_1_56; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2764 = 6'h39 == index ? 1'h0 : dirty_1_57; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2765 = 6'h3a == index ? 1'h0 : dirty_1_58; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2766 = 6'h3b == index ? 1'h0 : dirty_1_59; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2767 = 6'h3c == index ? 1'h0 : dirty_1_60; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2768 = 6'h3d == index ? 1'h0 : dirty_1_61; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2769 = 6'h3e == index ? 1'h0 : dirty_1_62; // @[d_cache.scala 178:{40,40} 27:26]
  wire  _GEN_2770 = 6'h3f == index ? 1'h0 : dirty_1_63; // @[d_cache.scala 178:{40,40} 27:26]
  wire [63:0] _GEN_3027 = _GEN_390 ? _GEN_712 : write_back_data; // @[d_cache.scala 173:47 174:41 31:34]
  wire [40:0] _GEN_3028 = _GEN_390 ? _write_back_addr_T_3 : {{9'd0}, write_back_addr}; // @[d_cache.scala 173:47 175:41 32:34]
  wire [63:0] _GEN_3029 = _GEN_390 ? _GEN_1680 : _GEN_1680; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3030 = _GEN_390 ? _GEN_1681 : _GEN_1681; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3031 = _GEN_390 ? _GEN_1682 : _GEN_1682; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3032 = _GEN_390 ? _GEN_1683 : _GEN_1683; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3033 = _GEN_390 ? _GEN_1684 : _GEN_1684; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3034 = _GEN_390 ? _GEN_1685 : _GEN_1685; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3035 = _GEN_390 ? _GEN_1686 : _GEN_1686; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3036 = _GEN_390 ? _GEN_1687 : _GEN_1687; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3037 = _GEN_390 ? _GEN_1688 : _GEN_1688; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3038 = _GEN_390 ? _GEN_1689 : _GEN_1689; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3039 = _GEN_390 ? _GEN_1690 : _GEN_1690; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3040 = _GEN_390 ? _GEN_1691 : _GEN_1691; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3041 = _GEN_390 ? _GEN_1692 : _GEN_1692; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3042 = _GEN_390 ? _GEN_1693 : _GEN_1693; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3043 = _GEN_390 ? _GEN_1694 : _GEN_1694; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3044 = _GEN_390 ? _GEN_1695 : _GEN_1695; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3045 = _GEN_390 ? _GEN_1696 : _GEN_1696; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3046 = _GEN_390 ? _GEN_1697 : _GEN_1697; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3047 = _GEN_390 ? _GEN_1698 : _GEN_1698; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3048 = _GEN_390 ? _GEN_1699 : _GEN_1699; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3049 = _GEN_390 ? _GEN_1700 : _GEN_1700; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3050 = _GEN_390 ? _GEN_1701 : _GEN_1701; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3051 = _GEN_390 ? _GEN_1702 : _GEN_1702; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3052 = _GEN_390 ? _GEN_1703 : _GEN_1703; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3053 = _GEN_390 ? _GEN_1704 : _GEN_1704; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3054 = _GEN_390 ? _GEN_1705 : _GEN_1705; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3055 = _GEN_390 ? _GEN_1706 : _GEN_1706; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3056 = _GEN_390 ? _GEN_1707 : _GEN_1707; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3057 = _GEN_390 ? _GEN_1708 : _GEN_1708; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3058 = _GEN_390 ? _GEN_1709 : _GEN_1709; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3059 = _GEN_390 ? _GEN_1710 : _GEN_1710; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3060 = _GEN_390 ? _GEN_1711 : _GEN_1711; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3061 = _GEN_390 ? _GEN_1712 : _GEN_1712; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3062 = _GEN_390 ? _GEN_1713 : _GEN_1713; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3063 = _GEN_390 ? _GEN_1714 : _GEN_1714; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3064 = _GEN_390 ? _GEN_1715 : _GEN_1715; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3065 = _GEN_390 ? _GEN_1716 : _GEN_1716; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3066 = _GEN_390 ? _GEN_1717 : _GEN_1717; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3067 = _GEN_390 ? _GEN_1718 : _GEN_1718; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3068 = _GEN_390 ? _GEN_1719 : _GEN_1719; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3069 = _GEN_390 ? _GEN_1720 : _GEN_1720; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3070 = _GEN_390 ? _GEN_1721 : _GEN_1721; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3071 = _GEN_390 ? _GEN_1722 : _GEN_1722; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3072 = _GEN_390 ? _GEN_1723 : _GEN_1723; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3073 = _GEN_390 ? _GEN_1724 : _GEN_1724; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3074 = _GEN_390 ? _GEN_1725 : _GEN_1725; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3075 = _GEN_390 ? _GEN_1726 : _GEN_1726; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3076 = _GEN_390 ? _GEN_1727 : _GEN_1727; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3077 = _GEN_390 ? _GEN_1728 : _GEN_1728; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3078 = _GEN_390 ? _GEN_1729 : _GEN_1729; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3079 = _GEN_390 ? _GEN_1730 : _GEN_1730; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3080 = _GEN_390 ? _GEN_1731 : _GEN_1731; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3081 = _GEN_390 ? _GEN_1732 : _GEN_1732; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3082 = _GEN_390 ? _GEN_1733 : _GEN_1733; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3083 = _GEN_390 ? _GEN_1734 : _GEN_1734; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3084 = _GEN_390 ? _GEN_1735 : _GEN_1735; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3085 = _GEN_390 ? _GEN_1736 : _GEN_1736; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3086 = _GEN_390 ? _GEN_1737 : _GEN_1737; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3087 = _GEN_390 ? _GEN_1738 : _GEN_1738; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3088 = _GEN_390 ? _GEN_1739 : _GEN_1739; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3089 = _GEN_390 ? _GEN_1740 : _GEN_1740; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3090 = _GEN_390 ? _GEN_1741 : _GEN_1741; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3091 = _GEN_390 ? _GEN_1742 : _GEN_1742; // @[d_cache.scala 173:47]
  wire [63:0] _GEN_3092 = _GEN_390 ? _GEN_1743 : _GEN_1743; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3093 = _GEN_390 ? _GEN_1744 : _GEN_1744; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3094 = _GEN_390 ? _GEN_1745 : _GEN_1745; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3095 = _GEN_390 ? _GEN_1746 : _GEN_1746; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3096 = _GEN_390 ? _GEN_1747 : _GEN_1747; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3097 = _GEN_390 ? _GEN_1748 : _GEN_1748; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3098 = _GEN_390 ? _GEN_1749 : _GEN_1749; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3099 = _GEN_390 ? _GEN_1750 : _GEN_1750; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3100 = _GEN_390 ? _GEN_1751 : _GEN_1751; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3101 = _GEN_390 ? _GEN_1752 : _GEN_1752; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3102 = _GEN_390 ? _GEN_1753 : _GEN_1753; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3103 = _GEN_390 ? _GEN_1754 : _GEN_1754; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3104 = _GEN_390 ? _GEN_1755 : _GEN_1755; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3105 = _GEN_390 ? _GEN_1756 : _GEN_1756; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3106 = _GEN_390 ? _GEN_1757 : _GEN_1757; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3107 = _GEN_390 ? _GEN_1758 : _GEN_1758; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3108 = _GEN_390 ? _GEN_1759 : _GEN_1759; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3109 = _GEN_390 ? _GEN_1760 : _GEN_1760; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3110 = _GEN_390 ? _GEN_1761 : _GEN_1761; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3111 = _GEN_390 ? _GEN_1762 : _GEN_1762; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3112 = _GEN_390 ? _GEN_1763 : _GEN_1763; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3113 = _GEN_390 ? _GEN_1764 : _GEN_1764; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3114 = _GEN_390 ? _GEN_1765 : _GEN_1765; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3115 = _GEN_390 ? _GEN_1766 : _GEN_1766; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3116 = _GEN_390 ? _GEN_1767 : _GEN_1767; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3117 = _GEN_390 ? _GEN_1768 : _GEN_1768; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3118 = _GEN_390 ? _GEN_1769 : _GEN_1769; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3119 = _GEN_390 ? _GEN_1770 : _GEN_1770; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3120 = _GEN_390 ? _GEN_1771 : _GEN_1771; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3121 = _GEN_390 ? _GEN_1772 : _GEN_1772; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3122 = _GEN_390 ? _GEN_1773 : _GEN_1773; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3123 = _GEN_390 ? _GEN_1774 : _GEN_1774; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3124 = _GEN_390 ? _GEN_1775 : _GEN_1775; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3125 = _GEN_390 ? _GEN_1776 : _GEN_1776; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3126 = _GEN_390 ? _GEN_1777 : _GEN_1777; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3127 = _GEN_390 ? _GEN_1778 : _GEN_1778; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3128 = _GEN_390 ? _GEN_1779 : _GEN_1779; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3129 = _GEN_390 ? _GEN_1780 : _GEN_1780; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3130 = _GEN_390 ? _GEN_1781 : _GEN_1781; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3131 = _GEN_390 ? _GEN_1782 : _GEN_1782; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3132 = _GEN_390 ? _GEN_1783 : _GEN_1783; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3133 = _GEN_390 ? _GEN_1784 : _GEN_1784; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3134 = _GEN_390 ? _GEN_1785 : _GEN_1785; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3135 = _GEN_390 ? _GEN_1786 : _GEN_1786; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3136 = _GEN_390 ? _GEN_1787 : _GEN_1787; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3137 = _GEN_390 ? _GEN_1788 : _GEN_1788; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3138 = _GEN_390 ? _GEN_1789 : _GEN_1789; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3139 = _GEN_390 ? _GEN_1790 : _GEN_1790; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3140 = _GEN_390 ? _GEN_1791 : _GEN_1791; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3141 = _GEN_390 ? _GEN_1792 : _GEN_1792; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3142 = _GEN_390 ? _GEN_1793 : _GEN_1793; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3143 = _GEN_390 ? _GEN_1794 : _GEN_1794; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3144 = _GEN_390 ? _GEN_1795 : _GEN_1795; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3145 = _GEN_390 ? _GEN_1796 : _GEN_1796; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3146 = _GEN_390 ? _GEN_1797 : _GEN_1797; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3147 = _GEN_390 ? _GEN_1798 : _GEN_1798; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3148 = _GEN_390 ? _GEN_1799 : _GEN_1799; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3149 = _GEN_390 ? _GEN_1800 : _GEN_1800; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3150 = _GEN_390 ? _GEN_1801 : _GEN_1801; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3151 = _GEN_390 ? _GEN_1802 : _GEN_1802; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3152 = _GEN_390 ? _GEN_1803 : _GEN_1803; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3153 = _GEN_390 ? _GEN_1804 : _GEN_1804; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3154 = _GEN_390 ? _GEN_1805 : _GEN_1805; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3155 = _GEN_390 ? _GEN_1806 : _GEN_1806; // @[d_cache.scala 173:47]
  wire [31:0] _GEN_3156 = _GEN_390 ? _GEN_1807 : _GEN_1807; // @[d_cache.scala 173:47]
  wire  _GEN_3157 = _GEN_390 ? _GEN_2707 : dirty_1_0; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3158 = _GEN_390 ? _GEN_2708 : dirty_1_1; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3159 = _GEN_390 ? _GEN_2709 : dirty_1_2; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3160 = _GEN_390 ? _GEN_2710 : dirty_1_3; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3161 = _GEN_390 ? _GEN_2711 : dirty_1_4; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3162 = _GEN_390 ? _GEN_2712 : dirty_1_5; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3163 = _GEN_390 ? _GEN_2713 : dirty_1_6; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3164 = _GEN_390 ? _GEN_2714 : dirty_1_7; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3165 = _GEN_390 ? _GEN_2715 : dirty_1_8; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3166 = _GEN_390 ? _GEN_2716 : dirty_1_9; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3167 = _GEN_390 ? _GEN_2717 : dirty_1_10; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3168 = _GEN_390 ? _GEN_2718 : dirty_1_11; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3169 = _GEN_390 ? _GEN_2719 : dirty_1_12; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3170 = _GEN_390 ? _GEN_2720 : dirty_1_13; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3171 = _GEN_390 ? _GEN_2721 : dirty_1_14; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3172 = _GEN_390 ? _GEN_2722 : dirty_1_15; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3173 = _GEN_390 ? _GEN_2723 : dirty_1_16; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3174 = _GEN_390 ? _GEN_2724 : dirty_1_17; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3175 = _GEN_390 ? _GEN_2725 : dirty_1_18; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3176 = _GEN_390 ? _GEN_2726 : dirty_1_19; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3177 = _GEN_390 ? _GEN_2727 : dirty_1_20; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3178 = _GEN_390 ? _GEN_2728 : dirty_1_21; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3179 = _GEN_390 ? _GEN_2729 : dirty_1_22; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3180 = _GEN_390 ? _GEN_2730 : dirty_1_23; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3181 = _GEN_390 ? _GEN_2731 : dirty_1_24; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3182 = _GEN_390 ? _GEN_2732 : dirty_1_25; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3183 = _GEN_390 ? _GEN_2733 : dirty_1_26; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3184 = _GEN_390 ? _GEN_2734 : dirty_1_27; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3185 = _GEN_390 ? _GEN_2735 : dirty_1_28; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3186 = _GEN_390 ? _GEN_2736 : dirty_1_29; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3187 = _GEN_390 ? _GEN_2737 : dirty_1_30; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3188 = _GEN_390 ? _GEN_2738 : dirty_1_31; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3189 = _GEN_390 ? _GEN_2739 : dirty_1_32; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3190 = _GEN_390 ? _GEN_2740 : dirty_1_33; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3191 = _GEN_390 ? _GEN_2741 : dirty_1_34; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3192 = _GEN_390 ? _GEN_2742 : dirty_1_35; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3193 = _GEN_390 ? _GEN_2743 : dirty_1_36; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3194 = _GEN_390 ? _GEN_2744 : dirty_1_37; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3195 = _GEN_390 ? _GEN_2745 : dirty_1_38; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3196 = _GEN_390 ? _GEN_2746 : dirty_1_39; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3197 = _GEN_390 ? _GEN_2747 : dirty_1_40; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3198 = _GEN_390 ? _GEN_2748 : dirty_1_41; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3199 = _GEN_390 ? _GEN_2749 : dirty_1_42; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3200 = _GEN_390 ? _GEN_2750 : dirty_1_43; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3201 = _GEN_390 ? _GEN_2751 : dirty_1_44; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3202 = _GEN_390 ? _GEN_2752 : dirty_1_45; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3203 = _GEN_390 ? _GEN_2753 : dirty_1_46; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3204 = _GEN_390 ? _GEN_2754 : dirty_1_47; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3205 = _GEN_390 ? _GEN_2755 : dirty_1_48; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3206 = _GEN_390 ? _GEN_2756 : dirty_1_49; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3207 = _GEN_390 ? _GEN_2757 : dirty_1_50; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3208 = _GEN_390 ? _GEN_2758 : dirty_1_51; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3209 = _GEN_390 ? _GEN_2759 : dirty_1_52; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3210 = _GEN_390 ? _GEN_2760 : dirty_1_53; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3211 = _GEN_390 ? _GEN_2761 : dirty_1_54; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3212 = _GEN_390 ? _GEN_2762 : dirty_1_55; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3213 = _GEN_390 ? _GEN_2763 : dirty_1_56; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3214 = _GEN_390 ? _GEN_2764 : dirty_1_57; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3215 = _GEN_390 ? _GEN_2765 : dirty_1_58; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3216 = _GEN_390 ? _GEN_2766 : dirty_1_59; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3217 = _GEN_390 ? _GEN_2767 : dirty_1_60; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3218 = _GEN_390 ? _GEN_2768 : dirty_1_61; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3219 = _GEN_390 ? _GEN_2769 : dirty_1_62; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3220 = _GEN_390 ? _GEN_2770 : dirty_1_63; // @[d_cache.scala 173:47 27:26]
  wire  _GEN_3221 = _GEN_390 ? _GEN_777 : _GEN_777; // @[d_cache.scala 173:47]
  wire  _GEN_3222 = _GEN_390 ? _GEN_778 : _GEN_778; // @[d_cache.scala 173:47]
  wire  _GEN_3223 = _GEN_390 ? _GEN_779 : _GEN_779; // @[d_cache.scala 173:47]
  wire  _GEN_3224 = _GEN_390 ? _GEN_780 : _GEN_780; // @[d_cache.scala 173:47]
  wire  _GEN_3225 = _GEN_390 ? _GEN_781 : _GEN_781; // @[d_cache.scala 173:47]
  wire  _GEN_3226 = _GEN_390 ? _GEN_782 : _GEN_782; // @[d_cache.scala 173:47]
  wire  _GEN_3227 = _GEN_390 ? _GEN_783 : _GEN_783; // @[d_cache.scala 173:47]
  wire  _GEN_3228 = _GEN_390 ? _GEN_784 : _GEN_784; // @[d_cache.scala 173:47]
  wire  _GEN_3229 = _GEN_390 ? _GEN_785 : _GEN_785; // @[d_cache.scala 173:47]
  wire  _GEN_3230 = _GEN_390 ? _GEN_786 : _GEN_786; // @[d_cache.scala 173:47]
  wire  _GEN_3231 = _GEN_390 ? _GEN_787 : _GEN_787; // @[d_cache.scala 173:47]
  wire  _GEN_3232 = _GEN_390 ? _GEN_788 : _GEN_788; // @[d_cache.scala 173:47]
  wire  _GEN_3233 = _GEN_390 ? _GEN_789 : _GEN_789; // @[d_cache.scala 173:47]
  wire  _GEN_3234 = _GEN_390 ? _GEN_790 : _GEN_790; // @[d_cache.scala 173:47]
  wire  _GEN_3235 = _GEN_390 ? _GEN_791 : _GEN_791; // @[d_cache.scala 173:47]
  wire  _GEN_3236 = _GEN_390 ? _GEN_792 : _GEN_792; // @[d_cache.scala 173:47]
  wire  _GEN_3237 = _GEN_390 ? _GEN_793 : _GEN_793; // @[d_cache.scala 173:47]
  wire  _GEN_3238 = _GEN_390 ? _GEN_794 : _GEN_794; // @[d_cache.scala 173:47]
  wire  _GEN_3239 = _GEN_390 ? _GEN_795 : _GEN_795; // @[d_cache.scala 173:47]
  wire  _GEN_3240 = _GEN_390 ? _GEN_796 : _GEN_796; // @[d_cache.scala 173:47]
  wire  _GEN_3241 = _GEN_390 ? _GEN_797 : _GEN_797; // @[d_cache.scala 173:47]
  wire  _GEN_3242 = _GEN_390 ? _GEN_798 : _GEN_798; // @[d_cache.scala 173:47]
  wire  _GEN_3243 = _GEN_390 ? _GEN_799 : _GEN_799; // @[d_cache.scala 173:47]
  wire  _GEN_3244 = _GEN_390 ? _GEN_800 : _GEN_800; // @[d_cache.scala 173:47]
  wire  _GEN_3245 = _GEN_390 ? _GEN_801 : _GEN_801; // @[d_cache.scala 173:47]
  wire  _GEN_3246 = _GEN_390 ? _GEN_802 : _GEN_802; // @[d_cache.scala 173:47]
  wire  _GEN_3247 = _GEN_390 ? _GEN_803 : _GEN_803; // @[d_cache.scala 173:47]
  wire  _GEN_3248 = _GEN_390 ? _GEN_804 : _GEN_804; // @[d_cache.scala 173:47]
  wire  _GEN_3249 = _GEN_390 ? _GEN_805 : _GEN_805; // @[d_cache.scala 173:47]
  wire  _GEN_3250 = _GEN_390 ? _GEN_806 : _GEN_806; // @[d_cache.scala 173:47]
  wire  _GEN_3251 = _GEN_390 ? _GEN_807 : _GEN_807; // @[d_cache.scala 173:47]
  wire  _GEN_3252 = _GEN_390 ? _GEN_808 : _GEN_808; // @[d_cache.scala 173:47]
  wire  _GEN_3253 = _GEN_390 ? _GEN_809 : _GEN_809; // @[d_cache.scala 173:47]
  wire  _GEN_3254 = _GEN_390 ? _GEN_810 : _GEN_810; // @[d_cache.scala 173:47]
  wire  _GEN_3255 = _GEN_390 ? _GEN_811 : _GEN_811; // @[d_cache.scala 173:47]
  wire  _GEN_3256 = _GEN_390 ? _GEN_812 : _GEN_812; // @[d_cache.scala 173:47]
  wire  _GEN_3257 = _GEN_390 ? _GEN_813 : _GEN_813; // @[d_cache.scala 173:47]
  wire  _GEN_3258 = _GEN_390 ? _GEN_814 : _GEN_814; // @[d_cache.scala 173:47]
  wire  _GEN_3259 = _GEN_390 ? _GEN_815 : _GEN_815; // @[d_cache.scala 173:47]
  wire  _GEN_3260 = _GEN_390 ? _GEN_816 : _GEN_816; // @[d_cache.scala 173:47]
  wire  _GEN_3261 = _GEN_390 ? _GEN_817 : _GEN_817; // @[d_cache.scala 173:47]
  wire  _GEN_3262 = _GEN_390 ? _GEN_818 : _GEN_818; // @[d_cache.scala 173:47]
  wire  _GEN_3263 = _GEN_390 ? _GEN_819 : _GEN_819; // @[d_cache.scala 173:47]
  wire  _GEN_3264 = _GEN_390 ? _GEN_820 : _GEN_820; // @[d_cache.scala 173:47]
  wire  _GEN_3265 = _GEN_390 ? _GEN_821 : _GEN_821; // @[d_cache.scala 173:47]
  wire  _GEN_3266 = _GEN_390 ? _GEN_822 : _GEN_822; // @[d_cache.scala 173:47]
  wire  _GEN_3267 = _GEN_390 ? _GEN_823 : _GEN_823; // @[d_cache.scala 173:47]
  wire  _GEN_3268 = _GEN_390 ? _GEN_824 : _GEN_824; // @[d_cache.scala 173:47]
  wire  _GEN_3269 = _GEN_390 ? _GEN_825 : _GEN_825; // @[d_cache.scala 173:47]
  wire  _GEN_3270 = _GEN_390 ? _GEN_826 : _GEN_826; // @[d_cache.scala 173:47]
  wire  _GEN_3271 = _GEN_390 ? _GEN_827 : _GEN_827; // @[d_cache.scala 173:47]
  wire  _GEN_3272 = _GEN_390 ? _GEN_828 : _GEN_828; // @[d_cache.scala 173:47]
  wire  _GEN_3273 = _GEN_390 ? _GEN_829 : _GEN_829; // @[d_cache.scala 173:47]
  wire  _GEN_3274 = _GEN_390 ? _GEN_830 : _GEN_830; // @[d_cache.scala 173:47]
  wire  _GEN_3275 = _GEN_390 ? _GEN_831 : _GEN_831; // @[d_cache.scala 173:47]
  wire  _GEN_3276 = _GEN_390 ? _GEN_832 : _GEN_832; // @[d_cache.scala 173:47]
  wire  _GEN_3277 = _GEN_390 ? _GEN_833 : _GEN_833; // @[d_cache.scala 173:47]
  wire  _GEN_3278 = _GEN_390 ? _GEN_834 : _GEN_834; // @[d_cache.scala 173:47]
  wire  _GEN_3279 = _GEN_390 ? _GEN_835 : _GEN_835; // @[d_cache.scala 173:47]
  wire  _GEN_3280 = _GEN_390 ? _GEN_836 : _GEN_836; // @[d_cache.scala 173:47]
  wire  _GEN_3281 = _GEN_390 ? _GEN_837 : _GEN_837; // @[d_cache.scala 173:47]
  wire  _GEN_3282 = _GEN_390 ? _GEN_838 : _GEN_838; // @[d_cache.scala 173:47]
  wire  _GEN_3283 = _GEN_390 ? _GEN_839 : _GEN_839; // @[d_cache.scala 173:47]
  wire  _GEN_3284 = _GEN_390 ? _GEN_840 : _GEN_840; // @[d_cache.scala 173:47]
  wire [2:0] _GEN_3285 = _GEN_390 ? 3'h6 : 3'h7; // @[d_cache.scala 173:47 180:31 183:31]
  wire [63:0] _GEN_3286 = ~quene ? _GEN_2320 : _GEN_3027; // @[d_cache.scala 154:34]
  wire [40:0] _GEN_3287 = ~quene ? _GEN_2321 : _GEN_3028; // @[d_cache.scala 154:34]
  wire [63:0] _GEN_3288 = ~quene ? _GEN_2322 : ram_0_0; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3289 = ~quene ? _GEN_2323 : ram_0_1; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3290 = ~quene ? _GEN_2324 : ram_0_2; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3291 = ~quene ? _GEN_2325 : ram_0_3; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3292 = ~quene ? _GEN_2326 : ram_0_4; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3293 = ~quene ? _GEN_2327 : ram_0_5; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3294 = ~quene ? _GEN_2328 : ram_0_6; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3295 = ~quene ? _GEN_2329 : ram_0_7; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3296 = ~quene ? _GEN_2330 : ram_0_8; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3297 = ~quene ? _GEN_2331 : ram_0_9; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3298 = ~quene ? _GEN_2332 : ram_0_10; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3299 = ~quene ? _GEN_2333 : ram_0_11; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3300 = ~quene ? _GEN_2334 : ram_0_12; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3301 = ~quene ? _GEN_2335 : ram_0_13; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3302 = ~quene ? _GEN_2336 : ram_0_14; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3303 = ~quene ? _GEN_2337 : ram_0_15; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3304 = ~quene ? _GEN_2338 : ram_0_16; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3305 = ~quene ? _GEN_2339 : ram_0_17; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3306 = ~quene ? _GEN_2340 : ram_0_18; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3307 = ~quene ? _GEN_2341 : ram_0_19; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3308 = ~quene ? _GEN_2342 : ram_0_20; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3309 = ~quene ? _GEN_2343 : ram_0_21; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3310 = ~quene ? _GEN_2344 : ram_0_22; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3311 = ~quene ? _GEN_2345 : ram_0_23; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3312 = ~quene ? _GEN_2346 : ram_0_24; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3313 = ~quene ? _GEN_2347 : ram_0_25; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3314 = ~quene ? _GEN_2348 : ram_0_26; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3315 = ~quene ? _GEN_2349 : ram_0_27; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3316 = ~quene ? _GEN_2350 : ram_0_28; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3317 = ~quene ? _GEN_2351 : ram_0_29; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3318 = ~quene ? _GEN_2352 : ram_0_30; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3319 = ~quene ? _GEN_2353 : ram_0_31; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3320 = ~quene ? _GEN_2354 : ram_0_32; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3321 = ~quene ? _GEN_2355 : ram_0_33; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3322 = ~quene ? _GEN_2356 : ram_0_34; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3323 = ~quene ? _GEN_2357 : ram_0_35; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3324 = ~quene ? _GEN_2358 : ram_0_36; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3325 = ~quene ? _GEN_2359 : ram_0_37; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3326 = ~quene ? _GEN_2360 : ram_0_38; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3327 = ~quene ? _GEN_2361 : ram_0_39; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3328 = ~quene ? _GEN_2362 : ram_0_40; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3329 = ~quene ? _GEN_2363 : ram_0_41; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3330 = ~quene ? _GEN_2364 : ram_0_42; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3331 = ~quene ? _GEN_2365 : ram_0_43; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3332 = ~quene ? _GEN_2366 : ram_0_44; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3333 = ~quene ? _GEN_2367 : ram_0_45; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3334 = ~quene ? _GEN_2368 : ram_0_46; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3335 = ~quene ? _GEN_2369 : ram_0_47; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3336 = ~quene ? _GEN_2370 : ram_0_48; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3337 = ~quene ? _GEN_2371 : ram_0_49; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3338 = ~quene ? _GEN_2372 : ram_0_50; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3339 = ~quene ? _GEN_2373 : ram_0_51; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3340 = ~quene ? _GEN_2374 : ram_0_52; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3341 = ~quene ? _GEN_2375 : ram_0_53; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3342 = ~quene ? _GEN_2376 : ram_0_54; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3343 = ~quene ? _GEN_2377 : ram_0_55; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3344 = ~quene ? _GEN_2378 : ram_0_56; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3345 = ~quene ? _GEN_2379 : ram_0_57; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3346 = ~quene ? _GEN_2380 : ram_0_58; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3347 = ~quene ? _GEN_2381 : ram_0_59; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3348 = ~quene ? _GEN_2382 : ram_0_60; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3349 = ~quene ? _GEN_2383 : ram_0_61; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3350 = ~quene ? _GEN_2384 : ram_0_62; // @[d_cache.scala 154:34 18:24]
  wire [63:0] _GEN_3351 = ~quene ? _GEN_2385 : ram_0_63; // @[d_cache.scala 154:34 18:24]
  wire [31:0] _GEN_3352 = ~quene ? _GEN_2386 : tag_0_0; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3353 = ~quene ? _GEN_2387 : tag_0_1; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3354 = ~quene ? _GEN_2388 : tag_0_2; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3355 = ~quene ? _GEN_2389 : tag_0_3; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3356 = ~quene ? _GEN_2390 : tag_0_4; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3357 = ~quene ? _GEN_2391 : tag_0_5; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3358 = ~quene ? _GEN_2392 : tag_0_6; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3359 = ~quene ? _GEN_2393 : tag_0_7; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3360 = ~quene ? _GEN_2394 : tag_0_8; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3361 = ~quene ? _GEN_2395 : tag_0_9; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3362 = ~quene ? _GEN_2396 : tag_0_10; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3363 = ~quene ? _GEN_2397 : tag_0_11; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3364 = ~quene ? _GEN_2398 : tag_0_12; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3365 = ~quene ? _GEN_2399 : tag_0_13; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3366 = ~quene ? _GEN_2400 : tag_0_14; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3367 = ~quene ? _GEN_2401 : tag_0_15; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3368 = ~quene ? _GEN_2402 : tag_0_16; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3369 = ~quene ? _GEN_2403 : tag_0_17; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3370 = ~quene ? _GEN_2404 : tag_0_18; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3371 = ~quene ? _GEN_2405 : tag_0_19; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3372 = ~quene ? _GEN_2406 : tag_0_20; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3373 = ~quene ? _GEN_2407 : tag_0_21; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3374 = ~quene ? _GEN_2408 : tag_0_22; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3375 = ~quene ? _GEN_2409 : tag_0_23; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3376 = ~quene ? _GEN_2410 : tag_0_24; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3377 = ~quene ? _GEN_2411 : tag_0_25; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3378 = ~quene ? _GEN_2412 : tag_0_26; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3379 = ~quene ? _GEN_2413 : tag_0_27; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3380 = ~quene ? _GEN_2414 : tag_0_28; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3381 = ~quene ? _GEN_2415 : tag_0_29; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3382 = ~quene ? _GEN_2416 : tag_0_30; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3383 = ~quene ? _GEN_2417 : tag_0_31; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3384 = ~quene ? _GEN_2418 : tag_0_32; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3385 = ~quene ? _GEN_2419 : tag_0_33; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3386 = ~quene ? _GEN_2420 : tag_0_34; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3387 = ~quene ? _GEN_2421 : tag_0_35; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3388 = ~quene ? _GEN_2422 : tag_0_36; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3389 = ~quene ? _GEN_2423 : tag_0_37; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3390 = ~quene ? _GEN_2424 : tag_0_38; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3391 = ~quene ? _GEN_2425 : tag_0_39; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3392 = ~quene ? _GEN_2426 : tag_0_40; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3393 = ~quene ? _GEN_2427 : tag_0_41; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3394 = ~quene ? _GEN_2428 : tag_0_42; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3395 = ~quene ? _GEN_2429 : tag_0_43; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3396 = ~quene ? _GEN_2430 : tag_0_44; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3397 = ~quene ? _GEN_2431 : tag_0_45; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3398 = ~quene ? _GEN_2432 : tag_0_46; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3399 = ~quene ? _GEN_2433 : tag_0_47; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3400 = ~quene ? _GEN_2434 : tag_0_48; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3401 = ~quene ? _GEN_2435 : tag_0_49; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3402 = ~quene ? _GEN_2436 : tag_0_50; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3403 = ~quene ? _GEN_2437 : tag_0_51; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3404 = ~quene ? _GEN_2438 : tag_0_52; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3405 = ~quene ? _GEN_2439 : tag_0_53; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3406 = ~quene ? _GEN_2440 : tag_0_54; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3407 = ~quene ? _GEN_2441 : tag_0_55; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3408 = ~quene ? _GEN_2442 : tag_0_56; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3409 = ~quene ? _GEN_2443 : tag_0_57; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3410 = ~quene ? _GEN_2444 : tag_0_58; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3411 = ~quene ? _GEN_2445 : tag_0_59; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3412 = ~quene ? _GEN_2446 : tag_0_60; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3413 = ~quene ? _GEN_2447 : tag_0_61; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3414 = ~quene ? _GEN_2448 : tag_0_62; // @[d_cache.scala 154:34 22:24]
  wire [31:0] _GEN_3415 = ~quene ? _GEN_2449 : tag_0_63; // @[d_cache.scala 154:34 22:24]
  wire  _GEN_3416 = ~quene ? _GEN_2450 : dirty_0_0; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3417 = ~quene ? _GEN_2451 : dirty_0_1; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3418 = ~quene ? _GEN_2452 : dirty_0_2; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3419 = ~quene ? _GEN_2453 : dirty_0_3; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3420 = ~quene ? _GEN_2454 : dirty_0_4; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3421 = ~quene ? _GEN_2455 : dirty_0_5; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3422 = ~quene ? _GEN_2456 : dirty_0_6; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3423 = ~quene ? _GEN_2457 : dirty_0_7; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3424 = ~quene ? _GEN_2458 : dirty_0_8; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3425 = ~quene ? _GEN_2459 : dirty_0_9; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3426 = ~quene ? _GEN_2460 : dirty_0_10; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3427 = ~quene ? _GEN_2461 : dirty_0_11; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3428 = ~quene ? _GEN_2462 : dirty_0_12; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3429 = ~quene ? _GEN_2463 : dirty_0_13; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3430 = ~quene ? _GEN_2464 : dirty_0_14; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3431 = ~quene ? _GEN_2465 : dirty_0_15; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3432 = ~quene ? _GEN_2466 : dirty_0_16; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3433 = ~quene ? _GEN_2467 : dirty_0_17; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3434 = ~quene ? _GEN_2468 : dirty_0_18; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3435 = ~quene ? _GEN_2469 : dirty_0_19; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3436 = ~quene ? _GEN_2470 : dirty_0_20; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3437 = ~quene ? _GEN_2471 : dirty_0_21; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3438 = ~quene ? _GEN_2472 : dirty_0_22; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3439 = ~quene ? _GEN_2473 : dirty_0_23; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3440 = ~quene ? _GEN_2474 : dirty_0_24; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3441 = ~quene ? _GEN_2475 : dirty_0_25; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3442 = ~quene ? _GEN_2476 : dirty_0_26; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3443 = ~quene ? _GEN_2477 : dirty_0_27; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3444 = ~quene ? _GEN_2478 : dirty_0_28; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3445 = ~quene ? _GEN_2479 : dirty_0_29; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3446 = ~quene ? _GEN_2480 : dirty_0_30; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3447 = ~quene ? _GEN_2481 : dirty_0_31; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3448 = ~quene ? _GEN_2482 : dirty_0_32; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3449 = ~quene ? _GEN_2483 : dirty_0_33; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3450 = ~quene ? _GEN_2484 : dirty_0_34; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3451 = ~quene ? _GEN_2485 : dirty_0_35; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3452 = ~quene ? _GEN_2486 : dirty_0_36; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3453 = ~quene ? _GEN_2487 : dirty_0_37; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3454 = ~quene ? _GEN_2488 : dirty_0_38; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3455 = ~quene ? _GEN_2489 : dirty_0_39; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3456 = ~quene ? _GEN_2490 : dirty_0_40; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3457 = ~quene ? _GEN_2491 : dirty_0_41; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3458 = ~quene ? _GEN_2492 : dirty_0_42; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3459 = ~quene ? _GEN_2493 : dirty_0_43; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3460 = ~quene ? _GEN_2494 : dirty_0_44; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3461 = ~quene ? _GEN_2495 : dirty_0_45; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3462 = ~quene ? _GEN_2496 : dirty_0_46; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3463 = ~quene ? _GEN_2497 : dirty_0_47; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3464 = ~quene ? _GEN_2498 : dirty_0_48; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3465 = ~quene ? _GEN_2499 : dirty_0_49; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3466 = ~quene ? _GEN_2500 : dirty_0_50; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3467 = ~quene ? _GEN_2501 : dirty_0_51; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3468 = ~quene ? _GEN_2502 : dirty_0_52; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3469 = ~quene ? _GEN_2503 : dirty_0_53; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3470 = ~quene ? _GEN_2504 : dirty_0_54; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3471 = ~quene ? _GEN_2505 : dirty_0_55; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3472 = ~quene ? _GEN_2506 : dirty_0_56; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3473 = ~quene ? _GEN_2507 : dirty_0_57; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3474 = ~quene ? _GEN_2508 : dirty_0_58; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3475 = ~quene ? _GEN_2509 : dirty_0_59; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3476 = ~quene ? _GEN_2510 : dirty_0_60; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3477 = ~quene ? _GEN_2511 : dirty_0_61; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3478 = ~quene ? _GEN_2512 : dirty_0_62; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3479 = ~quene ? _GEN_2513 : dirty_0_63; // @[d_cache.scala 154:34 26:26]
  wire  _GEN_3480 = ~quene ? _GEN_2514 : valid_0_0; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3481 = ~quene ? _GEN_2515 : valid_0_1; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3482 = ~quene ? _GEN_2516 : valid_0_2; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3483 = ~quene ? _GEN_2517 : valid_0_3; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3484 = ~quene ? _GEN_2518 : valid_0_4; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3485 = ~quene ? _GEN_2519 : valid_0_5; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3486 = ~quene ? _GEN_2520 : valid_0_6; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3487 = ~quene ? _GEN_2521 : valid_0_7; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3488 = ~quene ? _GEN_2522 : valid_0_8; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3489 = ~quene ? _GEN_2523 : valid_0_9; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3490 = ~quene ? _GEN_2524 : valid_0_10; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3491 = ~quene ? _GEN_2525 : valid_0_11; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3492 = ~quene ? _GEN_2526 : valid_0_12; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3493 = ~quene ? _GEN_2527 : valid_0_13; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3494 = ~quene ? _GEN_2528 : valid_0_14; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3495 = ~quene ? _GEN_2529 : valid_0_15; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3496 = ~quene ? _GEN_2530 : valid_0_16; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3497 = ~quene ? _GEN_2531 : valid_0_17; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3498 = ~quene ? _GEN_2532 : valid_0_18; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3499 = ~quene ? _GEN_2533 : valid_0_19; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3500 = ~quene ? _GEN_2534 : valid_0_20; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3501 = ~quene ? _GEN_2535 : valid_0_21; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3502 = ~quene ? _GEN_2536 : valid_0_22; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3503 = ~quene ? _GEN_2537 : valid_0_23; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3504 = ~quene ? _GEN_2538 : valid_0_24; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3505 = ~quene ? _GEN_2539 : valid_0_25; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3506 = ~quene ? _GEN_2540 : valid_0_26; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3507 = ~quene ? _GEN_2541 : valid_0_27; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3508 = ~quene ? _GEN_2542 : valid_0_28; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3509 = ~quene ? _GEN_2543 : valid_0_29; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3510 = ~quene ? _GEN_2544 : valid_0_30; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3511 = ~quene ? _GEN_2545 : valid_0_31; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3512 = ~quene ? _GEN_2546 : valid_0_32; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3513 = ~quene ? _GEN_2547 : valid_0_33; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3514 = ~quene ? _GEN_2548 : valid_0_34; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3515 = ~quene ? _GEN_2549 : valid_0_35; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3516 = ~quene ? _GEN_2550 : valid_0_36; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3517 = ~quene ? _GEN_2551 : valid_0_37; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3518 = ~quene ? _GEN_2552 : valid_0_38; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3519 = ~quene ? _GEN_2553 : valid_0_39; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3520 = ~quene ? _GEN_2554 : valid_0_40; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3521 = ~quene ? _GEN_2555 : valid_0_41; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3522 = ~quene ? _GEN_2556 : valid_0_42; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3523 = ~quene ? _GEN_2557 : valid_0_43; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3524 = ~quene ? _GEN_2558 : valid_0_44; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3525 = ~quene ? _GEN_2559 : valid_0_45; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3526 = ~quene ? _GEN_2560 : valid_0_46; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3527 = ~quene ? _GEN_2561 : valid_0_47; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3528 = ~quene ? _GEN_2562 : valid_0_48; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3529 = ~quene ? _GEN_2563 : valid_0_49; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3530 = ~quene ? _GEN_2564 : valid_0_50; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3531 = ~quene ? _GEN_2565 : valid_0_51; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3532 = ~quene ? _GEN_2566 : valid_0_52; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3533 = ~quene ? _GEN_2567 : valid_0_53; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3534 = ~quene ? _GEN_2568 : valid_0_54; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3535 = ~quene ? _GEN_2569 : valid_0_55; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3536 = ~quene ? _GEN_2570 : valid_0_56; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3537 = ~quene ? _GEN_2571 : valid_0_57; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3538 = ~quene ? _GEN_2572 : valid_0_58; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3539 = ~quene ? _GEN_2573 : valid_0_59; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3540 = ~quene ? _GEN_2574 : valid_0_60; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3541 = ~quene ? _GEN_2575 : valid_0_61; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3542 = ~quene ? _GEN_2576 : valid_0_62; // @[d_cache.scala 154:34 24:26]
  wire  _GEN_3543 = ~quene ? _GEN_2577 : valid_0_63; // @[d_cache.scala 154:34 24:26]
  wire [2:0] _GEN_3544 = ~quene ? _GEN_2578 : _GEN_3285; // @[d_cache.scala 154:34]
  wire [63:0] _GEN_3545 = ~quene ? ram_1_0 : _GEN_3029; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3546 = ~quene ? ram_1_1 : _GEN_3030; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3547 = ~quene ? ram_1_2 : _GEN_3031; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3548 = ~quene ? ram_1_3 : _GEN_3032; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3549 = ~quene ? ram_1_4 : _GEN_3033; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3550 = ~quene ? ram_1_5 : _GEN_3034; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3551 = ~quene ? ram_1_6 : _GEN_3035; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3552 = ~quene ? ram_1_7 : _GEN_3036; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3553 = ~quene ? ram_1_8 : _GEN_3037; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3554 = ~quene ? ram_1_9 : _GEN_3038; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3555 = ~quene ? ram_1_10 : _GEN_3039; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3556 = ~quene ? ram_1_11 : _GEN_3040; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3557 = ~quene ? ram_1_12 : _GEN_3041; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3558 = ~quene ? ram_1_13 : _GEN_3042; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3559 = ~quene ? ram_1_14 : _GEN_3043; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3560 = ~quene ? ram_1_15 : _GEN_3044; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3561 = ~quene ? ram_1_16 : _GEN_3045; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3562 = ~quene ? ram_1_17 : _GEN_3046; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3563 = ~quene ? ram_1_18 : _GEN_3047; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3564 = ~quene ? ram_1_19 : _GEN_3048; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3565 = ~quene ? ram_1_20 : _GEN_3049; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3566 = ~quene ? ram_1_21 : _GEN_3050; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3567 = ~quene ? ram_1_22 : _GEN_3051; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3568 = ~quene ? ram_1_23 : _GEN_3052; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3569 = ~quene ? ram_1_24 : _GEN_3053; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3570 = ~quene ? ram_1_25 : _GEN_3054; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3571 = ~quene ? ram_1_26 : _GEN_3055; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3572 = ~quene ? ram_1_27 : _GEN_3056; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3573 = ~quene ? ram_1_28 : _GEN_3057; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3574 = ~quene ? ram_1_29 : _GEN_3058; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3575 = ~quene ? ram_1_30 : _GEN_3059; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3576 = ~quene ? ram_1_31 : _GEN_3060; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3577 = ~quene ? ram_1_32 : _GEN_3061; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3578 = ~quene ? ram_1_33 : _GEN_3062; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3579 = ~quene ? ram_1_34 : _GEN_3063; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3580 = ~quene ? ram_1_35 : _GEN_3064; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3581 = ~quene ? ram_1_36 : _GEN_3065; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3582 = ~quene ? ram_1_37 : _GEN_3066; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3583 = ~quene ? ram_1_38 : _GEN_3067; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3584 = ~quene ? ram_1_39 : _GEN_3068; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3585 = ~quene ? ram_1_40 : _GEN_3069; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3586 = ~quene ? ram_1_41 : _GEN_3070; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3587 = ~quene ? ram_1_42 : _GEN_3071; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3588 = ~quene ? ram_1_43 : _GEN_3072; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3589 = ~quene ? ram_1_44 : _GEN_3073; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3590 = ~quene ? ram_1_45 : _GEN_3074; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3591 = ~quene ? ram_1_46 : _GEN_3075; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3592 = ~quene ? ram_1_47 : _GEN_3076; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3593 = ~quene ? ram_1_48 : _GEN_3077; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3594 = ~quene ? ram_1_49 : _GEN_3078; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3595 = ~quene ? ram_1_50 : _GEN_3079; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3596 = ~quene ? ram_1_51 : _GEN_3080; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3597 = ~quene ? ram_1_52 : _GEN_3081; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3598 = ~quene ? ram_1_53 : _GEN_3082; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3599 = ~quene ? ram_1_54 : _GEN_3083; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3600 = ~quene ? ram_1_55 : _GEN_3084; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3601 = ~quene ? ram_1_56 : _GEN_3085; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3602 = ~quene ? ram_1_57 : _GEN_3086; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3603 = ~quene ? ram_1_58 : _GEN_3087; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3604 = ~quene ? ram_1_59 : _GEN_3088; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3605 = ~quene ? ram_1_60 : _GEN_3089; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3606 = ~quene ? ram_1_61 : _GEN_3090; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3607 = ~quene ? ram_1_62 : _GEN_3091; // @[d_cache.scala 154:34 19:24]
  wire [63:0] _GEN_3608 = ~quene ? ram_1_63 : _GEN_3092; // @[d_cache.scala 154:34 19:24]
  wire [31:0] _GEN_3609 = ~quene ? tag_1_0 : _GEN_3093; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3610 = ~quene ? tag_1_1 : _GEN_3094; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3611 = ~quene ? tag_1_2 : _GEN_3095; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3612 = ~quene ? tag_1_3 : _GEN_3096; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3613 = ~quene ? tag_1_4 : _GEN_3097; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3614 = ~quene ? tag_1_5 : _GEN_3098; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3615 = ~quene ? tag_1_6 : _GEN_3099; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3616 = ~quene ? tag_1_7 : _GEN_3100; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3617 = ~quene ? tag_1_8 : _GEN_3101; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3618 = ~quene ? tag_1_9 : _GEN_3102; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3619 = ~quene ? tag_1_10 : _GEN_3103; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3620 = ~quene ? tag_1_11 : _GEN_3104; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3621 = ~quene ? tag_1_12 : _GEN_3105; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3622 = ~quene ? tag_1_13 : _GEN_3106; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3623 = ~quene ? tag_1_14 : _GEN_3107; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3624 = ~quene ? tag_1_15 : _GEN_3108; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3625 = ~quene ? tag_1_16 : _GEN_3109; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3626 = ~quene ? tag_1_17 : _GEN_3110; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3627 = ~quene ? tag_1_18 : _GEN_3111; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3628 = ~quene ? tag_1_19 : _GEN_3112; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3629 = ~quene ? tag_1_20 : _GEN_3113; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3630 = ~quene ? tag_1_21 : _GEN_3114; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3631 = ~quene ? tag_1_22 : _GEN_3115; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3632 = ~quene ? tag_1_23 : _GEN_3116; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3633 = ~quene ? tag_1_24 : _GEN_3117; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3634 = ~quene ? tag_1_25 : _GEN_3118; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3635 = ~quene ? tag_1_26 : _GEN_3119; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3636 = ~quene ? tag_1_27 : _GEN_3120; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3637 = ~quene ? tag_1_28 : _GEN_3121; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3638 = ~quene ? tag_1_29 : _GEN_3122; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3639 = ~quene ? tag_1_30 : _GEN_3123; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3640 = ~quene ? tag_1_31 : _GEN_3124; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3641 = ~quene ? tag_1_32 : _GEN_3125; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3642 = ~quene ? tag_1_33 : _GEN_3126; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3643 = ~quene ? tag_1_34 : _GEN_3127; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3644 = ~quene ? tag_1_35 : _GEN_3128; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3645 = ~quene ? tag_1_36 : _GEN_3129; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3646 = ~quene ? tag_1_37 : _GEN_3130; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3647 = ~quene ? tag_1_38 : _GEN_3131; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3648 = ~quene ? tag_1_39 : _GEN_3132; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3649 = ~quene ? tag_1_40 : _GEN_3133; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3650 = ~quene ? tag_1_41 : _GEN_3134; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3651 = ~quene ? tag_1_42 : _GEN_3135; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3652 = ~quene ? tag_1_43 : _GEN_3136; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3653 = ~quene ? tag_1_44 : _GEN_3137; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3654 = ~quene ? tag_1_45 : _GEN_3138; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3655 = ~quene ? tag_1_46 : _GEN_3139; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3656 = ~quene ? tag_1_47 : _GEN_3140; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3657 = ~quene ? tag_1_48 : _GEN_3141; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3658 = ~quene ? tag_1_49 : _GEN_3142; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3659 = ~quene ? tag_1_50 : _GEN_3143; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3660 = ~quene ? tag_1_51 : _GEN_3144; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3661 = ~quene ? tag_1_52 : _GEN_3145; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3662 = ~quene ? tag_1_53 : _GEN_3146; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3663 = ~quene ? tag_1_54 : _GEN_3147; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3664 = ~quene ? tag_1_55 : _GEN_3148; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3665 = ~quene ? tag_1_56 : _GEN_3149; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3666 = ~quene ? tag_1_57 : _GEN_3150; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3667 = ~quene ? tag_1_58 : _GEN_3151; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3668 = ~quene ? tag_1_59 : _GEN_3152; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3669 = ~quene ? tag_1_60 : _GEN_3153; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3670 = ~quene ? tag_1_61 : _GEN_3154; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3671 = ~quene ? tag_1_62 : _GEN_3155; // @[d_cache.scala 154:34 23:24]
  wire [31:0] _GEN_3672 = ~quene ? tag_1_63 : _GEN_3156; // @[d_cache.scala 154:34 23:24]
  wire  _GEN_3673 = ~quene ? dirty_1_0 : _GEN_3157; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3674 = ~quene ? dirty_1_1 : _GEN_3158; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3675 = ~quene ? dirty_1_2 : _GEN_3159; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3676 = ~quene ? dirty_1_3 : _GEN_3160; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3677 = ~quene ? dirty_1_4 : _GEN_3161; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3678 = ~quene ? dirty_1_5 : _GEN_3162; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3679 = ~quene ? dirty_1_6 : _GEN_3163; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3680 = ~quene ? dirty_1_7 : _GEN_3164; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3681 = ~quene ? dirty_1_8 : _GEN_3165; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3682 = ~quene ? dirty_1_9 : _GEN_3166; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3683 = ~quene ? dirty_1_10 : _GEN_3167; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3684 = ~quene ? dirty_1_11 : _GEN_3168; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3685 = ~quene ? dirty_1_12 : _GEN_3169; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3686 = ~quene ? dirty_1_13 : _GEN_3170; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3687 = ~quene ? dirty_1_14 : _GEN_3171; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3688 = ~quene ? dirty_1_15 : _GEN_3172; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3689 = ~quene ? dirty_1_16 : _GEN_3173; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3690 = ~quene ? dirty_1_17 : _GEN_3174; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3691 = ~quene ? dirty_1_18 : _GEN_3175; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3692 = ~quene ? dirty_1_19 : _GEN_3176; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3693 = ~quene ? dirty_1_20 : _GEN_3177; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3694 = ~quene ? dirty_1_21 : _GEN_3178; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3695 = ~quene ? dirty_1_22 : _GEN_3179; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3696 = ~quene ? dirty_1_23 : _GEN_3180; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3697 = ~quene ? dirty_1_24 : _GEN_3181; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3698 = ~quene ? dirty_1_25 : _GEN_3182; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3699 = ~quene ? dirty_1_26 : _GEN_3183; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3700 = ~quene ? dirty_1_27 : _GEN_3184; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3701 = ~quene ? dirty_1_28 : _GEN_3185; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3702 = ~quene ? dirty_1_29 : _GEN_3186; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3703 = ~quene ? dirty_1_30 : _GEN_3187; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3704 = ~quene ? dirty_1_31 : _GEN_3188; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3705 = ~quene ? dirty_1_32 : _GEN_3189; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3706 = ~quene ? dirty_1_33 : _GEN_3190; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3707 = ~quene ? dirty_1_34 : _GEN_3191; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3708 = ~quene ? dirty_1_35 : _GEN_3192; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3709 = ~quene ? dirty_1_36 : _GEN_3193; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3710 = ~quene ? dirty_1_37 : _GEN_3194; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3711 = ~quene ? dirty_1_38 : _GEN_3195; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3712 = ~quene ? dirty_1_39 : _GEN_3196; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3713 = ~quene ? dirty_1_40 : _GEN_3197; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3714 = ~quene ? dirty_1_41 : _GEN_3198; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3715 = ~quene ? dirty_1_42 : _GEN_3199; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3716 = ~quene ? dirty_1_43 : _GEN_3200; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3717 = ~quene ? dirty_1_44 : _GEN_3201; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3718 = ~quene ? dirty_1_45 : _GEN_3202; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3719 = ~quene ? dirty_1_46 : _GEN_3203; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3720 = ~quene ? dirty_1_47 : _GEN_3204; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3721 = ~quene ? dirty_1_48 : _GEN_3205; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3722 = ~quene ? dirty_1_49 : _GEN_3206; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3723 = ~quene ? dirty_1_50 : _GEN_3207; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3724 = ~quene ? dirty_1_51 : _GEN_3208; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3725 = ~quene ? dirty_1_52 : _GEN_3209; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3726 = ~quene ? dirty_1_53 : _GEN_3210; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3727 = ~quene ? dirty_1_54 : _GEN_3211; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3728 = ~quene ? dirty_1_55 : _GEN_3212; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3729 = ~quene ? dirty_1_56 : _GEN_3213; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3730 = ~quene ? dirty_1_57 : _GEN_3214; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3731 = ~quene ? dirty_1_58 : _GEN_3215; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3732 = ~quene ? dirty_1_59 : _GEN_3216; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3733 = ~quene ? dirty_1_60 : _GEN_3217; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3734 = ~quene ? dirty_1_61 : _GEN_3218; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3735 = ~quene ? dirty_1_62 : _GEN_3219; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3736 = ~quene ? dirty_1_63 : _GEN_3220; // @[d_cache.scala 154:34 27:26]
  wire  _GEN_3737 = ~quene ? valid_1_0 : _GEN_3221; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3738 = ~quene ? valid_1_1 : _GEN_3222; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3739 = ~quene ? valid_1_2 : _GEN_3223; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3740 = ~quene ? valid_1_3 : _GEN_3224; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3741 = ~quene ? valid_1_4 : _GEN_3225; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3742 = ~quene ? valid_1_5 : _GEN_3226; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3743 = ~quene ? valid_1_6 : _GEN_3227; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3744 = ~quene ? valid_1_7 : _GEN_3228; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3745 = ~quene ? valid_1_8 : _GEN_3229; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3746 = ~quene ? valid_1_9 : _GEN_3230; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3747 = ~quene ? valid_1_10 : _GEN_3231; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3748 = ~quene ? valid_1_11 : _GEN_3232; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3749 = ~quene ? valid_1_12 : _GEN_3233; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3750 = ~quene ? valid_1_13 : _GEN_3234; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3751 = ~quene ? valid_1_14 : _GEN_3235; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3752 = ~quene ? valid_1_15 : _GEN_3236; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3753 = ~quene ? valid_1_16 : _GEN_3237; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3754 = ~quene ? valid_1_17 : _GEN_3238; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3755 = ~quene ? valid_1_18 : _GEN_3239; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3756 = ~quene ? valid_1_19 : _GEN_3240; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3757 = ~quene ? valid_1_20 : _GEN_3241; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3758 = ~quene ? valid_1_21 : _GEN_3242; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3759 = ~quene ? valid_1_22 : _GEN_3243; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3760 = ~quene ? valid_1_23 : _GEN_3244; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3761 = ~quene ? valid_1_24 : _GEN_3245; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3762 = ~quene ? valid_1_25 : _GEN_3246; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3763 = ~quene ? valid_1_26 : _GEN_3247; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3764 = ~quene ? valid_1_27 : _GEN_3248; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3765 = ~quene ? valid_1_28 : _GEN_3249; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3766 = ~quene ? valid_1_29 : _GEN_3250; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3767 = ~quene ? valid_1_30 : _GEN_3251; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3768 = ~quene ? valid_1_31 : _GEN_3252; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3769 = ~quene ? valid_1_32 : _GEN_3253; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3770 = ~quene ? valid_1_33 : _GEN_3254; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3771 = ~quene ? valid_1_34 : _GEN_3255; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3772 = ~quene ? valid_1_35 : _GEN_3256; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3773 = ~quene ? valid_1_36 : _GEN_3257; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3774 = ~quene ? valid_1_37 : _GEN_3258; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3775 = ~quene ? valid_1_38 : _GEN_3259; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3776 = ~quene ? valid_1_39 : _GEN_3260; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3777 = ~quene ? valid_1_40 : _GEN_3261; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3778 = ~quene ? valid_1_41 : _GEN_3262; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3779 = ~quene ? valid_1_42 : _GEN_3263; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3780 = ~quene ? valid_1_43 : _GEN_3264; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3781 = ~quene ? valid_1_44 : _GEN_3265; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3782 = ~quene ? valid_1_45 : _GEN_3266; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3783 = ~quene ? valid_1_46 : _GEN_3267; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3784 = ~quene ? valid_1_47 : _GEN_3268; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3785 = ~quene ? valid_1_48 : _GEN_3269; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3786 = ~quene ? valid_1_49 : _GEN_3270; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3787 = ~quene ? valid_1_50 : _GEN_3271; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3788 = ~quene ? valid_1_51 : _GEN_3272; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3789 = ~quene ? valid_1_52 : _GEN_3273; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3790 = ~quene ? valid_1_53 : _GEN_3274; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3791 = ~quene ? valid_1_54 : _GEN_3275; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3792 = ~quene ? valid_1_55 : _GEN_3276; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3793 = ~quene ? valid_1_56 : _GEN_3277; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3794 = ~quene ? valid_1_57 : _GEN_3278; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3795 = ~quene ? valid_1_58 : _GEN_3279; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3796 = ~quene ? valid_1_59 : _GEN_3280; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3797 = ~quene ? valid_1_60 : _GEN_3281; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3798 = ~quene ? valid_1_61 : _GEN_3282; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3799 = ~quene ? valid_1_62 : _GEN_3283; // @[d_cache.scala 154:34 25:26]
  wire  _GEN_3800 = ~quene ? valid_1_63 : _GEN_3284; // @[d_cache.scala 154:34 25:26]
  wire [2:0] _GEN_3801 = unuse_way == 2'h2 ? 3'h7 : _GEN_3544; // @[d_cache.scala 147:40 148:23]
  wire [63:0] _GEN_3802 = unuse_way == 2'h2 ? _GEN_1680 : _GEN_3545; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3803 = unuse_way == 2'h2 ? _GEN_1681 : _GEN_3546; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3804 = unuse_way == 2'h2 ? _GEN_1682 : _GEN_3547; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3805 = unuse_way == 2'h2 ? _GEN_1683 : _GEN_3548; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3806 = unuse_way == 2'h2 ? _GEN_1684 : _GEN_3549; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3807 = unuse_way == 2'h2 ? _GEN_1685 : _GEN_3550; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3808 = unuse_way == 2'h2 ? _GEN_1686 : _GEN_3551; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3809 = unuse_way == 2'h2 ? _GEN_1687 : _GEN_3552; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3810 = unuse_way == 2'h2 ? _GEN_1688 : _GEN_3553; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3811 = unuse_way == 2'h2 ? _GEN_1689 : _GEN_3554; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3812 = unuse_way == 2'h2 ? _GEN_1690 : _GEN_3555; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3813 = unuse_way == 2'h2 ? _GEN_1691 : _GEN_3556; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3814 = unuse_way == 2'h2 ? _GEN_1692 : _GEN_3557; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3815 = unuse_way == 2'h2 ? _GEN_1693 : _GEN_3558; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3816 = unuse_way == 2'h2 ? _GEN_1694 : _GEN_3559; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3817 = unuse_way == 2'h2 ? _GEN_1695 : _GEN_3560; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3818 = unuse_way == 2'h2 ? _GEN_1696 : _GEN_3561; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3819 = unuse_way == 2'h2 ? _GEN_1697 : _GEN_3562; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3820 = unuse_way == 2'h2 ? _GEN_1698 : _GEN_3563; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3821 = unuse_way == 2'h2 ? _GEN_1699 : _GEN_3564; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3822 = unuse_way == 2'h2 ? _GEN_1700 : _GEN_3565; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3823 = unuse_way == 2'h2 ? _GEN_1701 : _GEN_3566; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3824 = unuse_way == 2'h2 ? _GEN_1702 : _GEN_3567; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3825 = unuse_way == 2'h2 ? _GEN_1703 : _GEN_3568; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3826 = unuse_way == 2'h2 ? _GEN_1704 : _GEN_3569; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3827 = unuse_way == 2'h2 ? _GEN_1705 : _GEN_3570; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3828 = unuse_way == 2'h2 ? _GEN_1706 : _GEN_3571; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3829 = unuse_way == 2'h2 ? _GEN_1707 : _GEN_3572; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3830 = unuse_way == 2'h2 ? _GEN_1708 : _GEN_3573; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3831 = unuse_way == 2'h2 ? _GEN_1709 : _GEN_3574; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3832 = unuse_way == 2'h2 ? _GEN_1710 : _GEN_3575; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3833 = unuse_way == 2'h2 ? _GEN_1711 : _GEN_3576; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3834 = unuse_way == 2'h2 ? _GEN_1712 : _GEN_3577; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3835 = unuse_way == 2'h2 ? _GEN_1713 : _GEN_3578; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3836 = unuse_way == 2'h2 ? _GEN_1714 : _GEN_3579; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3837 = unuse_way == 2'h2 ? _GEN_1715 : _GEN_3580; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3838 = unuse_way == 2'h2 ? _GEN_1716 : _GEN_3581; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3839 = unuse_way == 2'h2 ? _GEN_1717 : _GEN_3582; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3840 = unuse_way == 2'h2 ? _GEN_1718 : _GEN_3583; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3841 = unuse_way == 2'h2 ? _GEN_1719 : _GEN_3584; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3842 = unuse_way == 2'h2 ? _GEN_1720 : _GEN_3585; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3843 = unuse_way == 2'h2 ? _GEN_1721 : _GEN_3586; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3844 = unuse_way == 2'h2 ? _GEN_1722 : _GEN_3587; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3845 = unuse_way == 2'h2 ? _GEN_1723 : _GEN_3588; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3846 = unuse_way == 2'h2 ? _GEN_1724 : _GEN_3589; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3847 = unuse_way == 2'h2 ? _GEN_1725 : _GEN_3590; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3848 = unuse_way == 2'h2 ? _GEN_1726 : _GEN_3591; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3849 = unuse_way == 2'h2 ? _GEN_1727 : _GEN_3592; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3850 = unuse_way == 2'h2 ? _GEN_1728 : _GEN_3593; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3851 = unuse_way == 2'h2 ? _GEN_1729 : _GEN_3594; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3852 = unuse_way == 2'h2 ? _GEN_1730 : _GEN_3595; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3853 = unuse_way == 2'h2 ? _GEN_1731 : _GEN_3596; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3854 = unuse_way == 2'h2 ? _GEN_1732 : _GEN_3597; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3855 = unuse_way == 2'h2 ? _GEN_1733 : _GEN_3598; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3856 = unuse_way == 2'h2 ? _GEN_1734 : _GEN_3599; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3857 = unuse_way == 2'h2 ? _GEN_1735 : _GEN_3600; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3858 = unuse_way == 2'h2 ? _GEN_1736 : _GEN_3601; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3859 = unuse_way == 2'h2 ? _GEN_1737 : _GEN_3602; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3860 = unuse_way == 2'h2 ? _GEN_1738 : _GEN_3603; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3861 = unuse_way == 2'h2 ? _GEN_1739 : _GEN_3604; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3862 = unuse_way == 2'h2 ? _GEN_1740 : _GEN_3605; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3863 = unuse_way == 2'h2 ? _GEN_1741 : _GEN_3606; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3864 = unuse_way == 2'h2 ? _GEN_1742 : _GEN_3607; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3865 = unuse_way == 2'h2 ? _GEN_1743 : _GEN_3608; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3866 = unuse_way == 2'h2 ? _GEN_1744 : _GEN_3609; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3867 = unuse_way == 2'h2 ? _GEN_1745 : _GEN_3610; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3868 = unuse_way == 2'h2 ? _GEN_1746 : _GEN_3611; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3869 = unuse_way == 2'h2 ? _GEN_1747 : _GEN_3612; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3870 = unuse_way == 2'h2 ? _GEN_1748 : _GEN_3613; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3871 = unuse_way == 2'h2 ? _GEN_1749 : _GEN_3614; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3872 = unuse_way == 2'h2 ? _GEN_1750 : _GEN_3615; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3873 = unuse_way == 2'h2 ? _GEN_1751 : _GEN_3616; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3874 = unuse_way == 2'h2 ? _GEN_1752 : _GEN_3617; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3875 = unuse_way == 2'h2 ? _GEN_1753 : _GEN_3618; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3876 = unuse_way == 2'h2 ? _GEN_1754 : _GEN_3619; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3877 = unuse_way == 2'h2 ? _GEN_1755 : _GEN_3620; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3878 = unuse_way == 2'h2 ? _GEN_1756 : _GEN_3621; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3879 = unuse_way == 2'h2 ? _GEN_1757 : _GEN_3622; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3880 = unuse_way == 2'h2 ? _GEN_1758 : _GEN_3623; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3881 = unuse_way == 2'h2 ? _GEN_1759 : _GEN_3624; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3882 = unuse_way == 2'h2 ? _GEN_1760 : _GEN_3625; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3883 = unuse_way == 2'h2 ? _GEN_1761 : _GEN_3626; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3884 = unuse_way == 2'h2 ? _GEN_1762 : _GEN_3627; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3885 = unuse_way == 2'h2 ? _GEN_1763 : _GEN_3628; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3886 = unuse_way == 2'h2 ? _GEN_1764 : _GEN_3629; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3887 = unuse_way == 2'h2 ? _GEN_1765 : _GEN_3630; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3888 = unuse_way == 2'h2 ? _GEN_1766 : _GEN_3631; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3889 = unuse_way == 2'h2 ? _GEN_1767 : _GEN_3632; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3890 = unuse_way == 2'h2 ? _GEN_1768 : _GEN_3633; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3891 = unuse_way == 2'h2 ? _GEN_1769 : _GEN_3634; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3892 = unuse_way == 2'h2 ? _GEN_1770 : _GEN_3635; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3893 = unuse_way == 2'h2 ? _GEN_1771 : _GEN_3636; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3894 = unuse_way == 2'h2 ? _GEN_1772 : _GEN_3637; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3895 = unuse_way == 2'h2 ? _GEN_1773 : _GEN_3638; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3896 = unuse_way == 2'h2 ? _GEN_1774 : _GEN_3639; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3897 = unuse_way == 2'h2 ? _GEN_1775 : _GEN_3640; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3898 = unuse_way == 2'h2 ? _GEN_1776 : _GEN_3641; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3899 = unuse_way == 2'h2 ? _GEN_1777 : _GEN_3642; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3900 = unuse_way == 2'h2 ? _GEN_1778 : _GEN_3643; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3901 = unuse_way == 2'h2 ? _GEN_1779 : _GEN_3644; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3902 = unuse_way == 2'h2 ? _GEN_1780 : _GEN_3645; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3903 = unuse_way == 2'h2 ? _GEN_1781 : _GEN_3646; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3904 = unuse_way == 2'h2 ? _GEN_1782 : _GEN_3647; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3905 = unuse_way == 2'h2 ? _GEN_1783 : _GEN_3648; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3906 = unuse_way == 2'h2 ? _GEN_1784 : _GEN_3649; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3907 = unuse_way == 2'h2 ? _GEN_1785 : _GEN_3650; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3908 = unuse_way == 2'h2 ? _GEN_1786 : _GEN_3651; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3909 = unuse_way == 2'h2 ? _GEN_1787 : _GEN_3652; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3910 = unuse_way == 2'h2 ? _GEN_1788 : _GEN_3653; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3911 = unuse_way == 2'h2 ? _GEN_1789 : _GEN_3654; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3912 = unuse_way == 2'h2 ? _GEN_1790 : _GEN_3655; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3913 = unuse_way == 2'h2 ? _GEN_1791 : _GEN_3656; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3914 = unuse_way == 2'h2 ? _GEN_1792 : _GEN_3657; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3915 = unuse_way == 2'h2 ? _GEN_1793 : _GEN_3658; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3916 = unuse_way == 2'h2 ? _GEN_1794 : _GEN_3659; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3917 = unuse_way == 2'h2 ? _GEN_1795 : _GEN_3660; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3918 = unuse_way == 2'h2 ? _GEN_1796 : _GEN_3661; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3919 = unuse_way == 2'h2 ? _GEN_1797 : _GEN_3662; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3920 = unuse_way == 2'h2 ? _GEN_1798 : _GEN_3663; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3921 = unuse_way == 2'h2 ? _GEN_1799 : _GEN_3664; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3922 = unuse_way == 2'h2 ? _GEN_1800 : _GEN_3665; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3923 = unuse_way == 2'h2 ? _GEN_1801 : _GEN_3666; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3924 = unuse_way == 2'h2 ? _GEN_1802 : _GEN_3667; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3925 = unuse_way == 2'h2 ? _GEN_1803 : _GEN_3668; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3926 = unuse_way == 2'h2 ? _GEN_1804 : _GEN_3669; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3927 = unuse_way == 2'h2 ? _GEN_1805 : _GEN_3670; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3928 = unuse_way == 2'h2 ? _GEN_1806 : _GEN_3671; // @[d_cache.scala 147:40]
  wire [31:0] _GEN_3929 = unuse_way == 2'h2 ? _GEN_1807 : _GEN_3672; // @[d_cache.scala 147:40]
  wire  _GEN_3930 = unuse_way == 2'h2 ? _GEN_777 : _GEN_3737; // @[d_cache.scala 147:40]
  wire  _GEN_3931 = unuse_way == 2'h2 ? _GEN_778 : _GEN_3738; // @[d_cache.scala 147:40]
  wire  _GEN_3932 = unuse_way == 2'h2 ? _GEN_779 : _GEN_3739; // @[d_cache.scala 147:40]
  wire  _GEN_3933 = unuse_way == 2'h2 ? _GEN_780 : _GEN_3740; // @[d_cache.scala 147:40]
  wire  _GEN_3934 = unuse_way == 2'h2 ? _GEN_781 : _GEN_3741; // @[d_cache.scala 147:40]
  wire  _GEN_3935 = unuse_way == 2'h2 ? _GEN_782 : _GEN_3742; // @[d_cache.scala 147:40]
  wire  _GEN_3936 = unuse_way == 2'h2 ? _GEN_783 : _GEN_3743; // @[d_cache.scala 147:40]
  wire  _GEN_3937 = unuse_way == 2'h2 ? _GEN_784 : _GEN_3744; // @[d_cache.scala 147:40]
  wire  _GEN_3938 = unuse_way == 2'h2 ? _GEN_785 : _GEN_3745; // @[d_cache.scala 147:40]
  wire  _GEN_3939 = unuse_way == 2'h2 ? _GEN_786 : _GEN_3746; // @[d_cache.scala 147:40]
  wire  _GEN_3940 = unuse_way == 2'h2 ? _GEN_787 : _GEN_3747; // @[d_cache.scala 147:40]
  wire  _GEN_3941 = unuse_way == 2'h2 ? _GEN_788 : _GEN_3748; // @[d_cache.scala 147:40]
  wire  _GEN_3942 = unuse_way == 2'h2 ? _GEN_789 : _GEN_3749; // @[d_cache.scala 147:40]
  wire  _GEN_3943 = unuse_way == 2'h2 ? _GEN_790 : _GEN_3750; // @[d_cache.scala 147:40]
  wire  _GEN_3944 = unuse_way == 2'h2 ? _GEN_791 : _GEN_3751; // @[d_cache.scala 147:40]
  wire  _GEN_3945 = unuse_way == 2'h2 ? _GEN_792 : _GEN_3752; // @[d_cache.scala 147:40]
  wire  _GEN_3946 = unuse_way == 2'h2 ? _GEN_793 : _GEN_3753; // @[d_cache.scala 147:40]
  wire  _GEN_3947 = unuse_way == 2'h2 ? _GEN_794 : _GEN_3754; // @[d_cache.scala 147:40]
  wire  _GEN_3948 = unuse_way == 2'h2 ? _GEN_795 : _GEN_3755; // @[d_cache.scala 147:40]
  wire  _GEN_3949 = unuse_way == 2'h2 ? _GEN_796 : _GEN_3756; // @[d_cache.scala 147:40]
  wire  _GEN_3950 = unuse_way == 2'h2 ? _GEN_797 : _GEN_3757; // @[d_cache.scala 147:40]
  wire  _GEN_3951 = unuse_way == 2'h2 ? _GEN_798 : _GEN_3758; // @[d_cache.scala 147:40]
  wire  _GEN_3952 = unuse_way == 2'h2 ? _GEN_799 : _GEN_3759; // @[d_cache.scala 147:40]
  wire  _GEN_3953 = unuse_way == 2'h2 ? _GEN_800 : _GEN_3760; // @[d_cache.scala 147:40]
  wire  _GEN_3954 = unuse_way == 2'h2 ? _GEN_801 : _GEN_3761; // @[d_cache.scala 147:40]
  wire  _GEN_3955 = unuse_way == 2'h2 ? _GEN_802 : _GEN_3762; // @[d_cache.scala 147:40]
  wire  _GEN_3956 = unuse_way == 2'h2 ? _GEN_803 : _GEN_3763; // @[d_cache.scala 147:40]
  wire  _GEN_3957 = unuse_way == 2'h2 ? _GEN_804 : _GEN_3764; // @[d_cache.scala 147:40]
  wire  _GEN_3958 = unuse_way == 2'h2 ? _GEN_805 : _GEN_3765; // @[d_cache.scala 147:40]
  wire  _GEN_3959 = unuse_way == 2'h2 ? _GEN_806 : _GEN_3766; // @[d_cache.scala 147:40]
  wire  _GEN_3960 = unuse_way == 2'h2 ? _GEN_807 : _GEN_3767; // @[d_cache.scala 147:40]
  wire  _GEN_3961 = unuse_way == 2'h2 ? _GEN_808 : _GEN_3768; // @[d_cache.scala 147:40]
  wire  _GEN_3962 = unuse_way == 2'h2 ? _GEN_809 : _GEN_3769; // @[d_cache.scala 147:40]
  wire  _GEN_3963 = unuse_way == 2'h2 ? _GEN_810 : _GEN_3770; // @[d_cache.scala 147:40]
  wire  _GEN_3964 = unuse_way == 2'h2 ? _GEN_811 : _GEN_3771; // @[d_cache.scala 147:40]
  wire  _GEN_3965 = unuse_way == 2'h2 ? _GEN_812 : _GEN_3772; // @[d_cache.scala 147:40]
  wire  _GEN_3966 = unuse_way == 2'h2 ? _GEN_813 : _GEN_3773; // @[d_cache.scala 147:40]
  wire  _GEN_3967 = unuse_way == 2'h2 ? _GEN_814 : _GEN_3774; // @[d_cache.scala 147:40]
  wire  _GEN_3968 = unuse_way == 2'h2 ? _GEN_815 : _GEN_3775; // @[d_cache.scala 147:40]
  wire  _GEN_3969 = unuse_way == 2'h2 ? _GEN_816 : _GEN_3776; // @[d_cache.scala 147:40]
  wire  _GEN_3970 = unuse_way == 2'h2 ? _GEN_817 : _GEN_3777; // @[d_cache.scala 147:40]
  wire  _GEN_3971 = unuse_way == 2'h2 ? _GEN_818 : _GEN_3778; // @[d_cache.scala 147:40]
  wire  _GEN_3972 = unuse_way == 2'h2 ? _GEN_819 : _GEN_3779; // @[d_cache.scala 147:40]
  wire  _GEN_3973 = unuse_way == 2'h2 ? _GEN_820 : _GEN_3780; // @[d_cache.scala 147:40]
  wire  _GEN_3974 = unuse_way == 2'h2 ? _GEN_821 : _GEN_3781; // @[d_cache.scala 147:40]
  wire  _GEN_3975 = unuse_way == 2'h2 ? _GEN_822 : _GEN_3782; // @[d_cache.scala 147:40]
  wire  _GEN_3976 = unuse_way == 2'h2 ? _GEN_823 : _GEN_3783; // @[d_cache.scala 147:40]
  wire  _GEN_3977 = unuse_way == 2'h2 ? _GEN_824 : _GEN_3784; // @[d_cache.scala 147:40]
  wire  _GEN_3978 = unuse_way == 2'h2 ? _GEN_825 : _GEN_3785; // @[d_cache.scala 147:40]
  wire  _GEN_3979 = unuse_way == 2'h2 ? _GEN_826 : _GEN_3786; // @[d_cache.scala 147:40]
  wire  _GEN_3980 = unuse_way == 2'h2 ? _GEN_827 : _GEN_3787; // @[d_cache.scala 147:40]
  wire  _GEN_3981 = unuse_way == 2'h2 ? _GEN_828 : _GEN_3788; // @[d_cache.scala 147:40]
  wire  _GEN_3982 = unuse_way == 2'h2 ? _GEN_829 : _GEN_3789; // @[d_cache.scala 147:40]
  wire  _GEN_3983 = unuse_way == 2'h2 ? _GEN_830 : _GEN_3790; // @[d_cache.scala 147:40]
  wire  _GEN_3984 = unuse_way == 2'h2 ? _GEN_831 : _GEN_3791; // @[d_cache.scala 147:40]
  wire  _GEN_3985 = unuse_way == 2'h2 ? _GEN_832 : _GEN_3792; // @[d_cache.scala 147:40]
  wire  _GEN_3986 = unuse_way == 2'h2 ? _GEN_833 : _GEN_3793; // @[d_cache.scala 147:40]
  wire  _GEN_3987 = unuse_way == 2'h2 ? _GEN_834 : _GEN_3794; // @[d_cache.scala 147:40]
  wire  _GEN_3988 = unuse_way == 2'h2 ? _GEN_835 : _GEN_3795; // @[d_cache.scala 147:40]
  wire  _GEN_3989 = unuse_way == 2'h2 ? _GEN_836 : _GEN_3796; // @[d_cache.scala 147:40]
  wire  _GEN_3990 = unuse_way == 2'h2 ? _GEN_837 : _GEN_3797; // @[d_cache.scala 147:40]
  wire  _GEN_3991 = unuse_way == 2'h2 ? _GEN_838 : _GEN_3798; // @[d_cache.scala 147:40]
  wire  _GEN_3992 = unuse_way == 2'h2 ? _GEN_839 : _GEN_3799; // @[d_cache.scala 147:40]
  wire  _GEN_3993 = unuse_way == 2'h2 ? _GEN_840 : _GEN_3800; // @[d_cache.scala 147:40]
  wire [63:0] _GEN_3994 = unuse_way == 2'h2 ? write_back_data : _GEN_3286; // @[d_cache.scala 147:40 31:34]
  wire [40:0] _GEN_3995 = unuse_way == 2'h2 ? {{9'd0}, write_back_addr} : _GEN_3287; // @[d_cache.scala 147:40 32:34]
  wire [63:0] _GEN_3996 = unuse_way == 2'h2 ? ram_0_0 : _GEN_3288; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_3997 = unuse_way == 2'h2 ? ram_0_1 : _GEN_3289; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_3998 = unuse_way == 2'h2 ? ram_0_2 : _GEN_3290; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_3999 = unuse_way == 2'h2 ? ram_0_3 : _GEN_3291; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4000 = unuse_way == 2'h2 ? ram_0_4 : _GEN_3292; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4001 = unuse_way == 2'h2 ? ram_0_5 : _GEN_3293; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4002 = unuse_way == 2'h2 ? ram_0_6 : _GEN_3294; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4003 = unuse_way == 2'h2 ? ram_0_7 : _GEN_3295; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4004 = unuse_way == 2'h2 ? ram_0_8 : _GEN_3296; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4005 = unuse_way == 2'h2 ? ram_0_9 : _GEN_3297; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4006 = unuse_way == 2'h2 ? ram_0_10 : _GEN_3298; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4007 = unuse_way == 2'h2 ? ram_0_11 : _GEN_3299; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4008 = unuse_way == 2'h2 ? ram_0_12 : _GEN_3300; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4009 = unuse_way == 2'h2 ? ram_0_13 : _GEN_3301; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4010 = unuse_way == 2'h2 ? ram_0_14 : _GEN_3302; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4011 = unuse_way == 2'h2 ? ram_0_15 : _GEN_3303; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4012 = unuse_way == 2'h2 ? ram_0_16 : _GEN_3304; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4013 = unuse_way == 2'h2 ? ram_0_17 : _GEN_3305; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4014 = unuse_way == 2'h2 ? ram_0_18 : _GEN_3306; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4015 = unuse_way == 2'h2 ? ram_0_19 : _GEN_3307; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4016 = unuse_way == 2'h2 ? ram_0_20 : _GEN_3308; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4017 = unuse_way == 2'h2 ? ram_0_21 : _GEN_3309; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4018 = unuse_way == 2'h2 ? ram_0_22 : _GEN_3310; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4019 = unuse_way == 2'h2 ? ram_0_23 : _GEN_3311; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4020 = unuse_way == 2'h2 ? ram_0_24 : _GEN_3312; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4021 = unuse_way == 2'h2 ? ram_0_25 : _GEN_3313; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4022 = unuse_way == 2'h2 ? ram_0_26 : _GEN_3314; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4023 = unuse_way == 2'h2 ? ram_0_27 : _GEN_3315; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4024 = unuse_way == 2'h2 ? ram_0_28 : _GEN_3316; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4025 = unuse_way == 2'h2 ? ram_0_29 : _GEN_3317; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4026 = unuse_way == 2'h2 ? ram_0_30 : _GEN_3318; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4027 = unuse_way == 2'h2 ? ram_0_31 : _GEN_3319; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4028 = unuse_way == 2'h2 ? ram_0_32 : _GEN_3320; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4029 = unuse_way == 2'h2 ? ram_0_33 : _GEN_3321; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4030 = unuse_way == 2'h2 ? ram_0_34 : _GEN_3322; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4031 = unuse_way == 2'h2 ? ram_0_35 : _GEN_3323; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4032 = unuse_way == 2'h2 ? ram_0_36 : _GEN_3324; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4033 = unuse_way == 2'h2 ? ram_0_37 : _GEN_3325; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4034 = unuse_way == 2'h2 ? ram_0_38 : _GEN_3326; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4035 = unuse_way == 2'h2 ? ram_0_39 : _GEN_3327; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4036 = unuse_way == 2'h2 ? ram_0_40 : _GEN_3328; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4037 = unuse_way == 2'h2 ? ram_0_41 : _GEN_3329; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4038 = unuse_way == 2'h2 ? ram_0_42 : _GEN_3330; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4039 = unuse_way == 2'h2 ? ram_0_43 : _GEN_3331; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4040 = unuse_way == 2'h2 ? ram_0_44 : _GEN_3332; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4041 = unuse_way == 2'h2 ? ram_0_45 : _GEN_3333; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4042 = unuse_way == 2'h2 ? ram_0_46 : _GEN_3334; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4043 = unuse_way == 2'h2 ? ram_0_47 : _GEN_3335; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4044 = unuse_way == 2'h2 ? ram_0_48 : _GEN_3336; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4045 = unuse_way == 2'h2 ? ram_0_49 : _GEN_3337; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4046 = unuse_way == 2'h2 ? ram_0_50 : _GEN_3338; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4047 = unuse_way == 2'h2 ? ram_0_51 : _GEN_3339; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4048 = unuse_way == 2'h2 ? ram_0_52 : _GEN_3340; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4049 = unuse_way == 2'h2 ? ram_0_53 : _GEN_3341; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4050 = unuse_way == 2'h2 ? ram_0_54 : _GEN_3342; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4051 = unuse_way == 2'h2 ? ram_0_55 : _GEN_3343; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4052 = unuse_way == 2'h2 ? ram_0_56 : _GEN_3344; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4053 = unuse_way == 2'h2 ? ram_0_57 : _GEN_3345; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4054 = unuse_way == 2'h2 ? ram_0_58 : _GEN_3346; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4055 = unuse_way == 2'h2 ? ram_0_59 : _GEN_3347; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4056 = unuse_way == 2'h2 ? ram_0_60 : _GEN_3348; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4057 = unuse_way == 2'h2 ? ram_0_61 : _GEN_3349; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4058 = unuse_way == 2'h2 ? ram_0_62 : _GEN_3350; // @[d_cache.scala 147:40 18:24]
  wire [63:0] _GEN_4059 = unuse_way == 2'h2 ? ram_0_63 : _GEN_3351; // @[d_cache.scala 147:40 18:24]
  wire [31:0] _GEN_4060 = unuse_way == 2'h2 ? tag_0_0 : _GEN_3352; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4061 = unuse_way == 2'h2 ? tag_0_1 : _GEN_3353; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4062 = unuse_way == 2'h2 ? tag_0_2 : _GEN_3354; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4063 = unuse_way == 2'h2 ? tag_0_3 : _GEN_3355; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4064 = unuse_way == 2'h2 ? tag_0_4 : _GEN_3356; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4065 = unuse_way == 2'h2 ? tag_0_5 : _GEN_3357; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4066 = unuse_way == 2'h2 ? tag_0_6 : _GEN_3358; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4067 = unuse_way == 2'h2 ? tag_0_7 : _GEN_3359; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4068 = unuse_way == 2'h2 ? tag_0_8 : _GEN_3360; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4069 = unuse_way == 2'h2 ? tag_0_9 : _GEN_3361; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4070 = unuse_way == 2'h2 ? tag_0_10 : _GEN_3362; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4071 = unuse_way == 2'h2 ? tag_0_11 : _GEN_3363; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4072 = unuse_way == 2'h2 ? tag_0_12 : _GEN_3364; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4073 = unuse_way == 2'h2 ? tag_0_13 : _GEN_3365; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4074 = unuse_way == 2'h2 ? tag_0_14 : _GEN_3366; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4075 = unuse_way == 2'h2 ? tag_0_15 : _GEN_3367; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4076 = unuse_way == 2'h2 ? tag_0_16 : _GEN_3368; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4077 = unuse_way == 2'h2 ? tag_0_17 : _GEN_3369; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4078 = unuse_way == 2'h2 ? tag_0_18 : _GEN_3370; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4079 = unuse_way == 2'h2 ? tag_0_19 : _GEN_3371; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4080 = unuse_way == 2'h2 ? tag_0_20 : _GEN_3372; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4081 = unuse_way == 2'h2 ? tag_0_21 : _GEN_3373; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4082 = unuse_way == 2'h2 ? tag_0_22 : _GEN_3374; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4083 = unuse_way == 2'h2 ? tag_0_23 : _GEN_3375; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4084 = unuse_way == 2'h2 ? tag_0_24 : _GEN_3376; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4085 = unuse_way == 2'h2 ? tag_0_25 : _GEN_3377; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4086 = unuse_way == 2'h2 ? tag_0_26 : _GEN_3378; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4087 = unuse_way == 2'h2 ? tag_0_27 : _GEN_3379; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4088 = unuse_way == 2'h2 ? tag_0_28 : _GEN_3380; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4089 = unuse_way == 2'h2 ? tag_0_29 : _GEN_3381; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4090 = unuse_way == 2'h2 ? tag_0_30 : _GEN_3382; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4091 = unuse_way == 2'h2 ? tag_0_31 : _GEN_3383; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4092 = unuse_way == 2'h2 ? tag_0_32 : _GEN_3384; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4093 = unuse_way == 2'h2 ? tag_0_33 : _GEN_3385; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4094 = unuse_way == 2'h2 ? tag_0_34 : _GEN_3386; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4095 = unuse_way == 2'h2 ? tag_0_35 : _GEN_3387; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4096 = unuse_way == 2'h2 ? tag_0_36 : _GEN_3388; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4097 = unuse_way == 2'h2 ? tag_0_37 : _GEN_3389; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4098 = unuse_way == 2'h2 ? tag_0_38 : _GEN_3390; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4099 = unuse_way == 2'h2 ? tag_0_39 : _GEN_3391; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4100 = unuse_way == 2'h2 ? tag_0_40 : _GEN_3392; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4101 = unuse_way == 2'h2 ? tag_0_41 : _GEN_3393; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4102 = unuse_way == 2'h2 ? tag_0_42 : _GEN_3394; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4103 = unuse_way == 2'h2 ? tag_0_43 : _GEN_3395; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4104 = unuse_way == 2'h2 ? tag_0_44 : _GEN_3396; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4105 = unuse_way == 2'h2 ? tag_0_45 : _GEN_3397; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4106 = unuse_way == 2'h2 ? tag_0_46 : _GEN_3398; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4107 = unuse_way == 2'h2 ? tag_0_47 : _GEN_3399; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4108 = unuse_way == 2'h2 ? tag_0_48 : _GEN_3400; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4109 = unuse_way == 2'h2 ? tag_0_49 : _GEN_3401; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4110 = unuse_way == 2'h2 ? tag_0_50 : _GEN_3402; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4111 = unuse_way == 2'h2 ? tag_0_51 : _GEN_3403; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4112 = unuse_way == 2'h2 ? tag_0_52 : _GEN_3404; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4113 = unuse_way == 2'h2 ? tag_0_53 : _GEN_3405; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4114 = unuse_way == 2'h2 ? tag_0_54 : _GEN_3406; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4115 = unuse_way == 2'h2 ? tag_0_55 : _GEN_3407; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4116 = unuse_way == 2'h2 ? tag_0_56 : _GEN_3408; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4117 = unuse_way == 2'h2 ? tag_0_57 : _GEN_3409; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4118 = unuse_way == 2'h2 ? tag_0_58 : _GEN_3410; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4119 = unuse_way == 2'h2 ? tag_0_59 : _GEN_3411; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4120 = unuse_way == 2'h2 ? tag_0_60 : _GEN_3412; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4121 = unuse_way == 2'h2 ? tag_0_61 : _GEN_3413; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4122 = unuse_way == 2'h2 ? tag_0_62 : _GEN_3414; // @[d_cache.scala 147:40 22:24]
  wire [31:0] _GEN_4123 = unuse_way == 2'h2 ? tag_0_63 : _GEN_3415; // @[d_cache.scala 147:40 22:24]
  wire  _GEN_4124 = unuse_way == 2'h2 ? dirty_0_0 : _GEN_3416; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4125 = unuse_way == 2'h2 ? dirty_0_1 : _GEN_3417; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4126 = unuse_way == 2'h2 ? dirty_0_2 : _GEN_3418; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4127 = unuse_way == 2'h2 ? dirty_0_3 : _GEN_3419; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4128 = unuse_way == 2'h2 ? dirty_0_4 : _GEN_3420; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4129 = unuse_way == 2'h2 ? dirty_0_5 : _GEN_3421; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4130 = unuse_way == 2'h2 ? dirty_0_6 : _GEN_3422; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4131 = unuse_way == 2'h2 ? dirty_0_7 : _GEN_3423; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4132 = unuse_way == 2'h2 ? dirty_0_8 : _GEN_3424; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4133 = unuse_way == 2'h2 ? dirty_0_9 : _GEN_3425; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4134 = unuse_way == 2'h2 ? dirty_0_10 : _GEN_3426; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4135 = unuse_way == 2'h2 ? dirty_0_11 : _GEN_3427; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4136 = unuse_way == 2'h2 ? dirty_0_12 : _GEN_3428; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4137 = unuse_way == 2'h2 ? dirty_0_13 : _GEN_3429; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4138 = unuse_way == 2'h2 ? dirty_0_14 : _GEN_3430; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4139 = unuse_way == 2'h2 ? dirty_0_15 : _GEN_3431; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4140 = unuse_way == 2'h2 ? dirty_0_16 : _GEN_3432; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4141 = unuse_way == 2'h2 ? dirty_0_17 : _GEN_3433; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4142 = unuse_way == 2'h2 ? dirty_0_18 : _GEN_3434; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4143 = unuse_way == 2'h2 ? dirty_0_19 : _GEN_3435; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4144 = unuse_way == 2'h2 ? dirty_0_20 : _GEN_3436; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4145 = unuse_way == 2'h2 ? dirty_0_21 : _GEN_3437; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4146 = unuse_way == 2'h2 ? dirty_0_22 : _GEN_3438; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4147 = unuse_way == 2'h2 ? dirty_0_23 : _GEN_3439; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4148 = unuse_way == 2'h2 ? dirty_0_24 : _GEN_3440; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4149 = unuse_way == 2'h2 ? dirty_0_25 : _GEN_3441; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4150 = unuse_way == 2'h2 ? dirty_0_26 : _GEN_3442; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4151 = unuse_way == 2'h2 ? dirty_0_27 : _GEN_3443; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4152 = unuse_way == 2'h2 ? dirty_0_28 : _GEN_3444; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4153 = unuse_way == 2'h2 ? dirty_0_29 : _GEN_3445; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4154 = unuse_way == 2'h2 ? dirty_0_30 : _GEN_3446; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4155 = unuse_way == 2'h2 ? dirty_0_31 : _GEN_3447; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4156 = unuse_way == 2'h2 ? dirty_0_32 : _GEN_3448; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4157 = unuse_way == 2'h2 ? dirty_0_33 : _GEN_3449; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4158 = unuse_way == 2'h2 ? dirty_0_34 : _GEN_3450; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4159 = unuse_way == 2'h2 ? dirty_0_35 : _GEN_3451; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4160 = unuse_way == 2'h2 ? dirty_0_36 : _GEN_3452; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4161 = unuse_way == 2'h2 ? dirty_0_37 : _GEN_3453; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4162 = unuse_way == 2'h2 ? dirty_0_38 : _GEN_3454; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4163 = unuse_way == 2'h2 ? dirty_0_39 : _GEN_3455; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4164 = unuse_way == 2'h2 ? dirty_0_40 : _GEN_3456; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4165 = unuse_way == 2'h2 ? dirty_0_41 : _GEN_3457; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4166 = unuse_way == 2'h2 ? dirty_0_42 : _GEN_3458; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4167 = unuse_way == 2'h2 ? dirty_0_43 : _GEN_3459; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4168 = unuse_way == 2'h2 ? dirty_0_44 : _GEN_3460; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4169 = unuse_way == 2'h2 ? dirty_0_45 : _GEN_3461; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4170 = unuse_way == 2'h2 ? dirty_0_46 : _GEN_3462; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4171 = unuse_way == 2'h2 ? dirty_0_47 : _GEN_3463; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4172 = unuse_way == 2'h2 ? dirty_0_48 : _GEN_3464; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4173 = unuse_way == 2'h2 ? dirty_0_49 : _GEN_3465; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4174 = unuse_way == 2'h2 ? dirty_0_50 : _GEN_3466; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4175 = unuse_way == 2'h2 ? dirty_0_51 : _GEN_3467; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4176 = unuse_way == 2'h2 ? dirty_0_52 : _GEN_3468; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4177 = unuse_way == 2'h2 ? dirty_0_53 : _GEN_3469; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4178 = unuse_way == 2'h2 ? dirty_0_54 : _GEN_3470; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4179 = unuse_way == 2'h2 ? dirty_0_55 : _GEN_3471; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4180 = unuse_way == 2'h2 ? dirty_0_56 : _GEN_3472; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4181 = unuse_way == 2'h2 ? dirty_0_57 : _GEN_3473; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4182 = unuse_way == 2'h2 ? dirty_0_58 : _GEN_3474; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4183 = unuse_way == 2'h2 ? dirty_0_59 : _GEN_3475; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4184 = unuse_way == 2'h2 ? dirty_0_60 : _GEN_3476; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4185 = unuse_way == 2'h2 ? dirty_0_61 : _GEN_3477; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4186 = unuse_way == 2'h2 ? dirty_0_62 : _GEN_3478; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4187 = unuse_way == 2'h2 ? dirty_0_63 : _GEN_3479; // @[d_cache.scala 147:40 26:26]
  wire  _GEN_4188 = unuse_way == 2'h2 ? valid_0_0 : _GEN_3480; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4189 = unuse_way == 2'h2 ? valid_0_1 : _GEN_3481; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4190 = unuse_way == 2'h2 ? valid_0_2 : _GEN_3482; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4191 = unuse_way == 2'h2 ? valid_0_3 : _GEN_3483; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4192 = unuse_way == 2'h2 ? valid_0_4 : _GEN_3484; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4193 = unuse_way == 2'h2 ? valid_0_5 : _GEN_3485; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4194 = unuse_way == 2'h2 ? valid_0_6 : _GEN_3486; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4195 = unuse_way == 2'h2 ? valid_0_7 : _GEN_3487; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4196 = unuse_way == 2'h2 ? valid_0_8 : _GEN_3488; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4197 = unuse_way == 2'h2 ? valid_0_9 : _GEN_3489; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4198 = unuse_way == 2'h2 ? valid_0_10 : _GEN_3490; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4199 = unuse_way == 2'h2 ? valid_0_11 : _GEN_3491; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4200 = unuse_way == 2'h2 ? valid_0_12 : _GEN_3492; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4201 = unuse_way == 2'h2 ? valid_0_13 : _GEN_3493; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4202 = unuse_way == 2'h2 ? valid_0_14 : _GEN_3494; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4203 = unuse_way == 2'h2 ? valid_0_15 : _GEN_3495; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4204 = unuse_way == 2'h2 ? valid_0_16 : _GEN_3496; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4205 = unuse_way == 2'h2 ? valid_0_17 : _GEN_3497; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4206 = unuse_way == 2'h2 ? valid_0_18 : _GEN_3498; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4207 = unuse_way == 2'h2 ? valid_0_19 : _GEN_3499; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4208 = unuse_way == 2'h2 ? valid_0_20 : _GEN_3500; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4209 = unuse_way == 2'h2 ? valid_0_21 : _GEN_3501; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4210 = unuse_way == 2'h2 ? valid_0_22 : _GEN_3502; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4211 = unuse_way == 2'h2 ? valid_0_23 : _GEN_3503; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4212 = unuse_way == 2'h2 ? valid_0_24 : _GEN_3504; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4213 = unuse_way == 2'h2 ? valid_0_25 : _GEN_3505; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4214 = unuse_way == 2'h2 ? valid_0_26 : _GEN_3506; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4215 = unuse_way == 2'h2 ? valid_0_27 : _GEN_3507; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4216 = unuse_way == 2'h2 ? valid_0_28 : _GEN_3508; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4217 = unuse_way == 2'h2 ? valid_0_29 : _GEN_3509; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4218 = unuse_way == 2'h2 ? valid_0_30 : _GEN_3510; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4219 = unuse_way == 2'h2 ? valid_0_31 : _GEN_3511; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4220 = unuse_way == 2'h2 ? valid_0_32 : _GEN_3512; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4221 = unuse_way == 2'h2 ? valid_0_33 : _GEN_3513; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4222 = unuse_way == 2'h2 ? valid_0_34 : _GEN_3514; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4223 = unuse_way == 2'h2 ? valid_0_35 : _GEN_3515; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4224 = unuse_way == 2'h2 ? valid_0_36 : _GEN_3516; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4225 = unuse_way == 2'h2 ? valid_0_37 : _GEN_3517; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4226 = unuse_way == 2'h2 ? valid_0_38 : _GEN_3518; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4227 = unuse_way == 2'h2 ? valid_0_39 : _GEN_3519; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4228 = unuse_way == 2'h2 ? valid_0_40 : _GEN_3520; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4229 = unuse_way == 2'h2 ? valid_0_41 : _GEN_3521; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4230 = unuse_way == 2'h2 ? valid_0_42 : _GEN_3522; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4231 = unuse_way == 2'h2 ? valid_0_43 : _GEN_3523; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4232 = unuse_way == 2'h2 ? valid_0_44 : _GEN_3524; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4233 = unuse_way == 2'h2 ? valid_0_45 : _GEN_3525; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4234 = unuse_way == 2'h2 ? valid_0_46 : _GEN_3526; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4235 = unuse_way == 2'h2 ? valid_0_47 : _GEN_3527; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4236 = unuse_way == 2'h2 ? valid_0_48 : _GEN_3528; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4237 = unuse_way == 2'h2 ? valid_0_49 : _GEN_3529; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4238 = unuse_way == 2'h2 ? valid_0_50 : _GEN_3530; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4239 = unuse_way == 2'h2 ? valid_0_51 : _GEN_3531; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4240 = unuse_way == 2'h2 ? valid_0_52 : _GEN_3532; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4241 = unuse_way == 2'h2 ? valid_0_53 : _GEN_3533; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4242 = unuse_way == 2'h2 ? valid_0_54 : _GEN_3534; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4243 = unuse_way == 2'h2 ? valid_0_55 : _GEN_3535; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4244 = unuse_way == 2'h2 ? valid_0_56 : _GEN_3536; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4245 = unuse_way == 2'h2 ? valid_0_57 : _GEN_3537; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4246 = unuse_way == 2'h2 ? valid_0_58 : _GEN_3538; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4247 = unuse_way == 2'h2 ? valid_0_59 : _GEN_3539; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4248 = unuse_way == 2'h2 ? valid_0_60 : _GEN_3540; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4249 = unuse_way == 2'h2 ? valid_0_61 : _GEN_3541; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4250 = unuse_way == 2'h2 ? valid_0_62 : _GEN_3542; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4251 = unuse_way == 2'h2 ? valid_0_63 : _GEN_3543; // @[d_cache.scala 147:40 24:26]
  wire  _GEN_4252 = unuse_way == 2'h2 ? dirty_1_0 : _GEN_3673; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4253 = unuse_way == 2'h2 ? dirty_1_1 : _GEN_3674; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4254 = unuse_way == 2'h2 ? dirty_1_2 : _GEN_3675; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4255 = unuse_way == 2'h2 ? dirty_1_3 : _GEN_3676; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4256 = unuse_way == 2'h2 ? dirty_1_4 : _GEN_3677; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4257 = unuse_way == 2'h2 ? dirty_1_5 : _GEN_3678; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4258 = unuse_way == 2'h2 ? dirty_1_6 : _GEN_3679; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4259 = unuse_way == 2'h2 ? dirty_1_7 : _GEN_3680; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4260 = unuse_way == 2'h2 ? dirty_1_8 : _GEN_3681; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4261 = unuse_way == 2'h2 ? dirty_1_9 : _GEN_3682; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4262 = unuse_way == 2'h2 ? dirty_1_10 : _GEN_3683; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4263 = unuse_way == 2'h2 ? dirty_1_11 : _GEN_3684; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4264 = unuse_way == 2'h2 ? dirty_1_12 : _GEN_3685; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4265 = unuse_way == 2'h2 ? dirty_1_13 : _GEN_3686; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4266 = unuse_way == 2'h2 ? dirty_1_14 : _GEN_3687; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4267 = unuse_way == 2'h2 ? dirty_1_15 : _GEN_3688; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4268 = unuse_way == 2'h2 ? dirty_1_16 : _GEN_3689; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4269 = unuse_way == 2'h2 ? dirty_1_17 : _GEN_3690; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4270 = unuse_way == 2'h2 ? dirty_1_18 : _GEN_3691; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4271 = unuse_way == 2'h2 ? dirty_1_19 : _GEN_3692; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4272 = unuse_way == 2'h2 ? dirty_1_20 : _GEN_3693; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4273 = unuse_way == 2'h2 ? dirty_1_21 : _GEN_3694; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4274 = unuse_way == 2'h2 ? dirty_1_22 : _GEN_3695; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4275 = unuse_way == 2'h2 ? dirty_1_23 : _GEN_3696; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4276 = unuse_way == 2'h2 ? dirty_1_24 : _GEN_3697; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4277 = unuse_way == 2'h2 ? dirty_1_25 : _GEN_3698; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4278 = unuse_way == 2'h2 ? dirty_1_26 : _GEN_3699; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4279 = unuse_way == 2'h2 ? dirty_1_27 : _GEN_3700; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4280 = unuse_way == 2'h2 ? dirty_1_28 : _GEN_3701; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4281 = unuse_way == 2'h2 ? dirty_1_29 : _GEN_3702; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4282 = unuse_way == 2'h2 ? dirty_1_30 : _GEN_3703; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4283 = unuse_way == 2'h2 ? dirty_1_31 : _GEN_3704; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4284 = unuse_way == 2'h2 ? dirty_1_32 : _GEN_3705; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4285 = unuse_way == 2'h2 ? dirty_1_33 : _GEN_3706; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4286 = unuse_way == 2'h2 ? dirty_1_34 : _GEN_3707; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4287 = unuse_way == 2'h2 ? dirty_1_35 : _GEN_3708; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4288 = unuse_way == 2'h2 ? dirty_1_36 : _GEN_3709; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4289 = unuse_way == 2'h2 ? dirty_1_37 : _GEN_3710; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4290 = unuse_way == 2'h2 ? dirty_1_38 : _GEN_3711; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4291 = unuse_way == 2'h2 ? dirty_1_39 : _GEN_3712; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4292 = unuse_way == 2'h2 ? dirty_1_40 : _GEN_3713; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4293 = unuse_way == 2'h2 ? dirty_1_41 : _GEN_3714; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4294 = unuse_way == 2'h2 ? dirty_1_42 : _GEN_3715; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4295 = unuse_way == 2'h2 ? dirty_1_43 : _GEN_3716; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4296 = unuse_way == 2'h2 ? dirty_1_44 : _GEN_3717; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4297 = unuse_way == 2'h2 ? dirty_1_45 : _GEN_3718; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4298 = unuse_way == 2'h2 ? dirty_1_46 : _GEN_3719; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4299 = unuse_way == 2'h2 ? dirty_1_47 : _GEN_3720; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4300 = unuse_way == 2'h2 ? dirty_1_48 : _GEN_3721; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4301 = unuse_way == 2'h2 ? dirty_1_49 : _GEN_3722; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4302 = unuse_way == 2'h2 ? dirty_1_50 : _GEN_3723; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4303 = unuse_way == 2'h2 ? dirty_1_51 : _GEN_3724; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4304 = unuse_way == 2'h2 ? dirty_1_52 : _GEN_3725; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4305 = unuse_way == 2'h2 ? dirty_1_53 : _GEN_3726; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4306 = unuse_way == 2'h2 ? dirty_1_54 : _GEN_3727; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4307 = unuse_way == 2'h2 ? dirty_1_55 : _GEN_3728; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4308 = unuse_way == 2'h2 ? dirty_1_56 : _GEN_3729; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4309 = unuse_way == 2'h2 ? dirty_1_57 : _GEN_3730; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4310 = unuse_way == 2'h2 ? dirty_1_58 : _GEN_3731; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4311 = unuse_way == 2'h2 ? dirty_1_59 : _GEN_3732; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4312 = unuse_way == 2'h2 ? dirty_1_60 : _GEN_3733; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4313 = unuse_way == 2'h2 ? dirty_1_61 : _GEN_3734; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4314 = unuse_way == 2'h2 ? dirty_1_62 : _GEN_3735; // @[d_cache.scala 147:40 27:26]
  wire  _GEN_4315 = unuse_way == 2'h2 ? dirty_1_63 : _GEN_3736; // @[d_cache.scala 147:40 27:26]
  wire [2:0] _GEN_4316 = unuse_way == 2'h1 ? 3'h7 : _GEN_3801; // @[d_cache.scala 141:34 142:23]
  wire [63:0] _GEN_4317 = unuse_way == 2'h1 ? _GEN_1488 : _GEN_3996; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4318 = unuse_way == 2'h1 ? _GEN_1489 : _GEN_3997; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4319 = unuse_way == 2'h1 ? _GEN_1490 : _GEN_3998; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4320 = unuse_way == 2'h1 ? _GEN_1491 : _GEN_3999; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4321 = unuse_way == 2'h1 ? _GEN_1492 : _GEN_4000; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4322 = unuse_way == 2'h1 ? _GEN_1493 : _GEN_4001; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4323 = unuse_way == 2'h1 ? _GEN_1494 : _GEN_4002; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4324 = unuse_way == 2'h1 ? _GEN_1495 : _GEN_4003; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4325 = unuse_way == 2'h1 ? _GEN_1496 : _GEN_4004; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4326 = unuse_way == 2'h1 ? _GEN_1497 : _GEN_4005; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4327 = unuse_way == 2'h1 ? _GEN_1498 : _GEN_4006; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4328 = unuse_way == 2'h1 ? _GEN_1499 : _GEN_4007; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4329 = unuse_way == 2'h1 ? _GEN_1500 : _GEN_4008; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4330 = unuse_way == 2'h1 ? _GEN_1501 : _GEN_4009; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4331 = unuse_way == 2'h1 ? _GEN_1502 : _GEN_4010; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4332 = unuse_way == 2'h1 ? _GEN_1503 : _GEN_4011; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4333 = unuse_way == 2'h1 ? _GEN_1504 : _GEN_4012; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4334 = unuse_way == 2'h1 ? _GEN_1505 : _GEN_4013; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4335 = unuse_way == 2'h1 ? _GEN_1506 : _GEN_4014; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4336 = unuse_way == 2'h1 ? _GEN_1507 : _GEN_4015; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4337 = unuse_way == 2'h1 ? _GEN_1508 : _GEN_4016; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4338 = unuse_way == 2'h1 ? _GEN_1509 : _GEN_4017; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4339 = unuse_way == 2'h1 ? _GEN_1510 : _GEN_4018; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4340 = unuse_way == 2'h1 ? _GEN_1511 : _GEN_4019; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4341 = unuse_way == 2'h1 ? _GEN_1512 : _GEN_4020; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4342 = unuse_way == 2'h1 ? _GEN_1513 : _GEN_4021; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4343 = unuse_way == 2'h1 ? _GEN_1514 : _GEN_4022; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4344 = unuse_way == 2'h1 ? _GEN_1515 : _GEN_4023; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4345 = unuse_way == 2'h1 ? _GEN_1516 : _GEN_4024; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4346 = unuse_way == 2'h1 ? _GEN_1517 : _GEN_4025; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4347 = unuse_way == 2'h1 ? _GEN_1518 : _GEN_4026; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4348 = unuse_way == 2'h1 ? _GEN_1519 : _GEN_4027; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4349 = unuse_way == 2'h1 ? _GEN_1520 : _GEN_4028; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4350 = unuse_way == 2'h1 ? _GEN_1521 : _GEN_4029; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4351 = unuse_way == 2'h1 ? _GEN_1522 : _GEN_4030; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4352 = unuse_way == 2'h1 ? _GEN_1523 : _GEN_4031; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4353 = unuse_way == 2'h1 ? _GEN_1524 : _GEN_4032; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4354 = unuse_way == 2'h1 ? _GEN_1525 : _GEN_4033; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4355 = unuse_way == 2'h1 ? _GEN_1526 : _GEN_4034; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4356 = unuse_way == 2'h1 ? _GEN_1527 : _GEN_4035; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4357 = unuse_way == 2'h1 ? _GEN_1528 : _GEN_4036; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4358 = unuse_way == 2'h1 ? _GEN_1529 : _GEN_4037; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4359 = unuse_way == 2'h1 ? _GEN_1530 : _GEN_4038; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4360 = unuse_way == 2'h1 ? _GEN_1531 : _GEN_4039; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4361 = unuse_way == 2'h1 ? _GEN_1532 : _GEN_4040; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4362 = unuse_way == 2'h1 ? _GEN_1533 : _GEN_4041; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4363 = unuse_way == 2'h1 ? _GEN_1534 : _GEN_4042; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4364 = unuse_way == 2'h1 ? _GEN_1535 : _GEN_4043; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4365 = unuse_way == 2'h1 ? _GEN_1536 : _GEN_4044; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4366 = unuse_way == 2'h1 ? _GEN_1537 : _GEN_4045; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4367 = unuse_way == 2'h1 ? _GEN_1538 : _GEN_4046; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4368 = unuse_way == 2'h1 ? _GEN_1539 : _GEN_4047; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4369 = unuse_way == 2'h1 ? _GEN_1540 : _GEN_4048; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4370 = unuse_way == 2'h1 ? _GEN_1541 : _GEN_4049; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4371 = unuse_way == 2'h1 ? _GEN_1542 : _GEN_4050; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4372 = unuse_way == 2'h1 ? _GEN_1543 : _GEN_4051; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4373 = unuse_way == 2'h1 ? _GEN_1544 : _GEN_4052; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4374 = unuse_way == 2'h1 ? _GEN_1545 : _GEN_4053; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4375 = unuse_way == 2'h1 ? _GEN_1546 : _GEN_4054; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4376 = unuse_way == 2'h1 ? _GEN_1547 : _GEN_4055; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4377 = unuse_way == 2'h1 ? _GEN_1548 : _GEN_4056; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4378 = unuse_way == 2'h1 ? _GEN_1549 : _GEN_4057; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4379 = unuse_way == 2'h1 ? _GEN_1550 : _GEN_4058; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4380 = unuse_way == 2'h1 ? _GEN_1551 : _GEN_4059; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4381 = unuse_way == 2'h1 ? _GEN_1552 : _GEN_4060; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4382 = unuse_way == 2'h1 ? _GEN_1553 : _GEN_4061; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4383 = unuse_way == 2'h1 ? _GEN_1554 : _GEN_4062; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4384 = unuse_way == 2'h1 ? _GEN_1555 : _GEN_4063; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4385 = unuse_way == 2'h1 ? _GEN_1556 : _GEN_4064; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4386 = unuse_way == 2'h1 ? _GEN_1557 : _GEN_4065; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4387 = unuse_way == 2'h1 ? _GEN_1558 : _GEN_4066; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4388 = unuse_way == 2'h1 ? _GEN_1559 : _GEN_4067; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4389 = unuse_way == 2'h1 ? _GEN_1560 : _GEN_4068; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4390 = unuse_way == 2'h1 ? _GEN_1561 : _GEN_4069; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4391 = unuse_way == 2'h1 ? _GEN_1562 : _GEN_4070; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4392 = unuse_way == 2'h1 ? _GEN_1563 : _GEN_4071; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4393 = unuse_way == 2'h1 ? _GEN_1564 : _GEN_4072; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4394 = unuse_way == 2'h1 ? _GEN_1565 : _GEN_4073; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4395 = unuse_way == 2'h1 ? _GEN_1566 : _GEN_4074; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4396 = unuse_way == 2'h1 ? _GEN_1567 : _GEN_4075; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4397 = unuse_way == 2'h1 ? _GEN_1568 : _GEN_4076; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4398 = unuse_way == 2'h1 ? _GEN_1569 : _GEN_4077; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4399 = unuse_way == 2'h1 ? _GEN_1570 : _GEN_4078; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4400 = unuse_way == 2'h1 ? _GEN_1571 : _GEN_4079; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4401 = unuse_way == 2'h1 ? _GEN_1572 : _GEN_4080; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4402 = unuse_way == 2'h1 ? _GEN_1573 : _GEN_4081; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4403 = unuse_way == 2'h1 ? _GEN_1574 : _GEN_4082; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4404 = unuse_way == 2'h1 ? _GEN_1575 : _GEN_4083; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4405 = unuse_way == 2'h1 ? _GEN_1576 : _GEN_4084; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4406 = unuse_way == 2'h1 ? _GEN_1577 : _GEN_4085; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4407 = unuse_way == 2'h1 ? _GEN_1578 : _GEN_4086; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4408 = unuse_way == 2'h1 ? _GEN_1579 : _GEN_4087; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4409 = unuse_way == 2'h1 ? _GEN_1580 : _GEN_4088; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4410 = unuse_way == 2'h1 ? _GEN_1581 : _GEN_4089; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4411 = unuse_way == 2'h1 ? _GEN_1582 : _GEN_4090; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4412 = unuse_way == 2'h1 ? _GEN_1583 : _GEN_4091; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4413 = unuse_way == 2'h1 ? _GEN_1584 : _GEN_4092; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4414 = unuse_way == 2'h1 ? _GEN_1585 : _GEN_4093; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4415 = unuse_way == 2'h1 ? _GEN_1586 : _GEN_4094; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4416 = unuse_way == 2'h1 ? _GEN_1587 : _GEN_4095; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4417 = unuse_way == 2'h1 ? _GEN_1588 : _GEN_4096; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4418 = unuse_way == 2'h1 ? _GEN_1589 : _GEN_4097; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4419 = unuse_way == 2'h1 ? _GEN_1590 : _GEN_4098; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4420 = unuse_way == 2'h1 ? _GEN_1591 : _GEN_4099; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4421 = unuse_way == 2'h1 ? _GEN_1592 : _GEN_4100; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4422 = unuse_way == 2'h1 ? _GEN_1593 : _GEN_4101; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4423 = unuse_way == 2'h1 ? _GEN_1594 : _GEN_4102; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4424 = unuse_way == 2'h1 ? _GEN_1595 : _GEN_4103; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4425 = unuse_way == 2'h1 ? _GEN_1596 : _GEN_4104; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4426 = unuse_way == 2'h1 ? _GEN_1597 : _GEN_4105; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4427 = unuse_way == 2'h1 ? _GEN_1598 : _GEN_4106; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4428 = unuse_way == 2'h1 ? _GEN_1599 : _GEN_4107; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4429 = unuse_way == 2'h1 ? _GEN_1600 : _GEN_4108; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4430 = unuse_way == 2'h1 ? _GEN_1601 : _GEN_4109; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4431 = unuse_way == 2'h1 ? _GEN_1602 : _GEN_4110; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4432 = unuse_way == 2'h1 ? _GEN_1603 : _GEN_4111; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4433 = unuse_way == 2'h1 ? _GEN_1604 : _GEN_4112; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4434 = unuse_way == 2'h1 ? _GEN_1605 : _GEN_4113; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4435 = unuse_way == 2'h1 ? _GEN_1606 : _GEN_4114; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4436 = unuse_way == 2'h1 ? _GEN_1607 : _GEN_4115; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4437 = unuse_way == 2'h1 ? _GEN_1608 : _GEN_4116; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4438 = unuse_way == 2'h1 ? _GEN_1609 : _GEN_4117; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4439 = unuse_way == 2'h1 ? _GEN_1610 : _GEN_4118; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4440 = unuse_way == 2'h1 ? _GEN_1611 : _GEN_4119; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4441 = unuse_way == 2'h1 ? _GEN_1612 : _GEN_4120; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4442 = unuse_way == 2'h1 ? _GEN_1613 : _GEN_4121; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4443 = unuse_way == 2'h1 ? _GEN_1614 : _GEN_4122; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_4444 = unuse_way == 2'h1 ? _GEN_1615 : _GEN_4123; // @[d_cache.scala 141:34]
  wire  _GEN_4445 = unuse_way == 2'h1 ? _GEN_521 : _GEN_4188; // @[d_cache.scala 141:34]
  wire  _GEN_4446 = unuse_way == 2'h1 ? _GEN_522 : _GEN_4189; // @[d_cache.scala 141:34]
  wire  _GEN_4447 = unuse_way == 2'h1 ? _GEN_523 : _GEN_4190; // @[d_cache.scala 141:34]
  wire  _GEN_4448 = unuse_way == 2'h1 ? _GEN_524 : _GEN_4191; // @[d_cache.scala 141:34]
  wire  _GEN_4449 = unuse_way == 2'h1 ? _GEN_525 : _GEN_4192; // @[d_cache.scala 141:34]
  wire  _GEN_4450 = unuse_way == 2'h1 ? _GEN_526 : _GEN_4193; // @[d_cache.scala 141:34]
  wire  _GEN_4451 = unuse_way == 2'h1 ? _GEN_527 : _GEN_4194; // @[d_cache.scala 141:34]
  wire  _GEN_4452 = unuse_way == 2'h1 ? _GEN_528 : _GEN_4195; // @[d_cache.scala 141:34]
  wire  _GEN_4453 = unuse_way == 2'h1 ? _GEN_529 : _GEN_4196; // @[d_cache.scala 141:34]
  wire  _GEN_4454 = unuse_way == 2'h1 ? _GEN_530 : _GEN_4197; // @[d_cache.scala 141:34]
  wire  _GEN_4455 = unuse_way == 2'h1 ? _GEN_531 : _GEN_4198; // @[d_cache.scala 141:34]
  wire  _GEN_4456 = unuse_way == 2'h1 ? _GEN_532 : _GEN_4199; // @[d_cache.scala 141:34]
  wire  _GEN_4457 = unuse_way == 2'h1 ? _GEN_533 : _GEN_4200; // @[d_cache.scala 141:34]
  wire  _GEN_4458 = unuse_way == 2'h1 ? _GEN_534 : _GEN_4201; // @[d_cache.scala 141:34]
  wire  _GEN_4459 = unuse_way == 2'h1 ? _GEN_535 : _GEN_4202; // @[d_cache.scala 141:34]
  wire  _GEN_4460 = unuse_way == 2'h1 ? _GEN_536 : _GEN_4203; // @[d_cache.scala 141:34]
  wire  _GEN_4461 = unuse_way == 2'h1 ? _GEN_537 : _GEN_4204; // @[d_cache.scala 141:34]
  wire  _GEN_4462 = unuse_way == 2'h1 ? _GEN_538 : _GEN_4205; // @[d_cache.scala 141:34]
  wire  _GEN_4463 = unuse_way == 2'h1 ? _GEN_539 : _GEN_4206; // @[d_cache.scala 141:34]
  wire  _GEN_4464 = unuse_way == 2'h1 ? _GEN_540 : _GEN_4207; // @[d_cache.scala 141:34]
  wire  _GEN_4465 = unuse_way == 2'h1 ? _GEN_541 : _GEN_4208; // @[d_cache.scala 141:34]
  wire  _GEN_4466 = unuse_way == 2'h1 ? _GEN_542 : _GEN_4209; // @[d_cache.scala 141:34]
  wire  _GEN_4467 = unuse_way == 2'h1 ? _GEN_543 : _GEN_4210; // @[d_cache.scala 141:34]
  wire  _GEN_4468 = unuse_way == 2'h1 ? _GEN_544 : _GEN_4211; // @[d_cache.scala 141:34]
  wire  _GEN_4469 = unuse_way == 2'h1 ? _GEN_545 : _GEN_4212; // @[d_cache.scala 141:34]
  wire  _GEN_4470 = unuse_way == 2'h1 ? _GEN_546 : _GEN_4213; // @[d_cache.scala 141:34]
  wire  _GEN_4471 = unuse_way == 2'h1 ? _GEN_547 : _GEN_4214; // @[d_cache.scala 141:34]
  wire  _GEN_4472 = unuse_way == 2'h1 ? _GEN_548 : _GEN_4215; // @[d_cache.scala 141:34]
  wire  _GEN_4473 = unuse_way == 2'h1 ? _GEN_549 : _GEN_4216; // @[d_cache.scala 141:34]
  wire  _GEN_4474 = unuse_way == 2'h1 ? _GEN_550 : _GEN_4217; // @[d_cache.scala 141:34]
  wire  _GEN_4475 = unuse_way == 2'h1 ? _GEN_551 : _GEN_4218; // @[d_cache.scala 141:34]
  wire  _GEN_4476 = unuse_way == 2'h1 ? _GEN_552 : _GEN_4219; // @[d_cache.scala 141:34]
  wire  _GEN_4477 = unuse_way == 2'h1 ? _GEN_553 : _GEN_4220; // @[d_cache.scala 141:34]
  wire  _GEN_4478 = unuse_way == 2'h1 ? _GEN_554 : _GEN_4221; // @[d_cache.scala 141:34]
  wire  _GEN_4479 = unuse_way == 2'h1 ? _GEN_555 : _GEN_4222; // @[d_cache.scala 141:34]
  wire  _GEN_4480 = unuse_way == 2'h1 ? _GEN_556 : _GEN_4223; // @[d_cache.scala 141:34]
  wire  _GEN_4481 = unuse_way == 2'h1 ? _GEN_557 : _GEN_4224; // @[d_cache.scala 141:34]
  wire  _GEN_4482 = unuse_way == 2'h1 ? _GEN_558 : _GEN_4225; // @[d_cache.scala 141:34]
  wire  _GEN_4483 = unuse_way == 2'h1 ? _GEN_559 : _GEN_4226; // @[d_cache.scala 141:34]
  wire  _GEN_4484 = unuse_way == 2'h1 ? _GEN_560 : _GEN_4227; // @[d_cache.scala 141:34]
  wire  _GEN_4485 = unuse_way == 2'h1 ? _GEN_561 : _GEN_4228; // @[d_cache.scala 141:34]
  wire  _GEN_4486 = unuse_way == 2'h1 ? _GEN_562 : _GEN_4229; // @[d_cache.scala 141:34]
  wire  _GEN_4487 = unuse_way == 2'h1 ? _GEN_563 : _GEN_4230; // @[d_cache.scala 141:34]
  wire  _GEN_4488 = unuse_way == 2'h1 ? _GEN_564 : _GEN_4231; // @[d_cache.scala 141:34]
  wire  _GEN_4489 = unuse_way == 2'h1 ? _GEN_565 : _GEN_4232; // @[d_cache.scala 141:34]
  wire  _GEN_4490 = unuse_way == 2'h1 ? _GEN_566 : _GEN_4233; // @[d_cache.scala 141:34]
  wire  _GEN_4491 = unuse_way == 2'h1 ? _GEN_567 : _GEN_4234; // @[d_cache.scala 141:34]
  wire  _GEN_4492 = unuse_way == 2'h1 ? _GEN_568 : _GEN_4235; // @[d_cache.scala 141:34]
  wire  _GEN_4493 = unuse_way == 2'h1 ? _GEN_569 : _GEN_4236; // @[d_cache.scala 141:34]
  wire  _GEN_4494 = unuse_way == 2'h1 ? _GEN_570 : _GEN_4237; // @[d_cache.scala 141:34]
  wire  _GEN_4495 = unuse_way == 2'h1 ? _GEN_571 : _GEN_4238; // @[d_cache.scala 141:34]
  wire  _GEN_4496 = unuse_way == 2'h1 ? _GEN_572 : _GEN_4239; // @[d_cache.scala 141:34]
  wire  _GEN_4497 = unuse_way == 2'h1 ? _GEN_573 : _GEN_4240; // @[d_cache.scala 141:34]
  wire  _GEN_4498 = unuse_way == 2'h1 ? _GEN_574 : _GEN_4241; // @[d_cache.scala 141:34]
  wire  _GEN_4499 = unuse_way == 2'h1 ? _GEN_575 : _GEN_4242; // @[d_cache.scala 141:34]
  wire  _GEN_4500 = unuse_way == 2'h1 ? _GEN_576 : _GEN_4243; // @[d_cache.scala 141:34]
  wire  _GEN_4501 = unuse_way == 2'h1 ? _GEN_577 : _GEN_4244; // @[d_cache.scala 141:34]
  wire  _GEN_4502 = unuse_way == 2'h1 ? _GEN_578 : _GEN_4245; // @[d_cache.scala 141:34]
  wire  _GEN_4503 = unuse_way == 2'h1 ? _GEN_579 : _GEN_4246; // @[d_cache.scala 141:34]
  wire  _GEN_4504 = unuse_way == 2'h1 ? _GEN_580 : _GEN_4247; // @[d_cache.scala 141:34]
  wire  _GEN_4505 = unuse_way == 2'h1 ? _GEN_581 : _GEN_4248; // @[d_cache.scala 141:34]
  wire  _GEN_4506 = unuse_way == 2'h1 ? _GEN_582 : _GEN_4249; // @[d_cache.scala 141:34]
  wire  _GEN_4507 = unuse_way == 2'h1 ? _GEN_583 : _GEN_4250; // @[d_cache.scala 141:34]
  wire  _GEN_4508 = unuse_way == 2'h1 ? _GEN_584 : _GEN_4251; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_4509 = unuse_way == 2'h1 ? ram_1_0 : _GEN_3802; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4510 = unuse_way == 2'h1 ? ram_1_1 : _GEN_3803; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4511 = unuse_way == 2'h1 ? ram_1_2 : _GEN_3804; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4512 = unuse_way == 2'h1 ? ram_1_3 : _GEN_3805; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4513 = unuse_way == 2'h1 ? ram_1_4 : _GEN_3806; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4514 = unuse_way == 2'h1 ? ram_1_5 : _GEN_3807; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4515 = unuse_way == 2'h1 ? ram_1_6 : _GEN_3808; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4516 = unuse_way == 2'h1 ? ram_1_7 : _GEN_3809; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4517 = unuse_way == 2'h1 ? ram_1_8 : _GEN_3810; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4518 = unuse_way == 2'h1 ? ram_1_9 : _GEN_3811; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4519 = unuse_way == 2'h1 ? ram_1_10 : _GEN_3812; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4520 = unuse_way == 2'h1 ? ram_1_11 : _GEN_3813; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4521 = unuse_way == 2'h1 ? ram_1_12 : _GEN_3814; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4522 = unuse_way == 2'h1 ? ram_1_13 : _GEN_3815; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4523 = unuse_way == 2'h1 ? ram_1_14 : _GEN_3816; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4524 = unuse_way == 2'h1 ? ram_1_15 : _GEN_3817; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4525 = unuse_way == 2'h1 ? ram_1_16 : _GEN_3818; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4526 = unuse_way == 2'h1 ? ram_1_17 : _GEN_3819; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4527 = unuse_way == 2'h1 ? ram_1_18 : _GEN_3820; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4528 = unuse_way == 2'h1 ? ram_1_19 : _GEN_3821; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4529 = unuse_way == 2'h1 ? ram_1_20 : _GEN_3822; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4530 = unuse_way == 2'h1 ? ram_1_21 : _GEN_3823; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4531 = unuse_way == 2'h1 ? ram_1_22 : _GEN_3824; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4532 = unuse_way == 2'h1 ? ram_1_23 : _GEN_3825; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4533 = unuse_way == 2'h1 ? ram_1_24 : _GEN_3826; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4534 = unuse_way == 2'h1 ? ram_1_25 : _GEN_3827; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4535 = unuse_way == 2'h1 ? ram_1_26 : _GEN_3828; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4536 = unuse_way == 2'h1 ? ram_1_27 : _GEN_3829; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4537 = unuse_way == 2'h1 ? ram_1_28 : _GEN_3830; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4538 = unuse_way == 2'h1 ? ram_1_29 : _GEN_3831; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4539 = unuse_way == 2'h1 ? ram_1_30 : _GEN_3832; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4540 = unuse_way == 2'h1 ? ram_1_31 : _GEN_3833; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4541 = unuse_way == 2'h1 ? ram_1_32 : _GEN_3834; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4542 = unuse_way == 2'h1 ? ram_1_33 : _GEN_3835; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4543 = unuse_way == 2'h1 ? ram_1_34 : _GEN_3836; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4544 = unuse_way == 2'h1 ? ram_1_35 : _GEN_3837; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4545 = unuse_way == 2'h1 ? ram_1_36 : _GEN_3838; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4546 = unuse_way == 2'h1 ? ram_1_37 : _GEN_3839; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4547 = unuse_way == 2'h1 ? ram_1_38 : _GEN_3840; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4548 = unuse_way == 2'h1 ? ram_1_39 : _GEN_3841; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4549 = unuse_way == 2'h1 ? ram_1_40 : _GEN_3842; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4550 = unuse_way == 2'h1 ? ram_1_41 : _GEN_3843; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4551 = unuse_way == 2'h1 ? ram_1_42 : _GEN_3844; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4552 = unuse_way == 2'h1 ? ram_1_43 : _GEN_3845; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4553 = unuse_way == 2'h1 ? ram_1_44 : _GEN_3846; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4554 = unuse_way == 2'h1 ? ram_1_45 : _GEN_3847; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4555 = unuse_way == 2'h1 ? ram_1_46 : _GEN_3848; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4556 = unuse_way == 2'h1 ? ram_1_47 : _GEN_3849; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4557 = unuse_way == 2'h1 ? ram_1_48 : _GEN_3850; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4558 = unuse_way == 2'h1 ? ram_1_49 : _GEN_3851; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4559 = unuse_way == 2'h1 ? ram_1_50 : _GEN_3852; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4560 = unuse_way == 2'h1 ? ram_1_51 : _GEN_3853; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4561 = unuse_way == 2'h1 ? ram_1_52 : _GEN_3854; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4562 = unuse_way == 2'h1 ? ram_1_53 : _GEN_3855; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4563 = unuse_way == 2'h1 ? ram_1_54 : _GEN_3856; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4564 = unuse_way == 2'h1 ? ram_1_55 : _GEN_3857; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4565 = unuse_way == 2'h1 ? ram_1_56 : _GEN_3858; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4566 = unuse_way == 2'h1 ? ram_1_57 : _GEN_3859; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4567 = unuse_way == 2'h1 ? ram_1_58 : _GEN_3860; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4568 = unuse_way == 2'h1 ? ram_1_59 : _GEN_3861; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4569 = unuse_way == 2'h1 ? ram_1_60 : _GEN_3862; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4570 = unuse_way == 2'h1 ? ram_1_61 : _GEN_3863; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4571 = unuse_way == 2'h1 ? ram_1_62 : _GEN_3864; // @[d_cache.scala 141:34 19:24]
  wire [63:0] _GEN_4572 = unuse_way == 2'h1 ? ram_1_63 : _GEN_3865; // @[d_cache.scala 141:34 19:24]
  wire [31:0] _GEN_4573 = unuse_way == 2'h1 ? tag_1_0 : _GEN_3866; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4574 = unuse_way == 2'h1 ? tag_1_1 : _GEN_3867; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4575 = unuse_way == 2'h1 ? tag_1_2 : _GEN_3868; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4576 = unuse_way == 2'h1 ? tag_1_3 : _GEN_3869; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4577 = unuse_way == 2'h1 ? tag_1_4 : _GEN_3870; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4578 = unuse_way == 2'h1 ? tag_1_5 : _GEN_3871; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4579 = unuse_way == 2'h1 ? tag_1_6 : _GEN_3872; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4580 = unuse_way == 2'h1 ? tag_1_7 : _GEN_3873; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4581 = unuse_way == 2'h1 ? tag_1_8 : _GEN_3874; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4582 = unuse_way == 2'h1 ? tag_1_9 : _GEN_3875; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4583 = unuse_way == 2'h1 ? tag_1_10 : _GEN_3876; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4584 = unuse_way == 2'h1 ? tag_1_11 : _GEN_3877; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4585 = unuse_way == 2'h1 ? tag_1_12 : _GEN_3878; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4586 = unuse_way == 2'h1 ? tag_1_13 : _GEN_3879; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4587 = unuse_way == 2'h1 ? tag_1_14 : _GEN_3880; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4588 = unuse_way == 2'h1 ? tag_1_15 : _GEN_3881; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4589 = unuse_way == 2'h1 ? tag_1_16 : _GEN_3882; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4590 = unuse_way == 2'h1 ? tag_1_17 : _GEN_3883; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4591 = unuse_way == 2'h1 ? tag_1_18 : _GEN_3884; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4592 = unuse_way == 2'h1 ? tag_1_19 : _GEN_3885; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4593 = unuse_way == 2'h1 ? tag_1_20 : _GEN_3886; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4594 = unuse_way == 2'h1 ? tag_1_21 : _GEN_3887; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4595 = unuse_way == 2'h1 ? tag_1_22 : _GEN_3888; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4596 = unuse_way == 2'h1 ? tag_1_23 : _GEN_3889; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4597 = unuse_way == 2'h1 ? tag_1_24 : _GEN_3890; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4598 = unuse_way == 2'h1 ? tag_1_25 : _GEN_3891; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4599 = unuse_way == 2'h1 ? tag_1_26 : _GEN_3892; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4600 = unuse_way == 2'h1 ? tag_1_27 : _GEN_3893; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4601 = unuse_way == 2'h1 ? tag_1_28 : _GEN_3894; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4602 = unuse_way == 2'h1 ? tag_1_29 : _GEN_3895; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4603 = unuse_way == 2'h1 ? tag_1_30 : _GEN_3896; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4604 = unuse_way == 2'h1 ? tag_1_31 : _GEN_3897; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4605 = unuse_way == 2'h1 ? tag_1_32 : _GEN_3898; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4606 = unuse_way == 2'h1 ? tag_1_33 : _GEN_3899; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4607 = unuse_way == 2'h1 ? tag_1_34 : _GEN_3900; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4608 = unuse_way == 2'h1 ? tag_1_35 : _GEN_3901; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4609 = unuse_way == 2'h1 ? tag_1_36 : _GEN_3902; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4610 = unuse_way == 2'h1 ? tag_1_37 : _GEN_3903; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4611 = unuse_way == 2'h1 ? tag_1_38 : _GEN_3904; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4612 = unuse_way == 2'h1 ? tag_1_39 : _GEN_3905; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4613 = unuse_way == 2'h1 ? tag_1_40 : _GEN_3906; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4614 = unuse_way == 2'h1 ? tag_1_41 : _GEN_3907; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4615 = unuse_way == 2'h1 ? tag_1_42 : _GEN_3908; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4616 = unuse_way == 2'h1 ? tag_1_43 : _GEN_3909; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4617 = unuse_way == 2'h1 ? tag_1_44 : _GEN_3910; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4618 = unuse_way == 2'h1 ? tag_1_45 : _GEN_3911; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4619 = unuse_way == 2'h1 ? tag_1_46 : _GEN_3912; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4620 = unuse_way == 2'h1 ? tag_1_47 : _GEN_3913; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4621 = unuse_way == 2'h1 ? tag_1_48 : _GEN_3914; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4622 = unuse_way == 2'h1 ? tag_1_49 : _GEN_3915; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4623 = unuse_way == 2'h1 ? tag_1_50 : _GEN_3916; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4624 = unuse_way == 2'h1 ? tag_1_51 : _GEN_3917; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4625 = unuse_way == 2'h1 ? tag_1_52 : _GEN_3918; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4626 = unuse_way == 2'h1 ? tag_1_53 : _GEN_3919; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4627 = unuse_way == 2'h1 ? tag_1_54 : _GEN_3920; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4628 = unuse_way == 2'h1 ? tag_1_55 : _GEN_3921; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4629 = unuse_way == 2'h1 ? tag_1_56 : _GEN_3922; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4630 = unuse_way == 2'h1 ? tag_1_57 : _GEN_3923; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4631 = unuse_way == 2'h1 ? tag_1_58 : _GEN_3924; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4632 = unuse_way == 2'h1 ? tag_1_59 : _GEN_3925; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4633 = unuse_way == 2'h1 ? tag_1_60 : _GEN_3926; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4634 = unuse_way == 2'h1 ? tag_1_61 : _GEN_3927; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4635 = unuse_way == 2'h1 ? tag_1_62 : _GEN_3928; // @[d_cache.scala 141:34 23:24]
  wire [31:0] _GEN_4636 = unuse_way == 2'h1 ? tag_1_63 : _GEN_3929; // @[d_cache.scala 141:34 23:24]
  wire  _GEN_4637 = unuse_way == 2'h1 ? valid_1_0 : _GEN_3930; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4638 = unuse_way == 2'h1 ? valid_1_1 : _GEN_3931; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4639 = unuse_way == 2'h1 ? valid_1_2 : _GEN_3932; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4640 = unuse_way == 2'h1 ? valid_1_3 : _GEN_3933; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4641 = unuse_way == 2'h1 ? valid_1_4 : _GEN_3934; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4642 = unuse_way == 2'h1 ? valid_1_5 : _GEN_3935; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4643 = unuse_way == 2'h1 ? valid_1_6 : _GEN_3936; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4644 = unuse_way == 2'h1 ? valid_1_7 : _GEN_3937; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4645 = unuse_way == 2'h1 ? valid_1_8 : _GEN_3938; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4646 = unuse_way == 2'h1 ? valid_1_9 : _GEN_3939; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4647 = unuse_way == 2'h1 ? valid_1_10 : _GEN_3940; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4648 = unuse_way == 2'h1 ? valid_1_11 : _GEN_3941; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4649 = unuse_way == 2'h1 ? valid_1_12 : _GEN_3942; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4650 = unuse_way == 2'h1 ? valid_1_13 : _GEN_3943; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4651 = unuse_way == 2'h1 ? valid_1_14 : _GEN_3944; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4652 = unuse_way == 2'h1 ? valid_1_15 : _GEN_3945; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4653 = unuse_way == 2'h1 ? valid_1_16 : _GEN_3946; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4654 = unuse_way == 2'h1 ? valid_1_17 : _GEN_3947; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4655 = unuse_way == 2'h1 ? valid_1_18 : _GEN_3948; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4656 = unuse_way == 2'h1 ? valid_1_19 : _GEN_3949; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4657 = unuse_way == 2'h1 ? valid_1_20 : _GEN_3950; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4658 = unuse_way == 2'h1 ? valid_1_21 : _GEN_3951; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4659 = unuse_way == 2'h1 ? valid_1_22 : _GEN_3952; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4660 = unuse_way == 2'h1 ? valid_1_23 : _GEN_3953; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4661 = unuse_way == 2'h1 ? valid_1_24 : _GEN_3954; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4662 = unuse_way == 2'h1 ? valid_1_25 : _GEN_3955; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4663 = unuse_way == 2'h1 ? valid_1_26 : _GEN_3956; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4664 = unuse_way == 2'h1 ? valid_1_27 : _GEN_3957; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4665 = unuse_way == 2'h1 ? valid_1_28 : _GEN_3958; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4666 = unuse_way == 2'h1 ? valid_1_29 : _GEN_3959; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4667 = unuse_way == 2'h1 ? valid_1_30 : _GEN_3960; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4668 = unuse_way == 2'h1 ? valid_1_31 : _GEN_3961; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4669 = unuse_way == 2'h1 ? valid_1_32 : _GEN_3962; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4670 = unuse_way == 2'h1 ? valid_1_33 : _GEN_3963; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4671 = unuse_way == 2'h1 ? valid_1_34 : _GEN_3964; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4672 = unuse_way == 2'h1 ? valid_1_35 : _GEN_3965; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4673 = unuse_way == 2'h1 ? valid_1_36 : _GEN_3966; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4674 = unuse_way == 2'h1 ? valid_1_37 : _GEN_3967; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4675 = unuse_way == 2'h1 ? valid_1_38 : _GEN_3968; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4676 = unuse_way == 2'h1 ? valid_1_39 : _GEN_3969; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4677 = unuse_way == 2'h1 ? valid_1_40 : _GEN_3970; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4678 = unuse_way == 2'h1 ? valid_1_41 : _GEN_3971; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4679 = unuse_way == 2'h1 ? valid_1_42 : _GEN_3972; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4680 = unuse_way == 2'h1 ? valid_1_43 : _GEN_3973; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4681 = unuse_way == 2'h1 ? valid_1_44 : _GEN_3974; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4682 = unuse_way == 2'h1 ? valid_1_45 : _GEN_3975; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4683 = unuse_way == 2'h1 ? valid_1_46 : _GEN_3976; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4684 = unuse_way == 2'h1 ? valid_1_47 : _GEN_3977; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4685 = unuse_way == 2'h1 ? valid_1_48 : _GEN_3978; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4686 = unuse_way == 2'h1 ? valid_1_49 : _GEN_3979; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4687 = unuse_way == 2'h1 ? valid_1_50 : _GEN_3980; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4688 = unuse_way == 2'h1 ? valid_1_51 : _GEN_3981; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4689 = unuse_way == 2'h1 ? valid_1_52 : _GEN_3982; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4690 = unuse_way == 2'h1 ? valid_1_53 : _GEN_3983; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4691 = unuse_way == 2'h1 ? valid_1_54 : _GEN_3984; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4692 = unuse_way == 2'h1 ? valid_1_55 : _GEN_3985; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4693 = unuse_way == 2'h1 ? valid_1_56 : _GEN_3986; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4694 = unuse_way == 2'h1 ? valid_1_57 : _GEN_3987; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4695 = unuse_way == 2'h1 ? valid_1_58 : _GEN_3988; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4696 = unuse_way == 2'h1 ? valid_1_59 : _GEN_3989; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4697 = unuse_way == 2'h1 ? valid_1_60 : _GEN_3990; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4698 = unuse_way == 2'h1 ? valid_1_61 : _GEN_3991; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4699 = unuse_way == 2'h1 ? valid_1_62 : _GEN_3992; // @[d_cache.scala 141:34 25:26]
  wire  _GEN_4700 = unuse_way == 2'h1 ? valid_1_63 : _GEN_3993; // @[d_cache.scala 141:34 25:26]
  wire [63:0] _GEN_4701 = unuse_way == 2'h1 ? write_back_data : _GEN_3994; // @[d_cache.scala 141:34 31:34]
  wire [40:0] _GEN_4702 = unuse_way == 2'h1 ? {{9'd0}, write_back_addr} : _GEN_3995; // @[d_cache.scala 141:34 32:34]
  wire  _GEN_4703 = unuse_way == 2'h1 ? dirty_0_0 : _GEN_4124; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4704 = unuse_way == 2'h1 ? dirty_0_1 : _GEN_4125; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4705 = unuse_way == 2'h1 ? dirty_0_2 : _GEN_4126; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4706 = unuse_way == 2'h1 ? dirty_0_3 : _GEN_4127; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4707 = unuse_way == 2'h1 ? dirty_0_4 : _GEN_4128; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4708 = unuse_way == 2'h1 ? dirty_0_5 : _GEN_4129; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4709 = unuse_way == 2'h1 ? dirty_0_6 : _GEN_4130; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4710 = unuse_way == 2'h1 ? dirty_0_7 : _GEN_4131; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4711 = unuse_way == 2'h1 ? dirty_0_8 : _GEN_4132; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4712 = unuse_way == 2'h1 ? dirty_0_9 : _GEN_4133; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4713 = unuse_way == 2'h1 ? dirty_0_10 : _GEN_4134; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4714 = unuse_way == 2'h1 ? dirty_0_11 : _GEN_4135; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4715 = unuse_way == 2'h1 ? dirty_0_12 : _GEN_4136; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4716 = unuse_way == 2'h1 ? dirty_0_13 : _GEN_4137; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4717 = unuse_way == 2'h1 ? dirty_0_14 : _GEN_4138; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4718 = unuse_way == 2'h1 ? dirty_0_15 : _GEN_4139; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4719 = unuse_way == 2'h1 ? dirty_0_16 : _GEN_4140; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4720 = unuse_way == 2'h1 ? dirty_0_17 : _GEN_4141; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4721 = unuse_way == 2'h1 ? dirty_0_18 : _GEN_4142; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4722 = unuse_way == 2'h1 ? dirty_0_19 : _GEN_4143; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4723 = unuse_way == 2'h1 ? dirty_0_20 : _GEN_4144; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4724 = unuse_way == 2'h1 ? dirty_0_21 : _GEN_4145; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4725 = unuse_way == 2'h1 ? dirty_0_22 : _GEN_4146; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4726 = unuse_way == 2'h1 ? dirty_0_23 : _GEN_4147; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4727 = unuse_way == 2'h1 ? dirty_0_24 : _GEN_4148; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4728 = unuse_way == 2'h1 ? dirty_0_25 : _GEN_4149; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4729 = unuse_way == 2'h1 ? dirty_0_26 : _GEN_4150; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4730 = unuse_way == 2'h1 ? dirty_0_27 : _GEN_4151; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4731 = unuse_way == 2'h1 ? dirty_0_28 : _GEN_4152; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4732 = unuse_way == 2'h1 ? dirty_0_29 : _GEN_4153; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4733 = unuse_way == 2'h1 ? dirty_0_30 : _GEN_4154; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4734 = unuse_way == 2'h1 ? dirty_0_31 : _GEN_4155; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4735 = unuse_way == 2'h1 ? dirty_0_32 : _GEN_4156; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4736 = unuse_way == 2'h1 ? dirty_0_33 : _GEN_4157; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4737 = unuse_way == 2'h1 ? dirty_0_34 : _GEN_4158; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4738 = unuse_way == 2'h1 ? dirty_0_35 : _GEN_4159; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4739 = unuse_way == 2'h1 ? dirty_0_36 : _GEN_4160; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4740 = unuse_way == 2'h1 ? dirty_0_37 : _GEN_4161; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4741 = unuse_way == 2'h1 ? dirty_0_38 : _GEN_4162; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4742 = unuse_way == 2'h1 ? dirty_0_39 : _GEN_4163; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4743 = unuse_way == 2'h1 ? dirty_0_40 : _GEN_4164; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4744 = unuse_way == 2'h1 ? dirty_0_41 : _GEN_4165; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4745 = unuse_way == 2'h1 ? dirty_0_42 : _GEN_4166; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4746 = unuse_way == 2'h1 ? dirty_0_43 : _GEN_4167; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4747 = unuse_way == 2'h1 ? dirty_0_44 : _GEN_4168; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4748 = unuse_way == 2'h1 ? dirty_0_45 : _GEN_4169; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4749 = unuse_way == 2'h1 ? dirty_0_46 : _GEN_4170; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4750 = unuse_way == 2'h1 ? dirty_0_47 : _GEN_4171; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4751 = unuse_way == 2'h1 ? dirty_0_48 : _GEN_4172; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4752 = unuse_way == 2'h1 ? dirty_0_49 : _GEN_4173; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4753 = unuse_way == 2'h1 ? dirty_0_50 : _GEN_4174; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4754 = unuse_way == 2'h1 ? dirty_0_51 : _GEN_4175; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4755 = unuse_way == 2'h1 ? dirty_0_52 : _GEN_4176; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4756 = unuse_way == 2'h1 ? dirty_0_53 : _GEN_4177; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4757 = unuse_way == 2'h1 ? dirty_0_54 : _GEN_4178; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4758 = unuse_way == 2'h1 ? dirty_0_55 : _GEN_4179; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4759 = unuse_way == 2'h1 ? dirty_0_56 : _GEN_4180; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4760 = unuse_way == 2'h1 ? dirty_0_57 : _GEN_4181; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4761 = unuse_way == 2'h1 ? dirty_0_58 : _GEN_4182; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4762 = unuse_way == 2'h1 ? dirty_0_59 : _GEN_4183; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4763 = unuse_way == 2'h1 ? dirty_0_60 : _GEN_4184; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4764 = unuse_way == 2'h1 ? dirty_0_61 : _GEN_4185; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4765 = unuse_way == 2'h1 ? dirty_0_62 : _GEN_4186; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4766 = unuse_way == 2'h1 ? dirty_0_63 : _GEN_4187; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_4767 = unuse_way == 2'h1 ? dirty_1_0 : _GEN_4252; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4768 = unuse_way == 2'h1 ? dirty_1_1 : _GEN_4253; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4769 = unuse_way == 2'h1 ? dirty_1_2 : _GEN_4254; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4770 = unuse_way == 2'h1 ? dirty_1_3 : _GEN_4255; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4771 = unuse_way == 2'h1 ? dirty_1_4 : _GEN_4256; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4772 = unuse_way == 2'h1 ? dirty_1_5 : _GEN_4257; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4773 = unuse_way == 2'h1 ? dirty_1_6 : _GEN_4258; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4774 = unuse_way == 2'h1 ? dirty_1_7 : _GEN_4259; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4775 = unuse_way == 2'h1 ? dirty_1_8 : _GEN_4260; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4776 = unuse_way == 2'h1 ? dirty_1_9 : _GEN_4261; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4777 = unuse_way == 2'h1 ? dirty_1_10 : _GEN_4262; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4778 = unuse_way == 2'h1 ? dirty_1_11 : _GEN_4263; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4779 = unuse_way == 2'h1 ? dirty_1_12 : _GEN_4264; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4780 = unuse_way == 2'h1 ? dirty_1_13 : _GEN_4265; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4781 = unuse_way == 2'h1 ? dirty_1_14 : _GEN_4266; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4782 = unuse_way == 2'h1 ? dirty_1_15 : _GEN_4267; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4783 = unuse_way == 2'h1 ? dirty_1_16 : _GEN_4268; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4784 = unuse_way == 2'h1 ? dirty_1_17 : _GEN_4269; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4785 = unuse_way == 2'h1 ? dirty_1_18 : _GEN_4270; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4786 = unuse_way == 2'h1 ? dirty_1_19 : _GEN_4271; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4787 = unuse_way == 2'h1 ? dirty_1_20 : _GEN_4272; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4788 = unuse_way == 2'h1 ? dirty_1_21 : _GEN_4273; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4789 = unuse_way == 2'h1 ? dirty_1_22 : _GEN_4274; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4790 = unuse_way == 2'h1 ? dirty_1_23 : _GEN_4275; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4791 = unuse_way == 2'h1 ? dirty_1_24 : _GEN_4276; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4792 = unuse_way == 2'h1 ? dirty_1_25 : _GEN_4277; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4793 = unuse_way == 2'h1 ? dirty_1_26 : _GEN_4278; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4794 = unuse_way == 2'h1 ? dirty_1_27 : _GEN_4279; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4795 = unuse_way == 2'h1 ? dirty_1_28 : _GEN_4280; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4796 = unuse_way == 2'h1 ? dirty_1_29 : _GEN_4281; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4797 = unuse_way == 2'h1 ? dirty_1_30 : _GEN_4282; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4798 = unuse_way == 2'h1 ? dirty_1_31 : _GEN_4283; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4799 = unuse_way == 2'h1 ? dirty_1_32 : _GEN_4284; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4800 = unuse_way == 2'h1 ? dirty_1_33 : _GEN_4285; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4801 = unuse_way == 2'h1 ? dirty_1_34 : _GEN_4286; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4802 = unuse_way == 2'h1 ? dirty_1_35 : _GEN_4287; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4803 = unuse_way == 2'h1 ? dirty_1_36 : _GEN_4288; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4804 = unuse_way == 2'h1 ? dirty_1_37 : _GEN_4289; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4805 = unuse_way == 2'h1 ? dirty_1_38 : _GEN_4290; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4806 = unuse_way == 2'h1 ? dirty_1_39 : _GEN_4291; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4807 = unuse_way == 2'h1 ? dirty_1_40 : _GEN_4292; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4808 = unuse_way == 2'h1 ? dirty_1_41 : _GEN_4293; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4809 = unuse_way == 2'h1 ? dirty_1_42 : _GEN_4294; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4810 = unuse_way == 2'h1 ? dirty_1_43 : _GEN_4295; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4811 = unuse_way == 2'h1 ? dirty_1_44 : _GEN_4296; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4812 = unuse_way == 2'h1 ? dirty_1_45 : _GEN_4297; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4813 = unuse_way == 2'h1 ? dirty_1_46 : _GEN_4298; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4814 = unuse_way == 2'h1 ? dirty_1_47 : _GEN_4299; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4815 = unuse_way == 2'h1 ? dirty_1_48 : _GEN_4300; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4816 = unuse_way == 2'h1 ? dirty_1_49 : _GEN_4301; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4817 = unuse_way == 2'h1 ? dirty_1_50 : _GEN_4302; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4818 = unuse_way == 2'h1 ? dirty_1_51 : _GEN_4303; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4819 = unuse_way == 2'h1 ? dirty_1_52 : _GEN_4304; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4820 = unuse_way == 2'h1 ? dirty_1_53 : _GEN_4305; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4821 = unuse_way == 2'h1 ? dirty_1_54 : _GEN_4306; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4822 = unuse_way == 2'h1 ? dirty_1_55 : _GEN_4307; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4823 = unuse_way == 2'h1 ? dirty_1_56 : _GEN_4308; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4824 = unuse_way == 2'h1 ? dirty_1_57 : _GEN_4309; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4825 = unuse_way == 2'h1 ? dirty_1_58 : _GEN_4310; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4826 = unuse_way == 2'h1 ? dirty_1_59 : _GEN_4311; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4827 = unuse_way == 2'h1 ? dirty_1_60 : _GEN_4312; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4828 = unuse_way == 2'h1 ? dirty_1_61 : _GEN_4313; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4829 = unuse_way == 2'h1 ? dirty_1_62 : _GEN_4314; // @[d_cache.scala 141:34 27:26]
  wire  _GEN_4830 = unuse_way == 2'h1 ? dirty_1_63 : _GEN_4315; // @[d_cache.scala 141:34 27:26]
  wire [2:0] _GEN_4831 = io_from_axi_bvalid ? 3'h7 : state; // @[d_cache.scala 193:37 194:23 76:24]
  wire [2:0] _GEN_4832 = 3'h7 == state ? 3'h1 : state; // @[d_cache.scala 81:18 198:19 76:24]
  wire [2:0] _GEN_4833 = 3'h6 == state ? _GEN_4831 : _GEN_4832; // @[d_cache.scala 81:18]
  wire [2:0] _GEN_4834 = 3'h5 == state ? _GEN_4316 : _GEN_4833; // @[d_cache.scala 81:18]
  wire [63:0] _GEN_4835 = 3'h5 == state ? _GEN_4317 : ram_0_0; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4836 = 3'h5 == state ? _GEN_4318 : ram_0_1; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4837 = 3'h5 == state ? _GEN_4319 : ram_0_2; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4838 = 3'h5 == state ? _GEN_4320 : ram_0_3; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4839 = 3'h5 == state ? _GEN_4321 : ram_0_4; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4840 = 3'h5 == state ? _GEN_4322 : ram_0_5; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4841 = 3'h5 == state ? _GEN_4323 : ram_0_6; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4842 = 3'h5 == state ? _GEN_4324 : ram_0_7; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4843 = 3'h5 == state ? _GEN_4325 : ram_0_8; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4844 = 3'h5 == state ? _GEN_4326 : ram_0_9; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4845 = 3'h5 == state ? _GEN_4327 : ram_0_10; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4846 = 3'h5 == state ? _GEN_4328 : ram_0_11; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4847 = 3'h5 == state ? _GEN_4329 : ram_0_12; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4848 = 3'h5 == state ? _GEN_4330 : ram_0_13; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4849 = 3'h5 == state ? _GEN_4331 : ram_0_14; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4850 = 3'h5 == state ? _GEN_4332 : ram_0_15; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4851 = 3'h5 == state ? _GEN_4333 : ram_0_16; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4852 = 3'h5 == state ? _GEN_4334 : ram_0_17; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4853 = 3'h5 == state ? _GEN_4335 : ram_0_18; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4854 = 3'h5 == state ? _GEN_4336 : ram_0_19; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4855 = 3'h5 == state ? _GEN_4337 : ram_0_20; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4856 = 3'h5 == state ? _GEN_4338 : ram_0_21; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4857 = 3'h5 == state ? _GEN_4339 : ram_0_22; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4858 = 3'h5 == state ? _GEN_4340 : ram_0_23; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4859 = 3'h5 == state ? _GEN_4341 : ram_0_24; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4860 = 3'h5 == state ? _GEN_4342 : ram_0_25; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4861 = 3'h5 == state ? _GEN_4343 : ram_0_26; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4862 = 3'h5 == state ? _GEN_4344 : ram_0_27; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4863 = 3'h5 == state ? _GEN_4345 : ram_0_28; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4864 = 3'h5 == state ? _GEN_4346 : ram_0_29; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4865 = 3'h5 == state ? _GEN_4347 : ram_0_30; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4866 = 3'h5 == state ? _GEN_4348 : ram_0_31; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4867 = 3'h5 == state ? _GEN_4349 : ram_0_32; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4868 = 3'h5 == state ? _GEN_4350 : ram_0_33; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4869 = 3'h5 == state ? _GEN_4351 : ram_0_34; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4870 = 3'h5 == state ? _GEN_4352 : ram_0_35; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4871 = 3'h5 == state ? _GEN_4353 : ram_0_36; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4872 = 3'h5 == state ? _GEN_4354 : ram_0_37; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4873 = 3'h5 == state ? _GEN_4355 : ram_0_38; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4874 = 3'h5 == state ? _GEN_4356 : ram_0_39; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4875 = 3'h5 == state ? _GEN_4357 : ram_0_40; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4876 = 3'h5 == state ? _GEN_4358 : ram_0_41; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4877 = 3'h5 == state ? _GEN_4359 : ram_0_42; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4878 = 3'h5 == state ? _GEN_4360 : ram_0_43; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4879 = 3'h5 == state ? _GEN_4361 : ram_0_44; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4880 = 3'h5 == state ? _GEN_4362 : ram_0_45; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4881 = 3'h5 == state ? _GEN_4363 : ram_0_46; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4882 = 3'h5 == state ? _GEN_4364 : ram_0_47; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4883 = 3'h5 == state ? _GEN_4365 : ram_0_48; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4884 = 3'h5 == state ? _GEN_4366 : ram_0_49; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4885 = 3'h5 == state ? _GEN_4367 : ram_0_50; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4886 = 3'h5 == state ? _GEN_4368 : ram_0_51; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4887 = 3'h5 == state ? _GEN_4369 : ram_0_52; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4888 = 3'h5 == state ? _GEN_4370 : ram_0_53; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4889 = 3'h5 == state ? _GEN_4371 : ram_0_54; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4890 = 3'h5 == state ? _GEN_4372 : ram_0_55; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4891 = 3'h5 == state ? _GEN_4373 : ram_0_56; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4892 = 3'h5 == state ? _GEN_4374 : ram_0_57; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4893 = 3'h5 == state ? _GEN_4375 : ram_0_58; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4894 = 3'h5 == state ? _GEN_4376 : ram_0_59; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4895 = 3'h5 == state ? _GEN_4377 : ram_0_60; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4896 = 3'h5 == state ? _GEN_4378 : ram_0_61; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4897 = 3'h5 == state ? _GEN_4379 : ram_0_62; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_4898 = 3'h5 == state ? _GEN_4380 : ram_0_63; // @[d_cache.scala 81:18 18:24]
  wire [31:0] _GEN_4899 = 3'h5 == state ? _GEN_4381 : tag_0_0; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4900 = 3'h5 == state ? _GEN_4382 : tag_0_1; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4901 = 3'h5 == state ? _GEN_4383 : tag_0_2; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4902 = 3'h5 == state ? _GEN_4384 : tag_0_3; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4903 = 3'h5 == state ? _GEN_4385 : tag_0_4; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4904 = 3'h5 == state ? _GEN_4386 : tag_0_5; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4905 = 3'h5 == state ? _GEN_4387 : tag_0_6; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4906 = 3'h5 == state ? _GEN_4388 : tag_0_7; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4907 = 3'h5 == state ? _GEN_4389 : tag_0_8; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4908 = 3'h5 == state ? _GEN_4390 : tag_0_9; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4909 = 3'h5 == state ? _GEN_4391 : tag_0_10; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4910 = 3'h5 == state ? _GEN_4392 : tag_0_11; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4911 = 3'h5 == state ? _GEN_4393 : tag_0_12; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4912 = 3'h5 == state ? _GEN_4394 : tag_0_13; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4913 = 3'h5 == state ? _GEN_4395 : tag_0_14; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4914 = 3'h5 == state ? _GEN_4396 : tag_0_15; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4915 = 3'h5 == state ? _GEN_4397 : tag_0_16; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4916 = 3'h5 == state ? _GEN_4398 : tag_0_17; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4917 = 3'h5 == state ? _GEN_4399 : tag_0_18; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4918 = 3'h5 == state ? _GEN_4400 : tag_0_19; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4919 = 3'h5 == state ? _GEN_4401 : tag_0_20; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4920 = 3'h5 == state ? _GEN_4402 : tag_0_21; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4921 = 3'h5 == state ? _GEN_4403 : tag_0_22; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4922 = 3'h5 == state ? _GEN_4404 : tag_0_23; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4923 = 3'h5 == state ? _GEN_4405 : tag_0_24; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4924 = 3'h5 == state ? _GEN_4406 : tag_0_25; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4925 = 3'h5 == state ? _GEN_4407 : tag_0_26; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4926 = 3'h5 == state ? _GEN_4408 : tag_0_27; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4927 = 3'h5 == state ? _GEN_4409 : tag_0_28; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4928 = 3'h5 == state ? _GEN_4410 : tag_0_29; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4929 = 3'h5 == state ? _GEN_4411 : tag_0_30; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4930 = 3'h5 == state ? _GEN_4412 : tag_0_31; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4931 = 3'h5 == state ? _GEN_4413 : tag_0_32; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4932 = 3'h5 == state ? _GEN_4414 : tag_0_33; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4933 = 3'h5 == state ? _GEN_4415 : tag_0_34; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4934 = 3'h5 == state ? _GEN_4416 : tag_0_35; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4935 = 3'h5 == state ? _GEN_4417 : tag_0_36; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4936 = 3'h5 == state ? _GEN_4418 : tag_0_37; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4937 = 3'h5 == state ? _GEN_4419 : tag_0_38; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4938 = 3'h5 == state ? _GEN_4420 : tag_0_39; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4939 = 3'h5 == state ? _GEN_4421 : tag_0_40; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4940 = 3'h5 == state ? _GEN_4422 : tag_0_41; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4941 = 3'h5 == state ? _GEN_4423 : tag_0_42; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4942 = 3'h5 == state ? _GEN_4424 : tag_0_43; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4943 = 3'h5 == state ? _GEN_4425 : tag_0_44; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4944 = 3'h5 == state ? _GEN_4426 : tag_0_45; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4945 = 3'h5 == state ? _GEN_4427 : tag_0_46; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4946 = 3'h5 == state ? _GEN_4428 : tag_0_47; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4947 = 3'h5 == state ? _GEN_4429 : tag_0_48; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4948 = 3'h5 == state ? _GEN_4430 : tag_0_49; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4949 = 3'h5 == state ? _GEN_4431 : tag_0_50; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4950 = 3'h5 == state ? _GEN_4432 : tag_0_51; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4951 = 3'h5 == state ? _GEN_4433 : tag_0_52; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4952 = 3'h5 == state ? _GEN_4434 : tag_0_53; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4953 = 3'h5 == state ? _GEN_4435 : tag_0_54; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4954 = 3'h5 == state ? _GEN_4436 : tag_0_55; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4955 = 3'h5 == state ? _GEN_4437 : tag_0_56; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4956 = 3'h5 == state ? _GEN_4438 : tag_0_57; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4957 = 3'h5 == state ? _GEN_4439 : tag_0_58; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4958 = 3'h5 == state ? _GEN_4440 : tag_0_59; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4959 = 3'h5 == state ? _GEN_4441 : tag_0_60; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4960 = 3'h5 == state ? _GEN_4442 : tag_0_61; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4961 = 3'h5 == state ? _GEN_4443 : tag_0_62; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_4962 = 3'h5 == state ? _GEN_4444 : tag_0_63; // @[d_cache.scala 81:18 22:24]
  wire  _GEN_4963 = 3'h5 == state ? _GEN_4445 : valid_0_0; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4964 = 3'h5 == state ? _GEN_4446 : valid_0_1; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4965 = 3'h5 == state ? _GEN_4447 : valid_0_2; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4966 = 3'h5 == state ? _GEN_4448 : valid_0_3; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4967 = 3'h5 == state ? _GEN_4449 : valid_0_4; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4968 = 3'h5 == state ? _GEN_4450 : valid_0_5; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4969 = 3'h5 == state ? _GEN_4451 : valid_0_6; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4970 = 3'h5 == state ? _GEN_4452 : valid_0_7; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4971 = 3'h5 == state ? _GEN_4453 : valid_0_8; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4972 = 3'h5 == state ? _GEN_4454 : valid_0_9; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4973 = 3'h5 == state ? _GEN_4455 : valid_0_10; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4974 = 3'h5 == state ? _GEN_4456 : valid_0_11; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4975 = 3'h5 == state ? _GEN_4457 : valid_0_12; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4976 = 3'h5 == state ? _GEN_4458 : valid_0_13; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4977 = 3'h5 == state ? _GEN_4459 : valid_0_14; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4978 = 3'h5 == state ? _GEN_4460 : valid_0_15; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4979 = 3'h5 == state ? _GEN_4461 : valid_0_16; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4980 = 3'h5 == state ? _GEN_4462 : valid_0_17; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4981 = 3'h5 == state ? _GEN_4463 : valid_0_18; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4982 = 3'h5 == state ? _GEN_4464 : valid_0_19; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4983 = 3'h5 == state ? _GEN_4465 : valid_0_20; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4984 = 3'h5 == state ? _GEN_4466 : valid_0_21; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4985 = 3'h5 == state ? _GEN_4467 : valid_0_22; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4986 = 3'h5 == state ? _GEN_4468 : valid_0_23; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4987 = 3'h5 == state ? _GEN_4469 : valid_0_24; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4988 = 3'h5 == state ? _GEN_4470 : valid_0_25; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4989 = 3'h5 == state ? _GEN_4471 : valid_0_26; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4990 = 3'h5 == state ? _GEN_4472 : valid_0_27; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4991 = 3'h5 == state ? _GEN_4473 : valid_0_28; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4992 = 3'h5 == state ? _GEN_4474 : valid_0_29; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4993 = 3'h5 == state ? _GEN_4475 : valid_0_30; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4994 = 3'h5 == state ? _GEN_4476 : valid_0_31; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4995 = 3'h5 == state ? _GEN_4477 : valid_0_32; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4996 = 3'h5 == state ? _GEN_4478 : valid_0_33; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4997 = 3'h5 == state ? _GEN_4479 : valid_0_34; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4998 = 3'h5 == state ? _GEN_4480 : valid_0_35; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_4999 = 3'h5 == state ? _GEN_4481 : valid_0_36; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5000 = 3'h5 == state ? _GEN_4482 : valid_0_37; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5001 = 3'h5 == state ? _GEN_4483 : valid_0_38; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5002 = 3'h5 == state ? _GEN_4484 : valid_0_39; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5003 = 3'h5 == state ? _GEN_4485 : valid_0_40; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5004 = 3'h5 == state ? _GEN_4486 : valid_0_41; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5005 = 3'h5 == state ? _GEN_4487 : valid_0_42; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5006 = 3'h5 == state ? _GEN_4488 : valid_0_43; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5007 = 3'h5 == state ? _GEN_4489 : valid_0_44; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5008 = 3'h5 == state ? _GEN_4490 : valid_0_45; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5009 = 3'h5 == state ? _GEN_4491 : valid_0_46; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5010 = 3'h5 == state ? _GEN_4492 : valid_0_47; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5011 = 3'h5 == state ? _GEN_4493 : valid_0_48; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5012 = 3'h5 == state ? _GEN_4494 : valid_0_49; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5013 = 3'h5 == state ? _GEN_4495 : valid_0_50; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5014 = 3'h5 == state ? _GEN_4496 : valid_0_51; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5015 = 3'h5 == state ? _GEN_4497 : valid_0_52; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5016 = 3'h5 == state ? _GEN_4498 : valid_0_53; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5017 = 3'h5 == state ? _GEN_4499 : valid_0_54; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5018 = 3'h5 == state ? _GEN_4500 : valid_0_55; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5019 = 3'h5 == state ? _GEN_4501 : valid_0_56; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5020 = 3'h5 == state ? _GEN_4502 : valid_0_57; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5021 = 3'h5 == state ? _GEN_4503 : valid_0_58; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5022 = 3'h5 == state ? _GEN_4504 : valid_0_59; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5023 = 3'h5 == state ? _GEN_4505 : valid_0_60; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5024 = 3'h5 == state ? _GEN_4506 : valid_0_61; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5025 = 3'h5 == state ? _GEN_4507 : valid_0_62; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5026 = 3'h5 == state ? _GEN_4508 : valid_0_63; // @[d_cache.scala 81:18 24:26]
  wire [63:0] _GEN_5027 = 3'h5 == state ? _GEN_4509 : ram_1_0; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5028 = 3'h5 == state ? _GEN_4510 : ram_1_1; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5029 = 3'h5 == state ? _GEN_4511 : ram_1_2; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5030 = 3'h5 == state ? _GEN_4512 : ram_1_3; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5031 = 3'h5 == state ? _GEN_4513 : ram_1_4; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5032 = 3'h5 == state ? _GEN_4514 : ram_1_5; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5033 = 3'h5 == state ? _GEN_4515 : ram_1_6; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5034 = 3'h5 == state ? _GEN_4516 : ram_1_7; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5035 = 3'h5 == state ? _GEN_4517 : ram_1_8; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5036 = 3'h5 == state ? _GEN_4518 : ram_1_9; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5037 = 3'h5 == state ? _GEN_4519 : ram_1_10; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5038 = 3'h5 == state ? _GEN_4520 : ram_1_11; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5039 = 3'h5 == state ? _GEN_4521 : ram_1_12; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5040 = 3'h5 == state ? _GEN_4522 : ram_1_13; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5041 = 3'h5 == state ? _GEN_4523 : ram_1_14; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5042 = 3'h5 == state ? _GEN_4524 : ram_1_15; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5043 = 3'h5 == state ? _GEN_4525 : ram_1_16; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5044 = 3'h5 == state ? _GEN_4526 : ram_1_17; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5045 = 3'h5 == state ? _GEN_4527 : ram_1_18; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5046 = 3'h5 == state ? _GEN_4528 : ram_1_19; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5047 = 3'h5 == state ? _GEN_4529 : ram_1_20; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5048 = 3'h5 == state ? _GEN_4530 : ram_1_21; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5049 = 3'h5 == state ? _GEN_4531 : ram_1_22; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5050 = 3'h5 == state ? _GEN_4532 : ram_1_23; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5051 = 3'h5 == state ? _GEN_4533 : ram_1_24; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5052 = 3'h5 == state ? _GEN_4534 : ram_1_25; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5053 = 3'h5 == state ? _GEN_4535 : ram_1_26; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5054 = 3'h5 == state ? _GEN_4536 : ram_1_27; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5055 = 3'h5 == state ? _GEN_4537 : ram_1_28; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5056 = 3'h5 == state ? _GEN_4538 : ram_1_29; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5057 = 3'h5 == state ? _GEN_4539 : ram_1_30; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5058 = 3'h5 == state ? _GEN_4540 : ram_1_31; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5059 = 3'h5 == state ? _GEN_4541 : ram_1_32; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5060 = 3'h5 == state ? _GEN_4542 : ram_1_33; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5061 = 3'h5 == state ? _GEN_4543 : ram_1_34; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5062 = 3'h5 == state ? _GEN_4544 : ram_1_35; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5063 = 3'h5 == state ? _GEN_4545 : ram_1_36; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5064 = 3'h5 == state ? _GEN_4546 : ram_1_37; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5065 = 3'h5 == state ? _GEN_4547 : ram_1_38; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5066 = 3'h5 == state ? _GEN_4548 : ram_1_39; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5067 = 3'h5 == state ? _GEN_4549 : ram_1_40; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5068 = 3'h5 == state ? _GEN_4550 : ram_1_41; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5069 = 3'h5 == state ? _GEN_4551 : ram_1_42; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5070 = 3'h5 == state ? _GEN_4552 : ram_1_43; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5071 = 3'h5 == state ? _GEN_4553 : ram_1_44; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5072 = 3'h5 == state ? _GEN_4554 : ram_1_45; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5073 = 3'h5 == state ? _GEN_4555 : ram_1_46; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5074 = 3'h5 == state ? _GEN_4556 : ram_1_47; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5075 = 3'h5 == state ? _GEN_4557 : ram_1_48; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5076 = 3'h5 == state ? _GEN_4558 : ram_1_49; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5077 = 3'h5 == state ? _GEN_4559 : ram_1_50; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5078 = 3'h5 == state ? _GEN_4560 : ram_1_51; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5079 = 3'h5 == state ? _GEN_4561 : ram_1_52; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5080 = 3'h5 == state ? _GEN_4562 : ram_1_53; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5081 = 3'h5 == state ? _GEN_4563 : ram_1_54; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5082 = 3'h5 == state ? _GEN_4564 : ram_1_55; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5083 = 3'h5 == state ? _GEN_4565 : ram_1_56; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5084 = 3'h5 == state ? _GEN_4566 : ram_1_57; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5085 = 3'h5 == state ? _GEN_4567 : ram_1_58; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5086 = 3'h5 == state ? _GEN_4568 : ram_1_59; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5087 = 3'h5 == state ? _GEN_4569 : ram_1_60; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5088 = 3'h5 == state ? _GEN_4570 : ram_1_61; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5089 = 3'h5 == state ? _GEN_4571 : ram_1_62; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5090 = 3'h5 == state ? _GEN_4572 : ram_1_63; // @[d_cache.scala 81:18 19:24]
  wire [31:0] _GEN_5091 = 3'h5 == state ? _GEN_4573 : tag_1_0; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5092 = 3'h5 == state ? _GEN_4574 : tag_1_1; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5093 = 3'h5 == state ? _GEN_4575 : tag_1_2; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5094 = 3'h5 == state ? _GEN_4576 : tag_1_3; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5095 = 3'h5 == state ? _GEN_4577 : tag_1_4; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5096 = 3'h5 == state ? _GEN_4578 : tag_1_5; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5097 = 3'h5 == state ? _GEN_4579 : tag_1_6; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5098 = 3'h5 == state ? _GEN_4580 : tag_1_7; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5099 = 3'h5 == state ? _GEN_4581 : tag_1_8; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5100 = 3'h5 == state ? _GEN_4582 : tag_1_9; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5101 = 3'h5 == state ? _GEN_4583 : tag_1_10; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5102 = 3'h5 == state ? _GEN_4584 : tag_1_11; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5103 = 3'h5 == state ? _GEN_4585 : tag_1_12; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5104 = 3'h5 == state ? _GEN_4586 : tag_1_13; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5105 = 3'h5 == state ? _GEN_4587 : tag_1_14; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5106 = 3'h5 == state ? _GEN_4588 : tag_1_15; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5107 = 3'h5 == state ? _GEN_4589 : tag_1_16; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5108 = 3'h5 == state ? _GEN_4590 : tag_1_17; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5109 = 3'h5 == state ? _GEN_4591 : tag_1_18; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5110 = 3'h5 == state ? _GEN_4592 : tag_1_19; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5111 = 3'h5 == state ? _GEN_4593 : tag_1_20; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5112 = 3'h5 == state ? _GEN_4594 : tag_1_21; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5113 = 3'h5 == state ? _GEN_4595 : tag_1_22; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5114 = 3'h5 == state ? _GEN_4596 : tag_1_23; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5115 = 3'h5 == state ? _GEN_4597 : tag_1_24; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5116 = 3'h5 == state ? _GEN_4598 : tag_1_25; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5117 = 3'h5 == state ? _GEN_4599 : tag_1_26; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5118 = 3'h5 == state ? _GEN_4600 : tag_1_27; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5119 = 3'h5 == state ? _GEN_4601 : tag_1_28; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5120 = 3'h5 == state ? _GEN_4602 : tag_1_29; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5121 = 3'h5 == state ? _GEN_4603 : tag_1_30; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5122 = 3'h5 == state ? _GEN_4604 : tag_1_31; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5123 = 3'h5 == state ? _GEN_4605 : tag_1_32; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5124 = 3'h5 == state ? _GEN_4606 : tag_1_33; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5125 = 3'h5 == state ? _GEN_4607 : tag_1_34; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5126 = 3'h5 == state ? _GEN_4608 : tag_1_35; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5127 = 3'h5 == state ? _GEN_4609 : tag_1_36; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5128 = 3'h5 == state ? _GEN_4610 : tag_1_37; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5129 = 3'h5 == state ? _GEN_4611 : tag_1_38; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5130 = 3'h5 == state ? _GEN_4612 : tag_1_39; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5131 = 3'h5 == state ? _GEN_4613 : tag_1_40; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5132 = 3'h5 == state ? _GEN_4614 : tag_1_41; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5133 = 3'h5 == state ? _GEN_4615 : tag_1_42; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5134 = 3'h5 == state ? _GEN_4616 : tag_1_43; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5135 = 3'h5 == state ? _GEN_4617 : tag_1_44; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5136 = 3'h5 == state ? _GEN_4618 : tag_1_45; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5137 = 3'h5 == state ? _GEN_4619 : tag_1_46; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5138 = 3'h5 == state ? _GEN_4620 : tag_1_47; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5139 = 3'h5 == state ? _GEN_4621 : tag_1_48; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5140 = 3'h5 == state ? _GEN_4622 : tag_1_49; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5141 = 3'h5 == state ? _GEN_4623 : tag_1_50; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5142 = 3'h5 == state ? _GEN_4624 : tag_1_51; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5143 = 3'h5 == state ? _GEN_4625 : tag_1_52; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5144 = 3'h5 == state ? _GEN_4626 : tag_1_53; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5145 = 3'h5 == state ? _GEN_4627 : tag_1_54; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5146 = 3'h5 == state ? _GEN_4628 : tag_1_55; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5147 = 3'h5 == state ? _GEN_4629 : tag_1_56; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5148 = 3'h5 == state ? _GEN_4630 : tag_1_57; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5149 = 3'h5 == state ? _GEN_4631 : tag_1_58; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5150 = 3'h5 == state ? _GEN_4632 : tag_1_59; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5151 = 3'h5 == state ? _GEN_4633 : tag_1_60; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5152 = 3'h5 == state ? _GEN_4634 : tag_1_61; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5153 = 3'h5 == state ? _GEN_4635 : tag_1_62; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5154 = 3'h5 == state ? _GEN_4636 : tag_1_63; // @[d_cache.scala 81:18 23:24]
  wire  _GEN_5155 = 3'h5 == state ? _GEN_4637 : valid_1_0; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5156 = 3'h5 == state ? _GEN_4638 : valid_1_1; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5157 = 3'h5 == state ? _GEN_4639 : valid_1_2; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5158 = 3'h5 == state ? _GEN_4640 : valid_1_3; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5159 = 3'h5 == state ? _GEN_4641 : valid_1_4; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5160 = 3'h5 == state ? _GEN_4642 : valid_1_5; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5161 = 3'h5 == state ? _GEN_4643 : valid_1_6; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5162 = 3'h5 == state ? _GEN_4644 : valid_1_7; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5163 = 3'h5 == state ? _GEN_4645 : valid_1_8; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5164 = 3'h5 == state ? _GEN_4646 : valid_1_9; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5165 = 3'h5 == state ? _GEN_4647 : valid_1_10; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5166 = 3'h5 == state ? _GEN_4648 : valid_1_11; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5167 = 3'h5 == state ? _GEN_4649 : valid_1_12; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5168 = 3'h5 == state ? _GEN_4650 : valid_1_13; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5169 = 3'h5 == state ? _GEN_4651 : valid_1_14; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5170 = 3'h5 == state ? _GEN_4652 : valid_1_15; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5171 = 3'h5 == state ? _GEN_4653 : valid_1_16; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5172 = 3'h5 == state ? _GEN_4654 : valid_1_17; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5173 = 3'h5 == state ? _GEN_4655 : valid_1_18; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5174 = 3'h5 == state ? _GEN_4656 : valid_1_19; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5175 = 3'h5 == state ? _GEN_4657 : valid_1_20; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5176 = 3'h5 == state ? _GEN_4658 : valid_1_21; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5177 = 3'h5 == state ? _GEN_4659 : valid_1_22; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5178 = 3'h5 == state ? _GEN_4660 : valid_1_23; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5179 = 3'h5 == state ? _GEN_4661 : valid_1_24; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5180 = 3'h5 == state ? _GEN_4662 : valid_1_25; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5181 = 3'h5 == state ? _GEN_4663 : valid_1_26; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5182 = 3'h5 == state ? _GEN_4664 : valid_1_27; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5183 = 3'h5 == state ? _GEN_4665 : valid_1_28; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5184 = 3'h5 == state ? _GEN_4666 : valid_1_29; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5185 = 3'h5 == state ? _GEN_4667 : valid_1_30; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5186 = 3'h5 == state ? _GEN_4668 : valid_1_31; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5187 = 3'h5 == state ? _GEN_4669 : valid_1_32; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5188 = 3'h5 == state ? _GEN_4670 : valid_1_33; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5189 = 3'h5 == state ? _GEN_4671 : valid_1_34; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5190 = 3'h5 == state ? _GEN_4672 : valid_1_35; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5191 = 3'h5 == state ? _GEN_4673 : valid_1_36; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5192 = 3'h5 == state ? _GEN_4674 : valid_1_37; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5193 = 3'h5 == state ? _GEN_4675 : valid_1_38; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5194 = 3'h5 == state ? _GEN_4676 : valid_1_39; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5195 = 3'h5 == state ? _GEN_4677 : valid_1_40; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5196 = 3'h5 == state ? _GEN_4678 : valid_1_41; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5197 = 3'h5 == state ? _GEN_4679 : valid_1_42; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5198 = 3'h5 == state ? _GEN_4680 : valid_1_43; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5199 = 3'h5 == state ? _GEN_4681 : valid_1_44; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5200 = 3'h5 == state ? _GEN_4682 : valid_1_45; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5201 = 3'h5 == state ? _GEN_4683 : valid_1_46; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5202 = 3'h5 == state ? _GEN_4684 : valid_1_47; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5203 = 3'h5 == state ? _GEN_4685 : valid_1_48; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5204 = 3'h5 == state ? _GEN_4686 : valid_1_49; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5205 = 3'h5 == state ? _GEN_4687 : valid_1_50; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5206 = 3'h5 == state ? _GEN_4688 : valid_1_51; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5207 = 3'h5 == state ? _GEN_4689 : valid_1_52; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5208 = 3'h5 == state ? _GEN_4690 : valid_1_53; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5209 = 3'h5 == state ? _GEN_4691 : valid_1_54; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5210 = 3'h5 == state ? _GEN_4692 : valid_1_55; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5211 = 3'h5 == state ? _GEN_4693 : valid_1_56; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5212 = 3'h5 == state ? _GEN_4694 : valid_1_57; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5213 = 3'h5 == state ? _GEN_4695 : valid_1_58; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5214 = 3'h5 == state ? _GEN_4696 : valid_1_59; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5215 = 3'h5 == state ? _GEN_4697 : valid_1_60; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5216 = 3'h5 == state ? _GEN_4698 : valid_1_61; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5217 = 3'h5 == state ? _GEN_4699 : valid_1_62; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5218 = 3'h5 == state ? _GEN_4700 : valid_1_63; // @[d_cache.scala 81:18 25:26]
  wire [63:0] _GEN_5219 = 3'h5 == state ? _GEN_4701 : write_back_data; // @[d_cache.scala 81:18 31:34]
  wire [40:0] _GEN_5220 = 3'h5 == state ? _GEN_4702 : {{9'd0}, write_back_addr}; // @[d_cache.scala 81:18 32:34]
  wire  _GEN_5221 = 3'h5 == state ? _GEN_4703 : dirty_0_0; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5222 = 3'h5 == state ? _GEN_4704 : dirty_0_1; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5223 = 3'h5 == state ? _GEN_4705 : dirty_0_2; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5224 = 3'h5 == state ? _GEN_4706 : dirty_0_3; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5225 = 3'h5 == state ? _GEN_4707 : dirty_0_4; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5226 = 3'h5 == state ? _GEN_4708 : dirty_0_5; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5227 = 3'h5 == state ? _GEN_4709 : dirty_0_6; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5228 = 3'h5 == state ? _GEN_4710 : dirty_0_7; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5229 = 3'h5 == state ? _GEN_4711 : dirty_0_8; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5230 = 3'h5 == state ? _GEN_4712 : dirty_0_9; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5231 = 3'h5 == state ? _GEN_4713 : dirty_0_10; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5232 = 3'h5 == state ? _GEN_4714 : dirty_0_11; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5233 = 3'h5 == state ? _GEN_4715 : dirty_0_12; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5234 = 3'h5 == state ? _GEN_4716 : dirty_0_13; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5235 = 3'h5 == state ? _GEN_4717 : dirty_0_14; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5236 = 3'h5 == state ? _GEN_4718 : dirty_0_15; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5237 = 3'h5 == state ? _GEN_4719 : dirty_0_16; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5238 = 3'h5 == state ? _GEN_4720 : dirty_0_17; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5239 = 3'h5 == state ? _GEN_4721 : dirty_0_18; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5240 = 3'h5 == state ? _GEN_4722 : dirty_0_19; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5241 = 3'h5 == state ? _GEN_4723 : dirty_0_20; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5242 = 3'h5 == state ? _GEN_4724 : dirty_0_21; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5243 = 3'h5 == state ? _GEN_4725 : dirty_0_22; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5244 = 3'h5 == state ? _GEN_4726 : dirty_0_23; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5245 = 3'h5 == state ? _GEN_4727 : dirty_0_24; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5246 = 3'h5 == state ? _GEN_4728 : dirty_0_25; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5247 = 3'h5 == state ? _GEN_4729 : dirty_0_26; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5248 = 3'h5 == state ? _GEN_4730 : dirty_0_27; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5249 = 3'h5 == state ? _GEN_4731 : dirty_0_28; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5250 = 3'h5 == state ? _GEN_4732 : dirty_0_29; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5251 = 3'h5 == state ? _GEN_4733 : dirty_0_30; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5252 = 3'h5 == state ? _GEN_4734 : dirty_0_31; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5253 = 3'h5 == state ? _GEN_4735 : dirty_0_32; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5254 = 3'h5 == state ? _GEN_4736 : dirty_0_33; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5255 = 3'h5 == state ? _GEN_4737 : dirty_0_34; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5256 = 3'h5 == state ? _GEN_4738 : dirty_0_35; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5257 = 3'h5 == state ? _GEN_4739 : dirty_0_36; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5258 = 3'h5 == state ? _GEN_4740 : dirty_0_37; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5259 = 3'h5 == state ? _GEN_4741 : dirty_0_38; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5260 = 3'h5 == state ? _GEN_4742 : dirty_0_39; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5261 = 3'h5 == state ? _GEN_4743 : dirty_0_40; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5262 = 3'h5 == state ? _GEN_4744 : dirty_0_41; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5263 = 3'h5 == state ? _GEN_4745 : dirty_0_42; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5264 = 3'h5 == state ? _GEN_4746 : dirty_0_43; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5265 = 3'h5 == state ? _GEN_4747 : dirty_0_44; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5266 = 3'h5 == state ? _GEN_4748 : dirty_0_45; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5267 = 3'h5 == state ? _GEN_4749 : dirty_0_46; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5268 = 3'h5 == state ? _GEN_4750 : dirty_0_47; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5269 = 3'h5 == state ? _GEN_4751 : dirty_0_48; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5270 = 3'h5 == state ? _GEN_4752 : dirty_0_49; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5271 = 3'h5 == state ? _GEN_4753 : dirty_0_50; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5272 = 3'h5 == state ? _GEN_4754 : dirty_0_51; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5273 = 3'h5 == state ? _GEN_4755 : dirty_0_52; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5274 = 3'h5 == state ? _GEN_4756 : dirty_0_53; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5275 = 3'h5 == state ? _GEN_4757 : dirty_0_54; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5276 = 3'h5 == state ? _GEN_4758 : dirty_0_55; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5277 = 3'h5 == state ? _GEN_4759 : dirty_0_56; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5278 = 3'h5 == state ? _GEN_4760 : dirty_0_57; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5279 = 3'h5 == state ? _GEN_4761 : dirty_0_58; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5280 = 3'h5 == state ? _GEN_4762 : dirty_0_59; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5281 = 3'h5 == state ? _GEN_4763 : dirty_0_60; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5282 = 3'h5 == state ? _GEN_4764 : dirty_0_61; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5283 = 3'h5 == state ? _GEN_4765 : dirty_0_62; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5284 = 3'h5 == state ? _GEN_4766 : dirty_0_63; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5285 = 3'h5 == state ? _GEN_4767 : dirty_1_0; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5286 = 3'h5 == state ? _GEN_4768 : dirty_1_1; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5287 = 3'h5 == state ? _GEN_4769 : dirty_1_2; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5288 = 3'h5 == state ? _GEN_4770 : dirty_1_3; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5289 = 3'h5 == state ? _GEN_4771 : dirty_1_4; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5290 = 3'h5 == state ? _GEN_4772 : dirty_1_5; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5291 = 3'h5 == state ? _GEN_4773 : dirty_1_6; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5292 = 3'h5 == state ? _GEN_4774 : dirty_1_7; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5293 = 3'h5 == state ? _GEN_4775 : dirty_1_8; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5294 = 3'h5 == state ? _GEN_4776 : dirty_1_9; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5295 = 3'h5 == state ? _GEN_4777 : dirty_1_10; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5296 = 3'h5 == state ? _GEN_4778 : dirty_1_11; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5297 = 3'h5 == state ? _GEN_4779 : dirty_1_12; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5298 = 3'h5 == state ? _GEN_4780 : dirty_1_13; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5299 = 3'h5 == state ? _GEN_4781 : dirty_1_14; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5300 = 3'h5 == state ? _GEN_4782 : dirty_1_15; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5301 = 3'h5 == state ? _GEN_4783 : dirty_1_16; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5302 = 3'h5 == state ? _GEN_4784 : dirty_1_17; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5303 = 3'h5 == state ? _GEN_4785 : dirty_1_18; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5304 = 3'h5 == state ? _GEN_4786 : dirty_1_19; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5305 = 3'h5 == state ? _GEN_4787 : dirty_1_20; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5306 = 3'h5 == state ? _GEN_4788 : dirty_1_21; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5307 = 3'h5 == state ? _GEN_4789 : dirty_1_22; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5308 = 3'h5 == state ? _GEN_4790 : dirty_1_23; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5309 = 3'h5 == state ? _GEN_4791 : dirty_1_24; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5310 = 3'h5 == state ? _GEN_4792 : dirty_1_25; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5311 = 3'h5 == state ? _GEN_4793 : dirty_1_26; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5312 = 3'h5 == state ? _GEN_4794 : dirty_1_27; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5313 = 3'h5 == state ? _GEN_4795 : dirty_1_28; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5314 = 3'h5 == state ? _GEN_4796 : dirty_1_29; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5315 = 3'h5 == state ? _GEN_4797 : dirty_1_30; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5316 = 3'h5 == state ? _GEN_4798 : dirty_1_31; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5317 = 3'h5 == state ? _GEN_4799 : dirty_1_32; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5318 = 3'h5 == state ? _GEN_4800 : dirty_1_33; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5319 = 3'h5 == state ? _GEN_4801 : dirty_1_34; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5320 = 3'h5 == state ? _GEN_4802 : dirty_1_35; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5321 = 3'h5 == state ? _GEN_4803 : dirty_1_36; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5322 = 3'h5 == state ? _GEN_4804 : dirty_1_37; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5323 = 3'h5 == state ? _GEN_4805 : dirty_1_38; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5324 = 3'h5 == state ? _GEN_4806 : dirty_1_39; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5325 = 3'h5 == state ? _GEN_4807 : dirty_1_40; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5326 = 3'h5 == state ? _GEN_4808 : dirty_1_41; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5327 = 3'h5 == state ? _GEN_4809 : dirty_1_42; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5328 = 3'h5 == state ? _GEN_4810 : dirty_1_43; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5329 = 3'h5 == state ? _GEN_4811 : dirty_1_44; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5330 = 3'h5 == state ? _GEN_4812 : dirty_1_45; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5331 = 3'h5 == state ? _GEN_4813 : dirty_1_46; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5332 = 3'h5 == state ? _GEN_4814 : dirty_1_47; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5333 = 3'h5 == state ? _GEN_4815 : dirty_1_48; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5334 = 3'h5 == state ? _GEN_4816 : dirty_1_49; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5335 = 3'h5 == state ? _GEN_4817 : dirty_1_50; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5336 = 3'h5 == state ? _GEN_4818 : dirty_1_51; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5337 = 3'h5 == state ? _GEN_4819 : dirty_1_52; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5338 = 3'h5 == state ? _GEN_4820 : dirty_1_53; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5339 = 3'h5 == state ? _GEN_4821 : dirty_1_54; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5340 = 3'h5 == state ? _GEN_4822 : dirty_1_55; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5341 = 3'h5 == state ? _GEN_4823 : dirty_1_56; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5342 = 3'h5 == state ? _GEN_4824 : dirty_1_57; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5343 = 3'h5 == state ? _GEN_4825 : dirty_1_58; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5344 = 3'h5 == state ? _GEN_4826 : dirty_1_59; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5345 = 3'h5 == state ? _GEN_4827 : dirty_1_60; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5346 = 3'h5 == state ? _GEN_4828 : dirty_1_61; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5347 = 3'h5 == state ? _GEN_4829 : dirty_1_62; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5348 = 3'h5 == state ? _GEN_4830 : dirty_1_63; // @[d_cache.scala 81:18 27:26]
  wire [2:0] _GEN_5349 = 3'h4 == state ? _GEN_1487 : _GEN_4834; // @[d_cache.scala 81:18]
  wire [63:0] _GEN_5350 = 3'h4 == state ? ram_0_0 : _GEN_4835; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5351 = 3'h4 == state ? ram_0_1 : _GEN_4836; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5352 = 3'h4 == state ? ram_0_2 : _GEN_4837; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5353 = 3'h4 == state ? ram_0_3 : _GEN_4838; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5354 = 3'h4 == state ? ram_0_4 : _GEN_4839; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5355 = 3'h4 == state ? ram_0_5 : _GEN_4840; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5356 = 3'h4 == state ? ram_0_6 : _GEN_4841; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5357 = 3'h4 == state ? ram_0_7 : _GEN_4842; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5358 = 3'h4 == state ? ram_0_8 : _GEN_4843; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5359 = 3'h4 == state ? ram_0_9 : _GEN_4844; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5360 = 3'h4 == state ? ram_0_10 : _GEN_4845; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5361 = 3'h4 == state ? ram_0_11 : _GEN_4846; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5362 = 3'h4 == state ? ram_0_12 : _GEN_4847; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5363 = 3'h4 == state ? ram_0_13 : _GEN_4848; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5364 = 3'h4 == state ? ram_0_14 : _GEN_4849; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5365 = 3'h4 == state ? ram_0_15 : _GEN_4850; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5366 = 3'h4 == state ? ram_0_16 : _GEN_4851; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5367 = 3'h4 == state ? ram_0_17 : _GEN_4852; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5368 = 3'h4 == state ? ram_0_18 : _GEN_4853; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5369 = 3'h4 == state ? ram_0_19 : _GEN_4854; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5370 = 3'h4 == state ? ram_0_20 : _GEN_4855; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5371 = 3'h4 == state ? ram_0_21 : _GEN_4856; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5372 = 3'h4 == state ? ram_0_22 : _GEN_4857; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5373 = 3'h4 == state ? ram_0_23 : _GEN_4858; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5374 = 3'h4 == state ? ram_0_24 : _GEN_4859; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5375 = 3'h4 == state ? ram_0_25 : _GEN_4860; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5376 = 3'h4 == state ? ram_0_26 : _GEN_4861; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5377 = 3'h4 == state ? ram_0_27 : _GEN_4862; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5378 = 3'h4 == state ? ram_0_28 : _GEN_4863; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5379 = 3'h4 == state ? ram_0_29 : _GEN_4864; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5380 = 3'h4 == state ? ram_0_30 : _GEN_4865; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5381 = 3'h4 == state ? ram_0_31 : _GEN_4866; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5382 = 3'h4 == state ? ram_0_32 : _GEN_4867; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5383 = 3'h4 == state ? ram_0_33 : _GEN_4868; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5384 = 3'h4 == state ? ram_0_34 : _GEN_4869; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5385 = 3'h4 == state ? ram_0_35 : _GEN_4870; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5386 = 3'h4 == state ? ram_0_36 : _GEN_4871; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5387 = 3'h4 == state ? ram_0_37 : _GEN_4872; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5388 = 3'h4 == state ? ram_0_38 : _GEN_4873; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5389 = 3'h4 == state ? ram_0_39 : _GEN_4874; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5390 = 3'h4 == state ? ram_0_40 : _GEN_4875; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5391 = 3'h4 == state ? ram_0_41 : _GEN_4876; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5392 = 3'h4 == state ? ram_0_42 : _GEN_4877; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5393 = 3'h4 == state ? ram_0_43 : _GEN_4878; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5394 = 3'h4 == state ? ram_0_44 : _GEN_4879; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5395 = 3'h4 == state ? ram_0_45 : _GEN_4880; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5396 = 3'h4 == state ? ram_0_46 : _GEN_4881; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5397 = 3'h4 == state ? ram_0_47 : _GEN_4882; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5398 = 3'h4 == state ? ram_0_48 : _GEN_4883; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5399 = 3'h4 == state ? ram_0_49 : _GEN_4884; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5400 = 3'h4 == state ? ram_0_50 : _GEN_4885; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5401 = 3'h4 == state ? ram_0_51 : _GEN_4886; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5402 = 3'h4 == state ? ram_0_52 : _GEN_4887; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5403 = 3'h4 == state ? ram_0_53 : _GEN_4888; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5404 = 3'h4 == state ? ram_0_54 : _GEN_4889; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5405 = 3'h4 == state ? ram_0_55 : _GEN_4890; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5406 = 3'h4 == state ? ram_0_56 : _GEN_4891; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5407 = 3'h4 == state ? ram_0_57 : _GEN_4892; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5408 = 3'h4 == state ? ram_0_58 : _GEN_4893; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5409 = 3'h4 == state ? ram_0_59 : _GEN_4894; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5410 = 3'h4 == state ? ram_0_60 : _GEN_4895; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5411 = 3'h4 == state ? ram_0_61 : _GEN_4896; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5412 = 3'h4 == state ? ram_0_62 : _GEN_4897; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5413 = 3'h4 == state ? ram_0_63 : _GEN_4898; // @[d_cache.scala 81:18 18:24]
  wire [31:0] _GEN_5414 = 3'h4 == state ? tag_0_0 : _GEN_4899; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5415 = 3'h4 == state ? tag_0_1 : _GEN_4900; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5416 = 3'h4 == state ? tag_0_2 : _GEN_4901; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5417 = 3'h4 == state ? tag_0_3 : _GEN_4902; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5418 = 3'h4 == state ? tag_0_4 : _GEN_4903; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5419 = 3'h4 == state ? tag_0_5 : _GEN_4904; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5420 = 3'h4 == state ? tag_0_6 : _GEN_4905; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5421 = 3'h4 == state ? tag_0_7 : _GEN_4906; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5422 = 3'h4 == state ? tag_0_8 : _GEN_4907; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5423 = 3'h4 == state ? tag_0_9 : _GEN_4908; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5424 = 3'h4 == state ? tag_0_10 : _GEN_4909; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5425 = 3'h4 == state ? tag_0_11 : _GEN_4910; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5426 = 3'h4 == state ? tag_0_12 : _GEN_4911; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5427 = 3'h4 == state ? tag_0_13 : _GEN_4912; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5428 = 3'h4 == state ? tag_0_14 : _GEN_4913; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5429 = 3'h4 == state ? tag_0_15 : _GEN_4914; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5430 = 3'h4 == state ? tag_0_16 : _GEN_4915; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5431 = 3'h4 == state ? tag_0_17 : _GEN_4916; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5432 = 3'h4 == state ? tag_0_18 : _GEN_4917; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5433 = 3'h4 == state ? tag_0_19 : _GEN_4918; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5434 = 3'h4 == state ? tag_0_20 : _GEN_4919; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5435 = 3'h4 == state ? tag_0_21 : _GEN_4920; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5436 = 3'h4 == state ? tag_0_22 : _GEN_4921; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5437 = 3'h4 == state ? tag_0_23 : _GEN_4922; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5438 = 3'h4 == state ? tag_0_24 : _GEN_4923; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5439 = 3'h4 == state ? tag_0_25 : _GEN_4924; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5440 = 3'h4 == state ? tag_0_26 : _GEN_4925; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5441 = 3'h4 == state ? tag_0_27 : _GEN_4926; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5442 = 3'h4 == state ? tag_0_28 : _GEN_4927; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5443 = 3'h4 == state ? tag_0_29 : _GEN_4928; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5444 = 3'h4 == state ? tag_0_30 : _GEN_4929; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5445 = 3'h4 == state ? tag_0_31 : _GEN_4930; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5446 = 3'h4 == state ? tag_0_32 : _GEN_4931; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5447 = 3'h4 == state ? tag_0_33 : _GEN_4932; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5448 = 3'h4 == state ? tag_0_34 : _GEN_4933; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5449 = 3'h4 == state ? tag_0_35 : _GEN_4934; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5450 = 3'h4 == state ? tag_0_36 : _GEN_4935; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5451 = 3'h4 == state ? tag_0_37 : _GEN_4936; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5452 = 3'h4 == state ? tag_0_38 : _GEN_4937; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5453 = 3'h4 == state ? tag_0_39 : _GEN_4938; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5454 = 3'h4 == state ? tag_0_40 : _GEN_4939; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5455 = 3'h4 == state ? tag_0_41 : _GEN_4940; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5456 = 3'h4 == state ? tag_0_42 : _GEN_4941; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5457 = 3'h4 == state ? tag_0_43 : _GEN_4942; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5458 = 3'h4 == state ? tag_0_44 : _GEN_4943; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5459 = 3'h4 == state ? tag_0_45 : _GEN_4944; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5460 = 3'h4 == state ? tag_0_46 : _GEN_4945; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5461 = 3'h4 == state ? tag_0_47 : _GEN_4946; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5462 = 3'h4 == state ? tag_0_48 : _GEN_4947; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5463 = 3'h4 == state ? tag_0_49 : _GEN_4948; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5464 = 3'h4 == state ? tag_0_50 : _GEN_4949; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5465 = 3'h4 == state ? tag_0_51 : _GEN_4950; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5466 = 3'h4 == state ? tag_0_52 : _GEN_4951; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5467 = 3'h4 == state ? tag_0_53 : _GEN_4952; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5468 = 3'h4 == state ? tag_0_54 : _GEN_4953; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5469 = 3'h4 == state ? tag_0_55 : _GEN_4954; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5470 = 3'h4 == state ? tag_0_56 : _GEN_4955; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5471 = 3'h4 == state ? tag_0_57 : _GEN_4956; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5472 = 3'h4 == state ? tag_0_58 : _GEN_4957; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5473 = 3'h4 == state ? tag_0_59 : _GEN_4958; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5474 = 3'h4 == state ? tag_0_60 : _GEN_4959; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5475 = 3'h4 == state ? tag_0_61 : _GEN_4960; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5476 = 3'h4 == state ? tag_0_62 : _GEN_4961; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5477 = 3'h4 == state ? tag_0_63 : _GEN_4962; // @[d_cache.scala 81:18 22:24]
  wire  _GEN_5478 = 3'h4 == state ? valid_0_0 : _GEN_4963; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5479 = 3'h4 == state ? valid_0_1 : _GEN_4964; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5480 = 3'h4 == state ? valid_0_2 : _GEN_4965; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5481 = 3'h4 == state ? valid_0_3 : _GEN_4966; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5482 = 3'h4 == state ? valid_0_4 : _GEN_4967; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5483 = 3'h4 == state ? valid_0_5 : _GEN_4968; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5484 = 3'h4 == state ? valid_0_6 : _GEN_4969; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5485 = 3'h4 == state ? valid_0_7 : _GEN_4970; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5486 = 3'h4 == state ? valid_0_8 : _GEN_4971; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5487 = 3'h4 == state ? valid_0_9 : _GEN_4972; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5488 = 3'h4 == state ? valid_0_10 : _GEN_4973; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5489 = 3'h4 == state ? valid_0_11 : _GEN_4974; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5490 = 3'h4 == state ? valid_0_12 : _GEN_4975; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5491 = 3'h4 == state ? valid_0_13 : _GEN_4976; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5492 = 3'h4 == state ? valid_0_14 : _GEN_4977; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5493 = 3'h4 == state ? valid_0_15 : _GEN_4978; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5494 = 3'h4 == state ? valid_0_16 : _GEN_4979; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5495 = 3'h4 == state ? valid_0_17 : _GEN_4980; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5496 = 3'h4 == state ? valid_0_18 : _GEN_4981; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5497 = 3'h4 == state ? valid_0_19 : _GEN_4982; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5498 = 3'h4 == state ? valid_0_20 : _GEN_4983; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5499 = 3'h4 == state ? valid_0_21 : _GEN_4984; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5500 = 3'h4 == state ? valid_0_22 : _GEN_4985; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5501 = 3'h4 == state ? valid_0_23 : _GEN_4986; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5502 = 3'h4 == state ? valid_0_24 : _GEN_4987; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5503 = 3'h4 == state ? valid_0_25 : _GEN_4988; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5504 = 3'h4 == state ? valid_0_26 : _GEN_4989; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5505 = 3'h4 == state ? valid_0_27 : _GEN_4990; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5506 = 3'h4 == state ? valid_0_28 : _GEN_4991; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5507 = 3'h4 == state ? valid_0_29 : _GEN_4992; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5508 = 3'h4 == state ? valid_0_30 : _GEN_4993; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5509 = 3'h4 == state ? valid_0_31 : _GEN_4994; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5510 = 3'h4 == state ? valid_0_32 : _GEN_4995; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5511 = 3'h4 == state ? valid_0_33 : _GEN_4996; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5512 = 3'h4 == state ? valid_0_34 : _GEN_4997; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5513 = 3'h4 == state ? valid_0_35 : _GEN_4998; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5514 = 3'h4 == state ? valid_0_36 : _GEN_4999; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5515 = 3'h4 == state ? valid_0_37 : _GEN_5000; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5516 = 3'h4 == state ? valid_0_38 : _GEN_5001; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5517 = 3'h4 == state ? valid_0_39 : _GEN_5002; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5518 = 3'h4 == state ? valid_0_40 : _GEN_5003; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5519 = 3'h4 == state ? valid_0_41 : _GEN_5004; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5520 = 3'h4 == state ? valid_0_42 : _GEN_5005; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5521 = 3'h4 == state ? valid_0_43 : _GEN_5006; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5522 = 3'h4 == state ? valid_0_44 : _GEN_5007; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5523 = 3'h4 == state ? valid_0_45 : _GEN_5008; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5524 = 3'h4 == state ? valid_0_46 : _GEN_5009; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5525 = 3'h4 == state ? valid_0_47 : _GEN_5010; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5526 = 3'h4 == state ? valid_0_48 : _GEN_5011; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5527 = 3'h4 == state ? valid_0_49 : _GEN_5012; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5528 = 3'h4 == state ? valid_0_50 : _GEN_5013; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5529 = 3'h4 == state ? valid_0_51 : _GEN_5014; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5530 = 3'h4 == state ? valid_0_52 : _GEN_5015; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5531 = 3'h4 == state ? valid_0_53 : _GEN_5016; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5532 = 3'h4 == state ? valid_0_54 : _GEN_5017; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5533 = 3'h4 == state ? valid_0_55 : _GEN_5018; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5534 = 3'h4 == state ? valid_0_56 : _GEN_5019; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5535 = 3'h4 == state ? valid_0_57 : _GEN_5020; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5536 = 3'h4 == state ? valid_0_58 : _GEN_5021; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5537 = 3'h4 == state ? valid_0_59 : _GEN_5022; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5538 = 3'h4 == state ? valid_0_60 : _GEN_5023; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5539 = 3'h4 == state ? valid_0_61 : _GEN_5024; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5540 = 3'h4 == state ? valid_0_62 : _GEN_5025; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5541 = 3'h4 == state ? valid_0_63 : _GEN_5026; // @[d_cache.scala 81:18 24:26]
  wire [63:0] _GEN_5542 = 3'h4 == state ? ram_1_0 : _GEN_5027; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5543 = 3'h4 == state ? ram_1_1 : _GEN_5028; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5544 = 3'h4 == state ? ram_1_2 : _GEN_5029; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5545 = 3'h4 == state ? ram_1_3 : _GEN_5030; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5546 = 3'h4 == state ? ram_1_4 : _GEN_5031; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5547 = 3'h4 == state ? ram_1_5 : _GEN_5032; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5548 = 3'h4 == state ? ram_1_6 : _GEN_5033; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5549 = 3'h4 == state ? ram_1_7 : _GEN_5034; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5550 = 3'h4 == state ? ram_1_8 : _GEN_5035; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5551 = 3'h4 == state ? ram_1_9 : _GEN_5036; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5552 = 3'h4 == state ? ram_1_10 : _GEN_5037; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5553 = 3'h4 == state ? ram_1_11 : _GEN_5038; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5554 = 3'h4 == state ? ram_1_12 : _GEN_5039; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5555 = 3'h4 == state ? ram_1_13 : _GEN_5040; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5556 = 3'h4 == state ? ram_1_14 : _GEN_5041; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5557 = 3'h4 == state ? ram_1_15 : _GEN_5042; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5558 = 3'h4 == state ? ram_1_16 : _GEN_5043; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5559 = 3'h4 == state ? ram_1_17 : _GEN_5044; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5560 = 3'h4 == state ? ram_1_18 : _GEN_5045; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5561 = 3'h4 == state ? ram_1_19 : _GEN_5046; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5562 = 3'h4 == state ? ram_1_20 : _GEN_5047; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5563 = 3'h4 == state ? ram_1_21 : _GEN_5048; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5564 = 3'h4 == state ? ram_1_22 : _GEN_5049; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5565 = 3'h4 == state ? ram_1_23 : _GEN_5050; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5566 = 3'h4 == state ? ram_1_24 : _GEN_5051; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5567 = 3'h4 == state ? ram_1_25 : _GEN_5052; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5568 = 3'h4 == state ? ram_1_26 : _GEN_5053; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5569 = 3'h4 == state ? ram_1_27 : _GEN_5054; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5570 = 3'h4 == state ? ram_1_28 : _GEN_5055; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5571 = 3'h4 == state ? ram_1_29 : _GEN_5056; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5572 = 3'h4 == state ? ram_1_30 : _GEN_5057; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5573 = 3'h4 == state ? ram_1_31 : _GEN_5058; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5574 = 3'h4 == state ? ram_1_32 : _GEN_5059; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5575 = 3'h4 == state ? ram_1_33 : _GEN_5060; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5576 = 3'h4 == state ? ram_1_34 : _GEN_5061; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5577 = 3'h4 == state ? ram_1_35 : _GEN_5062; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5578 = 3'h4 == state ? ram_1_36 : _GEN_5063; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5579 = 3'h4 == state ? ram_1_37 : _GEN_5064; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5580 = 3'h4 == state ? ram_1_38 : _GEN_5065; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5581 = 3'h4 == state ? ram_1_39 : _GEN_5066; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5582 = 3'h4 == state ? ram_1_40 : _GEN_5067; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5583 = 3'h4 == state ? ram_1_41 : _GEN_5068; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5584 = 3'h4 == state ? ram_1_42 : _GEN_5069; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5585 = 3'h4 == state ? ram_1_43 : _GEN_5070; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5586 = 3'h4 == state ? ram_1_44 : _GEN_5071; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5587 = 3'h4 == state ? ram_1_45 : _GEN_5072; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5588 = 3'h4 == state ? ram_1_46 : _GEN_5073; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5589 = 3'h4 == state ? ram_1_47 : _GEN_5074; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5590 = 3'h4 == state ? ram_1_48 : _GEN_5075; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5591 = 3'h4 == state ? ram_1_49 : _GEN_5076; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5592 = 3'h4 == state ? ram_1_50 : _GEN_5077; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5593 = 3'h4 == state ? ram_1_51 : _GEN_5078; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5594 = 3'h4 == state ? ram_1_52 : _GEN_5079; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5595 = 3'h4 == state ? ram_1_53 : _GEN_5080; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5596 = 3'h4 == state ? ram_1_54 : _GEN_5081; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5597 = 3'h4 == state ? ram_1_55 : _GEN_5082; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5598 = 3'h4 == state ? ram_1_56 : _GEN_5083; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5599 = 3'h4 == state ? ram_1_57 : _GEN_5084; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5600 = 3'h4 == state ? ram_1_58 : _GEN_5085; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5601 = 3'h4 == state ? ram_1_59 : _GEN_5086; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5602 = 3'h4 == state ? ram_1_60 : _GEN_5087; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5603 = 3'h4 == state ? ram_1_61 : _GEN_5088; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5604 = 3'h4 == state ? ram_1_62 : _GEN_5089; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_5605 = 3'h4 == state ? ram_1_63 : _GEN_5090; // @[d_cache.scala 81:18 19:24]
  wire [31:0] _GEN_5606 = 3'h4 == state ? tag_1_0 : _GEN_5091; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5607 = 3'h4 == state ? tag_1_1 : _GEN_5092; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5608 = 3'h4 == state ? tag_1_2 : _GEN_5093; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5609 = 3'h4 == state ? tag_1_3 : _GEN_5094; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5610 = 3'h4 == state ? tag_1_4 : _GEN_5095; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5611 = 3'h4 == state ? tag_1_5 : _GEN_5096; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5612 = 3'h4 == state ? tag_1_6 : _GEN_5097; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5613 = 3'h4 == state ? tag_1_7 : _GEN_5098; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5614 = 3'h4 == state ? tag_1_8 : _GEN_5099; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5615 = 3'h4 == state ? tag_1_9 : _GEN_5100; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5616 = 3'h4 == state ? tag_1_10 : _GEN_5101; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5617 = 3'h4 == state ? tag_1_11 : _GEN_5102; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5618 = 3'h4 == state ? tag_1_12 : _GEN_5103; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5619 = 3'h4 == state ? tag_1_13 : _GEN_5104; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5620 = 3'h4 == state ? tag_1_14 : _GEN_5105; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5621 = 3'h4 == state ? tag_1_15 : _GEN_5106; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5622 = 3'h4 == state ? tag_1_16 : _GEN_5107; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5623 = 3'h4 == state ? tag_1_17 : _GEN_5108; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5624 = 3'h4 == state ? tag_1_18 : _GEN_5109; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5625 = 3'h4 == state ? tag_1_19 : _GEN_5110; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5626 = 3'h4 == state ? tag_1_20 : _GEN_5111; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5627 = 3'h4 == state ? tag_1_21 : _GEN_5112; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5628 = 3'h4 == state ? tag_1_22 : _GEN_5113; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5629 = 3'h4 == state ? tag_1_23 : _GEN_5114; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5630 = 3'h4 == state ? tag_1_24 : _GEN_5115; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5631 = 3'h4 == state ? tag_1_25 : _GEN_5116; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5632 = 3'h4 == state ? tag_1_26 : _GEN_5117; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5633 = 3'h4 == state ? tag_1_27 : _GEN_5118; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5634 = 3'h4 == state ? tag_1_28 : _GEN_5119; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5635 = 3'h4 == state ? tag_1_29 : _GEN_5120; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5636 = 3'h4 == state ? tag_1_30 : _GEN_5121; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5637 = 3'h4 == state ? tag_1_31 : _GEN_5122; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5638 = 3'h4 == state ? tag_1_32 : _GEN_5123; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5639 = 3'h4 == state ? tag_1_33 : _GEN_5124; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5640 = 3'h4 == state ? tag_1_34 : _GEN_5125; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5641 = 3'h4 == state ? tag_1_35 : _GEN_5126; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5642 = 3'h4 == state ? tag_1_36 : _GEN_5127; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5643 = 3'h4 == state ? tag_1_37 : _GEN_5128; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5644 = 3'h4 == state ? tag_1_38 : _GEN_5129; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5645 = 3'h4 == state ? tag_1_39 : _GEN_5130; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5646 = 3'h4 == state ? tag_1_40 : _GEN_5131; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5647 = 3'h4 == state ? tag_1_41 : _GEN_5132; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5648 = 3'h4 == state ? tag_1_42 : _GEN_5133; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5649 = 3'h4 == state ? tag_1_43 : _GEN_5134; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5650 = 3'h4 == state ? tag_1_44 : _GEN_5135; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5651 = 3'h4 == state ? tag_1_45 : _GEN_5136; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5652 = 3'h4 == state ? tag_1_46 : _GEN_5137; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5653 = 3'h4 == state ? tag_1_47 : _GEN_5138; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5654 = 3'h4 == state ? tag_1_48 : _GEN_5139; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5655 = 3'h4 == state ? tag_1_49 : _GEN_5140; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5656 = 3'h4 == state ? tag_1_50 : _GEN_5141; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5657 = 3'h4 == state ? tag_1_51 : _GEN_5142; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5658 = 3'h4 == state ? tag_1_52 : _GEN_5143; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5659 = 3'h4 == state ? tag_1_53 : _GEN_5144; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5660 = 3'h4 == state ? tag_1_54 : _GEN_5145; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5661 = 3'h4 == state ? tag_1_55 : _GEN_5146; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5662 = 3'h4 == state ? tag_1_56 : _GEN_5147; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5663 = 3'h4 == state ? tag_1_57 : _GEN_5148; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5664 = 3'h4 == state ? tag_1_58 : _GEN_5149; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5665 = 3'h4 == state ? tag_1_59 : _GEN_5150; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5666 = 3'h4 == state ? tag_1_60 : _GEN_5151; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5667 = 3'h4 == state ? tag_1_61 : _GEN_5152; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5668 = 3'h4 == state ? tag_1_62 : _GEN_5153; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_5669 = 3'h4 == state ? tag_1_63 : _GEN_5154; // @[d_cache.scala 81:18 23:24]
  wire  _GEN_5670 = 3'h4 == state ? valid_1_0 : _GEN_5155; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5671 = 3'h4 == state ? valid_1_1 : _GEN_5156; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5672 = 3'h4 == state ? valid_1_2 : _GEN_5157; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5673 = 3'h4 == state ? valid_1_3 : _GEN_5158; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5674 = 3'h4 == state ? valid_1_4 : _GEN_5159; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5675 = 3'h4 == state ? valid_1_5 : _GEN_5160; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5676 = 3'h4 == state ? valid_1_6 : _GEN_5161; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5677 = 3'h4 == state ? valid_1_7 : _GEN_5162; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5678 = 3'h4 == state ? valid_1_8 : _GEN_5163; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5679 = 3'h4 == state ? valid_1_9 : _GEN_5164; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5680 = 3'h4 == state ? valid_1_10 : _GEN_5165; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5681 = 3'h4 == state ? valid_1_11 : _GEN_5166; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5682 = 3'h4 == state ? valid_1_12 : _GEN_5167; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5683 = 3'h4 == state ? valid_1_13 : _GEN_5168; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5684 = 3'h4 == state ? valid_1_14 : _GEN_5169; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5685 = 3'h4 == state ? valid_1_15 : _GEN_5170; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5686 = 3'h4 == state ? valid_1_16 : _GEN_5171; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5687 = 3'h4 == state ? valid_1_17 : _GEN_5172; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5688 = 3'h4 == state ? valid_1_18 : _GEN_5173; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5689 = 3'h4 == state ? valid_1_19 : _GEN_5174; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5690 = 3'h4 == state ? valid_1_20 : _GEN_5175; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5691 = 3'h4 == state ? valid_1_21 : _GEN_5176; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5692 = 3'h4 == state ? valid_1_22 : _GEN_5177; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5693 = 3'h4 == state ? valid_1_23 : _GEN_5178; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5694 = 3'h4 == state ? valid_1_24 : _GEN_5179; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5695 = 3'h4 == state ? valid_1_25 : _GEN_5180; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5696 = 3'h4 == state ? valid_1_26 : _GEN_5181; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5697 = 3'h4 == state ? valid_1_27 : _GEN_5182; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5698 = 3'h4 == state ? valid_1_28 : _GEN_5183; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5699 = 3'h4 == state ? valid_1_29 : _GEN_5184; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5700 = 3'h4 == state ? valid_1_30 : _GEN_5185; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5701 = 3'h4 == state ? valid_1_31 : _GEN_5186; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5702 = 3'h4 == state ? valid_1_32 : _GEN_5187; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5703 = 3'h4 == state ? valid_1_33 : _GEN_5188; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5704 = 3'h4 == state ? valid_1_34 : _GEN_5189; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5705 = 3'h4 == state ? valid_1_35 : _GEN_5190; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5706 = 3'h4 == state ? valid_1_36 : _GEN_5191; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5707 = 3'h4 == state ? valid_1_37 : _GEN_5192; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5708 = 3'h4 == state ? valid_1_38 : _GEN_5193; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5709 = 3'h4 == state ? valid_1_39 : _GEN_5194; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5710 = 3'h4 == state ? valid_1_40 : _GEN_5195; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5711 = 3'h4 == state ? valid_1_41 : _GEN_5196; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5712 = 3'h4 == state ? valid_1_42 : _GEN_5197; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5713 = 3'h4 == state ? valid_1_43 : _GEN_5198; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5714 = 3'h4 == state ? valid_1_44 : _GEN_5199; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5715 = 3'h4 == state ? valid_1_45 : _GEN_5200; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5716 = 3'h4 == state ? valid_1_46 : _GEN_5201; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5717 = 3'h4 == state ? valid_1_47 : _GEN_5202; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5718 = 3'h4 == state ? valid_1_48 : _GEN_5203; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5719 = 3'h4 == state ? valid_1_49 : _GEN_5204; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5720 = 3'h4 == state ? valid_1_50 : _GEN_5205; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5721 = 3'h4 == state ? valid_1_51 : _GEN_5206; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5722 = 3'h4 == state ? valid_1_52 : _GEN_5207; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5723 = 3'h4 == state ? valid_1_53 : _GEN_5208; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5724 = 3'h4 == state ? valid_1_54 : _GEN_5209; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5725 = 3'h4 == state ? valid_1_55 : _GEN_5210; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5726 = 3'h4 == state ? valid_1_56 : _GEN_5211; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5727 = 3'h4 == state ? valid_1_57 : _GEN_5212; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5728 = 3'h4 == state ? valid_1_58 : _GEN_5213; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5729 = 3'h4 == state ? valid_1_59 : _GEN_5214; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5730 = 3'h4 == state ? valid_1_60 : _GEN_5215; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5731 = 3'h4 == state ? valid_1_61 : _GEN_5216; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5732 = 3'h4 == state ? valid_1_62 : _GEN_5217; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_5733 = 3'h4 == state ? valid_1_63 : _GEN_5218; // @[d_cache.scala 81:18 25:26]
  wire [63:0] _GEN_5734 = 3'h4 == state ? write_back_data : _GEN_5219; // @[d_cache.scala 81:18 31:34]
  wire [40:0] _GEN_5735 = 3'h4 == state ? {{9'd0}, write_back_addr} : _GEN_5220; // @[d_cache.scala 81:18 32:34]
  wire  _GEN_5736 = 3'h4 == state ? dirty_0_0 : _GEN_5221; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5737 = 3'h4 == state ? dirty_0_1 : _GEN_5222; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5738 = 3'h4 == state ? dirty_0_2 : _GEN_5223; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5739 = 3'h4 == state ? dirty_0_3 : _GEN_5224; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5740 = 3'h4 == state ? dirty_0_4 : _GEN_5225; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5741 = 3'h4 == state ? dirty_0_5 : _GEN_5226; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5742 = 3'h4 == state ? dirty_0_6 : _GEN_5227; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5743 = 3'h4 == state ? dirty_0_7 : _GEN_5228; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5744 = 3'h4 == state ? dirty_0_8 : _GEN_5229; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5745 = 3'h4 == state ? dirty_0_9 : _GEN_5230; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5746 = 3'h4 == state ? dirty_0_10 : _GEN_5231; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5747 = 3'h4 == state ? dirty_0_11 : _GEN_5232; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5748 = 3'h4 == state ? dirty_0_12 : _GEN_5233; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5749 = 3'h4 == state ? dirty_0_13 : _GEN_5234; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5750 = 3'h4 == state ? dirty_0_14 : _GEN_5235; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5751 = 3'h4 == state ? dirty_0_15 : _GEN_5236; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5752 = 3'h4 == state ? dirty_0_16 : _GEN_5237; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5753 = 3'h4 == state ? dirty_0_17 : _GEN_5238; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5754 = 3'h4 == state ? dirty_0_18 : _GEN_5239; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5755 = 3'h4 == state ? dirty_0_19 : _GEN_5240; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5756 = 3'h4 == state ? dirty_0_20 : _GEN_5241; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5757 = 3'h4 == state ? dirty_0_21 : _GEN_5242; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5758 = 3'h4 == state ? dirty_0_22 : _GEN_5243; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5759 = 3'h4 == state ? dirty_0_23 : _GEN_5244; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5760 = 3'h4 == state ? dirty_0_24 : _GEN_5245; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5761 = 3'h4 == state ? dirty_0_25 : _GEN_5246; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5762 = 3'h4 == state ? dirty_0_26 : _GEN_5247; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5763 = 3'h4 == state ? dirty_0_27 : _GEN_5248; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5764 = 3'h4 == state ? dirty_0_28 : _GEN_5249; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5765 = 3'h4 == state ? dirty_0_29 : _GEN_5250; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5766 = 3'h4 == state ? dirty_0_30 : _GEN_5251; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5767 = 3'h4 == state ? dirty_0_31 : _GEN_5252; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5768 = 3'h4 == state ? dirty_0_32 : _GEN_5253; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5769 = 3'h4 == state ? dirty_0_33 : _GEN_5254; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5770 = 3'h4 == state ? dirty_0_34 : _GEN_5255; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5771 = 3'h4 == state ? dirty_0_35 : _GEN_5256; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5772 = 3'h4 == state ? dirty_0_36 : _GEN_5257; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5773 = 3'h4 == state ? dirty_0_37 : _GEN_5258; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5774 = 3'h4 == state ? dirty_0_38 : _GEN_5259; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5775 = 3'h4 == state ? dirty_0_39 : _GEN_5260; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5776 = 3'h4 == state ? dirty_0_40 : _GEN_5261; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5777 = 3'h4 == state ? dirty_0_41 : _GEN_5262; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5778 = 3'h4 == state ? dirty_0_42 : _GEN_5263; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5779 = 3'h4 == state ? dirty_0_43 : _GEN_5264; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5780 = 3'h4 == state ? dirty_0_44 : _GEN_5265; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5781 = 3'h4 == state ? dirty_0_45 : _GEN_5266; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5782 = 3'h4 == state ? dirty_0_46 : _GEN_5267; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5783 = 3'h4 == state ? dirty_0_47 : _GEN_5268; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5784 = 3'h4 == state ? dirty_0_48 : _GEN_5269; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5785 = 3'h4 == state ? dirty_0_49 : _GEN_5270; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5786 = 3'h4 == state ? dirty_0_50 : _GEN_5271; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5787 = 3'h4 == state ? dirty_0_51 : _GEN_5272; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5788 = 3'h4 == state ? dirty_0_52 : _GEN_5273; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5789 = 3'h4 == state ? dirty_0_53 : _GEN_5274; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5790 = 3'h4 == state ? dirty_0_54 : _GEN_5275; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5791 = 3'h4 == state ? dirty_0_55 : _GEN_5276; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5792 = 3'h4 == state ? dirty_0_56 : _GEN_5277; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5793 = 3'h4 == state ? dirty_0_57 : _GEN_5278; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5794 = 3'h4 == state ? dirty_0_58 : _GEN_5279; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5795 = 3'h4 == state ? dirty_0_59 : _GEN_5280; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5796 = 3'h4 == state ? dirty_0_60 : _GEN_5281; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5797 = 3'h4 == state ? dirty_0_61 : _GEN_5282; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5798 = 3'h4 == state ? dirty_0_62 : _GEN_5283; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5799 = 3'h4 == state ? dirty_0_63 : _GEN_5284; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_5800 = 3'h4 == state ? dirty_1_0 : _GEN_5285; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5801 = 3'h4 == state ? dirty_1_1 : _GEN_5286; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5802 = 3'h4 == state ? dirty_1_2 : _GEN_5287; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5803 = 3'h4 == state ? dirty_1_3 : _GEN_5288; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5804 = 3'h4 == state ? dirty_1_4 : _GEN_5289; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5805 = 3'h4 == state ? dirty_1_5 : _GEN_5290; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5806 = 3'h4 == state ? dirty_1_6 : _GEN_5291; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5807 = 3'h4 == state ? dirty_1_7 : _GEN_5292; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5808 = 3'h4 == state ? dirty_1_8 : _GEN_5293; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5809 = 3'h4 == state ? dirty_1_9 : _GEN_5294; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5810 = 3'h4 == state ? dirty_1_10 : _GEN_5295; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5811 = 3'h4 == state ? dirty_1_11 : _GEN_5296; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5812 = 3'h4 == state ? dirty_1_12 : _GEN_5297; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5813 = 3'h4 == state ? dirty_1_13 : _GEN_5298; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5814 = 3'h4 == state ? dirty_1_14 : _GEN_5299; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5815 = 3'h4 == state ? dirty_1_15 : _GEN_5300; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5816 = 3'h4 == state ? dirty_1_16 : _GEN_5301; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5817 = 3'h4 == state ? dirty_1_17 : _GEN_5302; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5818 = 3'h4 == state ? dirty_1_18 : _GEN_5303; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5819 = 3'h4 == state ? dirty_1_19 : _GEN_5304; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5820 = 3'h4 == state ? dirty_1_20 : _GEN_5305; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5821 = 3'h4 == state ? dirty_1_21 : _GEN_5306; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5822 = 3'h4 == state ? dirty_1_22 : _GEN_5307; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5823 = 3'h4 == state ? dirty_1_23 : _GEN_5308; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5824 = 3'h4 == state ? dirty_1_24 : _GEN_5309; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5825 = 3'h4 == state ? dirty_1_25 : _GEN_5310; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5826 = 3'h4 == state ? dirty_1_26 : _GEN_5311; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5827 = 3'h4 == state ? dirty_1_27 : _GEN_5312; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5828 = 3'h4 == state ? dirty_1_28 : _GEN_5313; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5829 = 3'h4 == state ? dirty_1_29 : _GEN_5314; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5830 = 3'h4 == state ? dirty_1_30 : _GEN_5315; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5831 = 3'h4 == state ? dirty_1_31 : _GEN_5316; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5832 = 3'h4 == state ? dirty_1_32 : _GEN_5317; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5833 = 3'h4 == state ? dirty_1_33 : _GEN_5318; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5834 = 3'h4 == state ? dirty_1_34 : _GEN_5319; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5835 = 3'h4 == state ? dirty_1_35 : _GEN_5320; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5836 = 3'h4 == state ? dirty_1_36 : _GEN_5321; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5837 = 3'h4 == state ? dirty_1_37 : _GEN_5322; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5838 = 3'h4 == state ? dirty_1_38 : _GEN_5323; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5839 = 3'h4 == state ? dirty_1_39 : _GEN_5324; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5840 = 3'h4 == state ? dirty_1_40 : _GEN_5325; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5841 = 3'h4 == state ? dirty_1_41 : _GEN_5326; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5842 = 3'h4 == state ? dirty_1_42 : _GEN_5327; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5843 = 3'h4 == state ? dirty_1_43 : _GEN_5328; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5844 = 3'h4 == state ? dirty_1_44 : _GEN_5329; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5845 = 3'h4 == state ? dirty_1_45 : _GEN_5330; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5846 = 3'h4 == state ? dirty_1_46 : _GEN_5331; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5847 = 3'h4 == state ? dirty_1_47 : _GEN_5332; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5848 = 3'h4 == state ? dirty_1_48 : _GEN_5333; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5849 = 3'h4 == state ? dirty_1_49 : _GEN_5334; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5850 = 3'h4 == state ? dirty_1_50 : _GEN_5335; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5851 = 3'h4 == state ? dirty_1_51 : _GEN_5336; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5852 = 3'h4 == state ? dirty_1_52 : _GEN_5337; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5853 = 3'h4 == state ? dirty_1_53 : _GEN_5338; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5854 = 3'h4 == state ? dirty_1_54 : _GEN_5339; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5855 = 3'h4 == state ? dirty_1_55 : _GEN_5340; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5856 = 3'h4 == state ? dirty_1_56 : _GEN_5341; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5857 = 3'h4 == state ? dirty_1_57 : _GEN_5342; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5858 = 3'h4 == state ? dirty_1_58 : _GEN_5343; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5859 = 3'h4 == state ? dirty_1_59 : _GEN_5344; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5860 = 3'h4 == state ? dirty_1_60 : _GEN_5345; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5861 = 3'h4 == state ? dirty_1_61 : _GEN_5346; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5862 = 3'h4 == state ? dirty_1_62 : _GEN_5347; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_5863 = 3'h4 == state ? dirty_1_63 : _GEN_5348; // @[d_cache.scala 81:18 27:26]
  wire [2:0] _GEN_5864 = 3'h3 == state ? _GEN_1485 : _GEN_5349; // @[d_cache.scala 81:18]
  wire [63:0] _GEN_5865 = 3'h3 == state ? _GEN_1486 : receive_data; // @[d_cache.scala 81:18 36:31]
  wire [63:0] _GEN_5866 = 3'h3 == state ? ram_0_0 : _GEN_5350; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5867 = 3'h3 == state ? ram_0_1 : _GEN_5351; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5868 = 3'h3 == state ? ram_0_2 : _GEN_5352; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5869 = 3'h3 == state ? ram_0_3 : _GEN_5353; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5870 = 3'h3 == state ? ram_0_4 : _GEN_5354; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5871 = 3'h3 == state ? ram_0_5 : _GEN_5355; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5872 = 3'h3 == state ? ram_0_6 : _GEN_5356; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5873 = 3'h3 == state ? ram_0_7 : _GEN_5357; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5874 = 3'h3 == state ? ram_0_8 : _GEN_5358; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5875 = 3'h3 == state ? ram_0_9 : _GEN_5359; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5876 = 3'h3 == state ? ram_0_10 : _GEN_5360; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5877 = 3'h3 == state ? ram_0_11 : _GEN_5361; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5878 = 3'h3 == state ? ram_0_12 : _GEN_5362; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5879 = 3'h3 == state ? ram_0_13 : _GEN_5363; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5880 = 3'h3 == state ? ram_0_14 : _GEN_5364; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5881 = 3'h3 == state ? ram_0_15 : _GEN_5365; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5882 = 3'h3 == state ? ram_0_16 : _GEN_5366; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5883 = 3'h3 == state ? ram_0_17 : _GEN_5367; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5884 = 3'h3 == state ? ram_0_18 : _GEN_5368; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5885 = 3'h3 == state ? ram_0_19 : _GEN_5369; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5886 = 3'h3 == state ? ram_0_20 : _GEN_5370; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5887 = 3'h3 == state ? ram_0_21 : _GEN_5371; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5888 = 3'h3 == state ? ram_0_22 : _GEN_5372; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5889 = 3'h3 == state ? ram_0_23 : _GEN_5373; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5890 = 3'h3 == state ? ram_0_24 : _GEN_5374; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5891 = 3'h3 == state ? ram_0_25 : _GEN_5375; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5892 = 3'h3 == state ? ram_0_26 : _GEN_5376; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5893 = 3'h3 == state ? ram_0_27 : _GEN_5377; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5894 = 3'h3 == state ? ram_0_28 : _GEN_5378; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5895 = 3'h3 == state ? ram_0_29 : _GEN_5379; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5896 = 3'h3 == state ? ram_0_30 : _GEN_5380; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5897 = 3'h3 == state ? ram_0_31 : _GEN_5381; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5898 = 3'h3 == state ? ram_0_32 : _GEN_5382; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5899 = 3'h3 == state ? ram_0_33 : _GEN_5383; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5900 = 3'h3 == state ? ram_0_34 : _GEN_5384; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5901 = 3'h3 == state ? ram_0_35 : _GEN_5385; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5902 = 3'h3 == state ? ram_0_36 : _GEN_5386; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5903 = 3'h3 == state ? ram_0_37 : _GEN_5387; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5904 = 3'h3 == state ? ram_0_38 : _GEN_5388; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5905 = 3'h3 == state ? ram_0_39 : _GEN_5389; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5906 = 3'h3 == state ? ram_0_40 : _GEN_5390; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5907 = 3'h3 == state ? ram_0_41 : _GEN_5391; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5908 = 3'h3 == state ? ram_0_42 : _GEN_5392; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5909 = 3'h3 == state ? ram_0_43 : _GEN_5393; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5910 = 3'h3 == state ? ram_0_44 : _GEN_5394; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5911 = 3'h3 == state ? ram_0_45 : _GEN_5395; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5912 = 3'h3 == state ? ram_0_46 : _GEN_5396; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5913 = 3'h3 == state ? ram_0_47 : _GEN_5397; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5914 = 3'h3 == state ? ram_0_48 : _GEN_5398; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5915 = 3'h3 == state ? ram_0_49 : _GEN_5399; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5916 = 3'h3 == state ? ram_0_50 : _GEN_5400; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5917 = 3'h3 == state ? ram_0_51 : _GEN_5401; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5918 = 3'h3 == state ? ram_0_52 : _GEN_5402; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5919 = 3'h3 == state ? ram_0_53 : _GEN_5403; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5920 = 3'h3 == state ? ram_0_54 : _GEN_5404; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5921 = 3'h3 == state ? ram_0_55 : _GEN_5405; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5922 = 3'h3 == state ? ram_0_56 : _GEN_5406; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5923 = 3'h3 == state ? ram_0_57 : _GEN_5407; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5924 = 3'h3 == state ? ram_0_58 : _GEN_5408; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5925 = 3'h3 == state ? ram_0_59 : _GEN_5409; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5926 = 3'h3 == state ? ram_0_60 : _GEN_5410; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5927 = 3'h3 == state ? ram_0_61 : _GEN_5411; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5928 = 3'h3 == state ? ram_0_62 : _GEN_5412; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_5929 = 3'h3 == state ? ram_0_63 : _GEN_5413; // @[d_cache.scala 81:18 18:24]
  wire [31:0] _GEN_5930 = 3'h3 == state ? tag_0_0 : _GEN_5414; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5931 = 3'h3 == state ? tag_0_1 : _GEN_5415; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5932 = 3'h3 == state ? tag_0_2 : _GEN_5416; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5933 = 3'h3 == state ? tag_0_3 : _GEN_5417; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5934 = 3'h3 == state ? tag_0_4 : _GEN_5418; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5935 = 3'h3 == state ? tag_0_5 : _GEN_5419; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5936 = 3'h3 == state ? tag_0_6 : _GEN_5420; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5937 = 3'h3 == state ? tag_0_7 : _GEN_5421; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5938 = 3'h3 == state ? tag_0_8 : _GEN_5422; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5939 = 3'h3 == state ? tag_0_9 : _GEN_5423; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5940 = 3'h3 == state ? tag_0_10 : _GEN_5424; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5941 = 3'h3 == state ? tag_0_11 : _GEN_5425; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5942 = 3'h3 == state ? tag_0_12 : _GEN_5426; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5943 = 3'h3 == state ? tag_0_13 : _GEN_5427; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5944 = 3'h3 == state ? tag_0_14 : _GEN_5428; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5945 = 3'h3 == state ? tag_0_15 : _GEN_5429; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5946 = 3'h3 == state ? tag_0_16 : _GEN_5430; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5947 = 3'h3 == state ? tag_0_17 : _GEN_5431; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5948 = 3'h3 == state ? tag_0_18 : _GEN_5432; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5949 = 3'h3 == state ? tag_0_19 : _GEN_5433; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5950 = 3'h3 == state ? tag_0_20 : _GEN_5434; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5951 = 3'h3 == state ? tag_0_21 : _GEN_5435; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5952 = 3'h3 == state ? tag_0_22 : _GEN_5436; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5953 = 3'h3 == state ? tag_0_23 : _GEN_5437; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5954 = 3'h3 == state ? tag_0_24 : _GEN_5438; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5955 = 3'h3 == state ? tag_0_25 : _GEN_5439; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5956 = 3'h3 == state ? tag_0_26 : _GEN_5440; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5957 = 3'h3 == state ? tag_0_27 : _GEN_5441; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5958 = 3'h3 == state ? tag_0_28 : _GEN_5442; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5959 = 3'h3 == state ? tag_0_29 : _GEN_5443; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5960 = 3'h3 == state ? tag_0_30 : _GEN_5444; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5961 = 3'h3 == state ? tag_0_31 : _GEN_5445; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5962 = 3'h3 == state ? tag_0_32 : _GEN_5446; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5963 = 3'h3 == state ? tag_0_33 : _GEN_5447; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5964 = 3'h3 == state ? tag_0_34 : _GEN_5448; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5965 = 3'h3 == state ? tag_0_35 : _GEN_5449; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5966 = 3'h3 == state ? tag_0_36 : _GEN_5450; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5967 = 3'h3 == state ? tag_0_37 : _GEN_5451; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5968 = 3'h3 == state ? tag_0_38 : _GEN_5452; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5969 = 3'h3 == state ? tag_0_39 : _GEN_5453; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5970 = 3'h3 == state ? tag_0_40 : _GEN_5454; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5971 = 3'h3 == state ? tag_0_41 : _GEN_5455; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5972 = 3'h3 == state ? tag_0_42 : _GEN_5456; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5973 = 3'h3 == state ? tag_0_43 : _GEN_5457; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5974 = 3'h3 == state ? tag_0_44 : _GEN_5458; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5975 = 3'h3 == state ? tag_0_45 : _GEN_5459; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5976 = 3'h3 == state ? tag_0_46 : _GEN_5460; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5977 = 3'h3 == state ? tag_0_47 : _GEN_5461; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5978 = 3'h3 == state ? tag_0_48 : _GEN_5462; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5979 = 3'h3 == state ? tag_0_49 : _GEN_5463; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5980 = 3'h3 == state ? tag_0_50 : _GEN_5464; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5981 = 3'h3 == state ? tag_0_51 : _GEN_5465; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5982 = 3'h3 == state ? tag_0_52 : _GEN_5466; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5983 = 3'h3 == state ? tag_0_53 : _GEN_5467; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5984 = 3'h3 == state ? tag_0_54 : _GEN_5468; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5985 = 3'h3 == state ? tag_0_55 : _GEN_5469; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5986 = 3'h3 == state ? tag_0_56 : _GEN_5470; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5987 = 3'h3 == state ? tag_0_57 : _GEN_5471; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5988 = 3'h3 == state ? tag_0_58 : _GEN_5472; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5989 = 3'h3 == state ? tag_0_59 : _GEN_5473; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5990 = 3'h3 == state ? tag_0_60 : _GEN_5474; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5991 = 3'h3 == state ? tag_0_61 : _GEN_5475; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5992 = 3'h3 == state ? tag_0_62 : _GEN_5476; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_5993 = 3'h3 == state ? tag_0_63 : _GEN_5477; // @[d_cache.scala 81:18 22:24]
  wire  _GEN_5994 = 3'h3 == state ? valid_0_0 : _GEN_5478; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5995 = 3'h3 == state ? valid_0_1 : _GEN_5479; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5996 = 3'h3 == state ? valid_0_2 : _GEN_5480; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5997 = 3'h3 == state ? valid_0_3 : _GEN_5481; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5998 = 3'h3 == state ? valid_0_4 : _GEN_5482; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_5999 = 3'h3 == state ? valid_0_5 : _GEN_5483; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6000 = 3'h3 == state ? valid_0_6 : _GEN_5484; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6001 = 3'h3 == state ? valid_0_7 : _GEN_5485; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6002 = 3'h3 == state ? valid_0_8 : _GEN_5486; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6003 = 3'h3 == state ? valid_0_9 : _GEN_5487; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6004 = 3'h3 == state ? valid_0_10 : _GEN_5488; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6005 = 3'h3 == state ? valid_0_11 : _GEN_5489; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6006 = 3'h3 == state ? valid_0_12 : _GEN_5490; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6007 = 3'h3 == state ? valid_0_13 : _GEN_5491; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6008 = 3'h3 == state ? valid_0_14 : _GEN_5492; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6009 = 3'h3 == state ? valid_0_15 : _GEN_5493; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6010 = 3'h3 == state ? valid_0_16 : _GEN_5494; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6011 = 3'h3 == state ? valid_0_17 : _GEN_5495; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6012 = 3'h3 == state ? valid_0_18 : _GEN_5496; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6013 = 3'h3 == state ? valid_0_19 : _GEN_5497; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6014 = 3'h3 == state ? valid_0_20 : _GEN_5498; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6015 = 3'h3 == state ? valid_0_21 : _GEN_5499; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6016 = 3'h3 == state ? valid_0_22 : _GEN_5500; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6017 = 3'h3 == state ? valid_0_23 : _GEN_5501; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6018 = 3'h3 == state ? valid_0_24 : _GEN_5502; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6019 = 3'h3 == state ? valid_0_25 : _GEN_5503; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6020 = 3'h3 == state ? valid_0_26 : _GEN_5504; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6021 = 3'h3 == state ? valid_0_27 : _GEN_5505; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6022 = 3'h3 == state ? valid_0_28 : _GEN_5506; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6023 = 3'h3 == state ? valid_0_29 : _GEN_5507; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6024 = 3'h3 == state ? valid_0_30 : _GEN_5508; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6025 = 3'h3 == state ? valid_0_31 : _GEN_5509; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6026 = 3'h3 == state ? valid_0_32 : _GEN_5510; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6027 = 3'h3 == state ? valid_0_33 : _GEN_5511; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6028 = 3'h3 == state ? valid_0_34 : _GEN_5512; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6029 = 3'h3 == state ? valid_0_35 : _GEN_5513; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6030 = 3'h3 == state ? valid_0_36 : _GEN_5514; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6031 = 3'h3 == state ? valid_0_37 : _GEN_5515; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6032 = 3'h3 == state ? valid_0_38 : _GEN_5516; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6033 = 3'h3 == state ? valid_0_39 : _GEN_5517; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6034 = 3'h3 == state ? valid_0_40 : _GEN_5518; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6035 = 3'h3 == state ? valid_0_41 : _GEN_5519; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6036 = 3'h3 == state ? valid_0_42 : _GEN_5520; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6037 = 3'h3 == state ? valid_0_43 : _GEN_5521; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6038 = 3'h3 == state ? valid_0_44 : _GEN_5522; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6039 = 3'h3 == state ? valid_0_45 : _GEN_5523; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6040 = 3'h3 == state ? valid_0_46 : _GEN_5524; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6041 = 3'h3 == state ? valid_0_47 : _GEN_5525; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6042 = 3'h3 == state ? valid_0_48 : _GEN_5526; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6043 = 3'h3 == state ? valid_0_49 : _GEN_5527; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6044 = 3'h3 == state ? valid_0_50 : _GEN_5528; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6045 = 3'h3 == state ? valid_0_51 : _GEN_5529; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6046 = 3'h3 == state ? valid_0_52 : _GEN_5530; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6047 = 3'h3 == state ? valid_0_53 : _GEN_5531; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6048 = 3'h3 == state ? valid_0_54 : _GEN_5532; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6049 = 3'h3 == state ? valid_0_55 : _GEN_5533; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6050 = 3'h3 == state ? valid_0_56 : _GEN_5534; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6051 = 3'h3 == state ? valid_0_57 : _GEN_5535; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6052 = 3'h3 == state ? valid_0_58 : _GEN_5536; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6053 = 3'h3 == state ? valid_0_59 : _GEN_5537; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6054 = 3'h3 == state ? valid_0_60 : _GEN_5538; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6055 = 3'h3 == state ? valid_0_61 : _GEN_5539; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6056 = 3'h3 == state ? valid_0_62 : _GEN_5540; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_6057 = 3'h3 == state ? valid_0_63 : _GEN_5541; // @[d_cache.scala 81:18 24:26]
  wire [63:0] _GEN_6058 = 3'h3 == state ? ram_1_0 : _GEN_5542; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6059 = 3'h3 == state ? ram_1_1 : _GEN_5543; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6060 = 3'h3 == state ? ram_1_2 : _GEN_5544; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6061 = 3'h3 == state ? ram_1_3 : _GEN_5545; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6062 = 3'h3 == state ? ram_1_4 : _GEN_5546; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6063 = 3'h3 == state ? ram_1_5 : _GEN_5547; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6064 = 3'h3 == state ? ram_1_6 : _GEN_5548; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6065 = 3'h3 == state ? ram_1_7 : _GEN_5549; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6066 = 3'h3 == state ? ram_1_8 : _GEN_5550; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6067 = 3'h3 == state ? ram_1_9 : _GEN_5551; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6068 = 3'h3 == state ? ram_1_10 : _GEN_5552; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6069 = 3'h3 == state ? ram_1_11 : _GEN_5553; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6070 = 3'h3 == state ? ram_1_12 : _GEN_5554; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6071 = 3'h3 == state ? ram_1_13 : _GEN_5555; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6072 = 3'h3 == state ? ram_1_14 : _GEN_5556; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6073 = 3'h3 == state ? ram_1_15 : _GEN_5557; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6074 = 3'h3 == state ? ram_1_16 : _GEN_5558; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6075 = 3'h3 == state ? ram_1_17 : _GEN_5559; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6076 = 3'h3 == state ? ram_1_18 : _GEN_5560; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6077 = 3'h3 == state ? ram_1_19 : _GEN_5561; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6078 = 3'h3 == state ? ram_1_20 : _GEN_5562; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6079 = 3'h3 == state ? ram_1_21 : _GEN_5563; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6080 = 3'h3 == state ? ram_1_22 : _GEN_5564; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6081 = 3'h3 == state ? ram_1_23 : _GEN_5565; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6082 = 3'h3 == state ? ram_1_24 : _GEN_5566; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6083 = 3'h3 == state ? ram_1_25 : _GEN_5567; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6084 = 3'h3 == state ? ram_1_26 : _GEN_5568; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6085 = 3'h3 == state ? ram_1_27 : _GEN_5569; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6086 = 3'h3 == state ? ram_1_28 : _GEN_5570; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6087 = 3'h3 == state ? ram_1_29 : _GEN_5571; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6088 = 3'h3 == state ? ram_1_30 : _GEN_5572; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6089 = 3'h3 == state ? ram_1_31 : _GEN_5573; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6090 = 3'h3 == state ? ram_1_32 : _GEN_5574; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6091 = 3'h3 == state ? ram_1_33 : _GEN_5575; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6092 = 3'h3 == state ? ram_1_34 : _GEN_5576; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6093 = 3'h3 == state ? ram_1_35 : _GEN_5577; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6094 = 3'h3 == state ? ram_1_36 : _GEN_5578; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6095 = 3'h3 == state ? ram_1_37 : _GEN_5579; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6096 = 3'h3 == state ? ram_1_38 : _GEN_5580; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6097 = 3'h3 == state ? ram_1_39 : _GEN_5581; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6098 = 3'h3 == state ? ram_1_40 : _GEN_5582; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6099 = 3'h3 == state ? ram_1_41 : _GEN_5583; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6100 = 3'h3 == state ? ram_1_42 : _GEN_5584; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6101 = 3'h3 == state ? ram_1_43 : _GEN_5585; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6102 = 3'h3 == state ? ram_1_44 : _GEN_5586; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6103 = 3'h3 == state ? ram_1_45 : _GEN_5587; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6104 = 3'h3 == state ? ram_1_46 : _GEN_5588; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6105 = 3'h3 == state ? ram_1_47 : _GEN_5589; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6106 = 3'h3 == state ? ram_1_48 : _GEN_5590; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6107 = 3'h3 == state ? ram_1_49 : _GEN_5591; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6108 = 3'h3 == state ? ram_1_50 : _GEN_5592; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6109 = 3'h3 == state ? ram_1_51 : _GEN_5593; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6110 = 3'h3 == state ? ram_1_52 : _GEN_5594; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6111 = 3'h3 == state ? ram_1_53 : _GEN_5595; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6112 = 3'h3 == state ? ram_1_54 : _GEN_5596; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6113 = 3'h3 == state ? ram_1_55 : _GEN_5597; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6114 = 3'h3 == state ? ram_1_56 : _GEN_5598; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6115 = 3'h3 == state ? ram_1_57 : _GEN_5599; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6116 = 3'h3 == state ? ram_1_58 : _GEN_5600; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6117 = 3'h3 == state ? ram_1_59 : _GEN_5601; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6118 = 3'h3 == state ? ram_1_60 : _GEN_5602; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6119 = 3'h3 == state ? ram_1_61 : _GEN_5603; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6120 = 3'h3 == state ? ram_1_62 : _GEN_5604; // @[d_cache.scala 81:18 19:24]
  wire [63:0] _GEN_6121 = 3'h3 == state ? ram_1_63 : _GEN_5605; // @[d_cache.scala 81:18 19:24]
  wire [31:0] _GEN_6122 = 3'h3 == state ? tag_1_0 : _GEN_5606; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6123 = 3'h3 == state ? tag_1_1 : _GEN_5607; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6124 = 3'h3 == state ? tag_1_2 : _GEN_5608; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6125 = 3'h3 == state ? tag_1_3 : _GEN_5609; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6126 = 3'h3 == state ? tag_1_4 : _GEN_5610; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6127 = 3'h3 == state ? tag_1_5 : _GEN_5611; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6128 = 3'h3 == state ? tag_1_6 : _GEN_5612; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6129 = 3'h3 == state ? tag_1_7 : _GEN_5613; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6130 = 3'h3 == state ? tag_1_8 : _GEN_5614; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6131 = 3'h3 == state ? tag_1_9 : _GEN_5615; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6132 = 3'h3 == state ? tag_1_10 : _GEN_5616; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6133 = 3'h3 == state ? tag_1_11 : _GEN_5617; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6134 = 3'h3 == state ? tag_1_12 : _GEN_5618; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6135 = 3'h3 == state ? tag_1_13 : _GEN_5619; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6136 = 3'h3 == state ? tag_1_14 : _GEN_5620; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6137 = 3'h3 == state ? tag_1_15 : _GEN_5621; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6138 = 3'h3 == state ? tag_1_16 : _GEN_5622; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6139 = 3'h3 == state ? tag_1_17 : _GEN_5623; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6140 = 3'h3 == state ? tag_1_18 : _GEN_5624; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6141 = 3'h3 == state ? tag_1_19 : _GEN_5625; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6142 = 3'h3 == state ? tag_1_20 : _GEN_5626; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6143 = 3'h3 == state ? tag_1_21 : _GEN_5627; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6144 = 3'h3 == state ? tag_1_22 : _GEN_5628; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6145 = 3'h3 == state ? tag_1_23 : _GEN_5629; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6146 = 3'h3 == state ? tag_1_24 : _GEN_5630; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6147 = 3'h3 == state ? tag_1_25 : _GEN_5631; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6148 = 3'h3 == state ? tag_1_26 : _GEN_5632; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6149 = 3'h3 == state ? tag_1_27 : _GEN_5633; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6150 = 3'h3 == state ? tag_1_28 : _GEN_5634; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6151 = 3'h3 == state ? tag_1_29 : _GEN_5635; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6152 = 3'h3 == state ? tag_1_30 : _GEN_5636; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6153 = 3'h3 == state ? tag_1_31 : _GEN_5637; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6154 = 3'h3 == state ? tag_1_32 : _GEN_5638; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6155 = 3'h3 == state ? tag_1_33 : _GEN_5639; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6156 = 3'h3 == state ? tag_1_34 : _GEN_5640; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6157 = 3'h3 == state ? tag_1_35 : _GEN_5641; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6158 = 3'h3 == state ? tag_1_36 : _GEN_5642; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6159 = 3'h3 == state ? tag_1_37 : _GEN_5643; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6160 = 3'h3 == state ? tag_1_38 : _GEN_5644; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6161 = 3'h3 == state ? tag_1_39 : _GEN_5645; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6162 = 3'h3 == state ? tag_1_40 : _GEN_5646; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6163 = 3'h3 == state ? tag_1_41 : _GEN_5647; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6164 = 3'h3 == state ? tag_1_42 : _GEN_5648; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6165 = 3'h3 == state ? tag_1_43 : _GEN_5649; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6166 = 3'h3 == state ? tag_1_44 : _GEN_5650; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6167 = 3'h3 == state ? tag_1_45 : _GEN_5651; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6168 = 3'h3 == state ? tag_1_46 : _GEN_5652; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6169 = 3'h3 == state ? tag_1_47 : _GEN_5653; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6170 = 3'h3 == state ? tag_1_48 : _GEN_5654; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6171 = 3'h3 == state ? tag_1_49 : _GEN_5655; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6172 = 3'h3 == state ? tag_1_50 : _GEN_5656; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6173 = 3'h3 == state ? tag_1_51 : _GEN_5657; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6174 = 3'h3 == state ? tag_1_52 : _GEN_5658; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6175 = 3'h3 == state ? tag_1_53 : _GEN_5659; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6176 = 3'h3 == state ? tag_1_54 : _GEN_5660; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6177 = 3'h3 == state ? tag_1_55 : _GEN_5661; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6178 = 3'h3 == state ? tag_1_56 : _GEN_5662; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6179 = 3'h3 == state ? tag_1_57 : _GEN_5663; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6180 = 3'h3 == state ? tag_1_58 : _GEN_5664; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6181 = 3'h3 == state ? tag_1_59 : _GEN_5665; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6182 = 3'h3 == state ? tag_1_60 : _GEN_5666; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6183 = 3'h3 == state ? tag_1_61 : _GEN_5667; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6184 = 3'h3 == state ? tag_1_62 : _GEN_5668; // @[d_cache.scala 81:18 23:24]
  wire [31:0] _GEN_6185 = 3'h3 == state ? tag_1_63 : _GEN_5669; // @[d_cache.scala 81:18 23:24]
  wire  _GEN_6186 = 3'h3 == state ? valid_1_0 : _GEN_5670; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6187 = 3'h3 == state ? valid_1_1 : _GEN_5671; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6188 = 3'h3 == state ? valid_1_2 : _GEN_5672; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6189 = 3'h3 == state ? valid_1_3 : _GEN_5673; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6190 = 3'h3 == state ? valid_1_4 : _GEN_5674; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6191 = 3'h3 == state ? valid_1_5 : _GEN_5675; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6192 = 3'h3 == state ? valid_1_6 : _GEN_5676; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6193 = 3'h3 == state ? valid_1_7 : _GEN_5677; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6194 = 3'h3 == state ? valid_1_8 : _GEN_5678; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6195 = 3'h3 == state ? valid_1_9 : _GEN_5679; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6196 = 3'h3 == state ? valid_1_10 : _GEN_5680; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6197 = 3'h3 == state ? valid_1_11 : _GEN_5681; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6198 = 3'h3 == state ? valid_1_12 : _GEN_5682; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6199 = 3'h3 == state ? valid_1_13 : _GEN_5683; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6200 = 3'h3 == state ? valid_1_14 : _GEN_5684; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6201 = 3'h3 == state ? valid_1_15 : _GEN_5685; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6202 = 3'h3 == state ? valid_1_16 : _GEN_5686; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6203 = 3'h3 == state ? valid_1_17 : _GEN_5687; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6204 = 3'h3 == state ? valid_1_18 : _GEN_5688; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6205 = 3'h3 == state ? valid_1_19 : _GEN_5689; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6206 = 3'h3 == state ? valid_1_20 : _GEN_5690; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6207 = 3'h3 == state ? valid_1_21 : _GEN_5691; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6208 = 3'h3 == state ? valid_1_22 : _GEN_5692; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6209 = 3'h3 == state ? valid_1_23 : _GEN_5693; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6210 = 3'h3 == state ? valid_1_24 : _GEN_5694; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6211 = 3'h3 == state ? valid_1_25 : _GEN_5695; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6212 = 3'h3 == state ? valid_1_26 : _GEN_5696; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6213 = 3'h3 == state ? valid_1_27 : _GEN_5697; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6214 = 3'h3 == state ? valid_1_28 : _GEN_5698; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6215 = 3'h3 == state ? valid_1_29 : _GEN_5699; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6216 = 3'h3 == state ? valid_1_30 : _GEN_5700; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6217 = 3'h3 == state ? valid_1_31 : _GEN_5701; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6218 = 3'h3 == state ? valid_1_32 : _GEN_5702; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6219 = 3'h3 == state ? valid_1_33 : _GEN_5703; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6220 = 3'h3 == state ? valid_1_34 : _GEN_5704; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6221 = 3'h3 == state ? valid_1_35 : _GEN_5705; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6222 = 3'h3 == state ? valid_1_36 : _GEN_5706; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6223 = 3'h3 == state ? valid_1_37 : _GEN_5707; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6224 = 3'h3 == state ? valid_1_38 : _GEN_5708; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6225 = 3'h3 == state ? valid_1_39 : _GEN_5709; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6226 = 3'h3 == state ? valid_1_40 : _GEN_5710; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6227 = 3'h3 == state ? valid_1_41 : _GEN_5711; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6228 = 3'h3 == state ? valid_1_42 : _GEN_5712; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6229 = 3'h3 == state ? valid_1_43 : _GEN_5713; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6230 = 3'h3 == state ? valid_1_44 : _GEN_5714; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6231 = 3'h3 == state ? valid_1_45 : _GEN_5715; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6232 = 3'h3 == state ? valid_1_46 : _GEN_5716; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6233 = 3'h3 == state ? valid_1_47 : _GEN_5717; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6234 = 3'h3 == state ? valid_1_48 : _GEN_5718; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6235 = 3'h3 == state ? valid_1_49 : _GEN_5719; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6236 = 3'h3 == state ? valid_1_50 : _GEN_5720; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6237 = 3'h3 == state ? valid_1_51 : _GEN_5721; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6238 = 3'h3 == state ? valid_1_52 : _GEN_5722; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6239 = 3'h3 == state ? valid_1_53 : _GEN_5723; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6240 = 3'h3 == state ? valid_1_54 : _GEN_5724; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6241 = 3'h3 == state ? valid_1_55 : _GEN_5725; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6242 = 3'h3 == state ? valid_1_56 : _GEN_5726; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6243 = 3'h3 == state ? valid_1_57 : _GEN_5727; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6244 = 3'h3 == state ? valid_1_58 : _GEN_5728; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6245 = 3'h3 == state ? valid_1_59 : _GEN_5729; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6246 = 3'h3 == state ? valid_1_60 : _GEN_5730; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6247 = 3'h3 == state ? valid_1_61 : _GEN_5731; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6248 = 3'h3 == state ? valid_1_62 : _GEN_5732; // @[d_cache.scala 81:18 25:26]
  wire  _GEN_6249 = 3'h3 == state ? valid_1_63 : _GEN_5733; // @[d_cache.scala 81:18 25:26]
  wire [63:0] _GEN_6250 = 3'h3 == state ? write_back_data : _GEN_5734; // @[d_cache.scala 81:18 31:34]
  wire [40:0] _GEN_6251 = 3'h3 == state ? {{9'd0}, write_back_addr} : _GEN_5735; // @[d_cache.scala 81:18 32:34]
  wire  _GEN_6252 = 3'h3 == state ? dirty_0_0 : _GEN_5736; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6253 = 3'h3 == state ? dirty_0_1 : _GEN_5737; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6254 = 3'h3 == state ? dirty_0_2 : _GEN_5738; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6255 = 3'h3 == state ? dirty_0_3 : _GEN_5739; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6256 = 3'h3 == state ? dirty_0_4 : _GEN_5740; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6257 = 3'h3 == state ? dirty_0_5 : _GEN_5741; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6258 = 3'h3 == state ? dirty_0_6 : _GEN_5742; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6259 = 3'h3 == state ? dirty_0_7 : _GEN_5743; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6260 = 3'h3 == state ? dirty_0_8 : _GEN_5744; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6261 = 3'h3 == state ? dirty_0_9 : _GEN_5745; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6262 = 3'h3 == state ? dirty_0_10 : _GEN_5746; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6263 = 3'h3 == state ? dirty_0_11 : _GEN_5747; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6264 = 3'h3 == state ? dirty_0_12 : _GEN_5748; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6265 = 3'h3 == state ? dirty_0_13 : _GEN_5749; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6266 = 3'h3 == state ? dirty_0_14 : _GEN_5750; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6267 = 3'h3 == state ? dirty_0_15 : _GEN_5751; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6268 = 3'h3 == state ? dirty_0_16 : _GEN_5752; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6269 = 3'h3 == state ? dirty_0_17 : _GEN_5753; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6270 = 3'h3 == state ? dirty_0_18 : _GEN_5754; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6271 = 3'h3 == state ? dirty_0_19 : _GEN_5755; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6272 = 3'h3 == state ? dirty_0_20 : _GEN_5756; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6273 = 3'h3 == state ? dirty_0_21 : _GEN_5757; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6274 = 3'h3 == state ? dirty_0_22 : _GEN_5758; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6275 = 3'h3 == state ? dirty_0_23 : _GEN_5759; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6276 = 3'h3 == state ? dirty_0_24 : _GEN_5760; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6277 = 3'h3 == state ? dirty_0_25 : _GEN_5761; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6278 = 3'h3 == state ? dirty_0_26 : _GEN_5762; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6279 = 3'h3 == state ? dirty_0_27 : _GEN_5763; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6280 = 3'h3 == state ? dirty_0_28 : _GEN_5764; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6281 = 3'h3 == state ? dirty_0_29 : _GEN_5765; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6282 = 3'h3 == state ? dirty_0_30 : _GEN_5766; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6283 = 3'h3 == state ? dirty_0_31 : _GEN_5767; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6284 = 3'h3 == state ? dirty_0_32 : _GEN_5768; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6285 = 3'h3 == state ? dirty_0_33 : _GEN_5769; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6286 = 3'h3 == state ? dirty_0_34 : _GEN_5770; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6287 = 3'h3 == state ? dirty_0_35 : _GEN_5771; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6288 = 3'h3 == state ? dirty_0_36 : _GEN_5772; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6289 = 3'h3 == state ? dirty_0_37 : _GEN_5773; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6290 = 3'h3 == state ? dirty_0_38 : _GEN_5774; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6291 = 3'h3 == state ? dirty_0_39 : _GEN_5775; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6292 = 3'h3 == state ? dirty_0_40 : _GEN_5776; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6293 = 3'h3 == state ? dirty_0_41 : _GEN_5777; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6294 = 3'h3 == state ? dirty_0_42 : _GEN_5778; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6295 = 3'h3 == state ? dirty_0_43 : _GEN_5779; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6296 = 3'h3 == state ? dirty_0_44 : _GEN_5780; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6297 = 3'h3 == state ? dirty_0_45 : _GEN_5781; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6298 = 3'h3 == state ? dirty_0_46 : _GEN_5782; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6299 = 3'h3 == state ? dirty_0_47 : _GEN_5783; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6300 = 3'h3 == state ? dirty_0_48 : _GEN_5784; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6301 = 3'h3 == state ? dirty_0_49 : _GEN_5785; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6302 = 3'h3 == state ? dirty_0_50 : _GEN_5786; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6303 = 3'h3 == state ? dirty_0_51 : _GEN_5787; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6304 = 3'h3 == state ? dirty_0_52 : _GEN_5788; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6305 = 3'h3 == state ? dirty_0_53 : _GEN_5789; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6306 = 3'h3 == state ? dirty_0_54 : _GEN_5790; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6307 = 3'h3 == state ? dirty_0_55 : _GEN_5791; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6308 = 3'h3 == state ? dirty_0_56 : _GEN_5792; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6309 = 3'h3 == state ? dirty_0_57 : _GEN_5793; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6310 = 3'h3 == state ? dirty_0_58 : _GEN_5794; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6311 = 3'h3 == state ? dirty_0_59 : _GEN_5795; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6312 = 3'h3 == state ? dirty_0_60 : _GEN_5796; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6313 = 3'h3 == state ? dirty_0_61 : _GEN_5797; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6314 = 3'h3 == state ? dirty_0_62 : _GEN_5798; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6315 = 3'h3 == state ? dirty_0_63 : _GEN_5799; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_6316 = 3'h3 == state ? dirty_1_0 : _GEN_5800; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6317 = 3'h3 == state ? dirty_1_1 : _GEN_5801; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6318 = 3'h3 == state ? dirty_1_2 : _GEN_5802; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6319 = 3'h3 == state ? dirty_1_3 : _GEN_5803; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6320 = 3'h3 == state ? dirty_1_4 : _GEN_5804; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6321 = 3'h3 == state ? dirty_1_5 : _GEN_5805; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6322 = 3'h3 == state ? dirty_1_6 : _GEN_5806; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6323 = 3'h3 == state ? dirty_1_7 : _GEN_5807; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6324 = 3'h3 == state ? dirty_1_8 : _GEN_5808; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6325 = 3'h3 == state ? dirty_1_9 : _GEN_5809; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6326 = 3'h3 == state ? dirty_1_10 : _GEN_5810; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6327 = 3'h3 == state ? dirty_1_11 : _GEN_5811; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6328 = 3'h3 == state ? dirty_1_12 : _GEN_5812; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6329 = 3'h3 == state ? dirty_1_13 : _GEN_5813; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6330 = 3'h3 == state ? dirty_1_14 : _GEN_5814; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6331 = 3'h3 == state ? dirty_1_15 : _GEN_5815; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6332 = 3'h3 == state ? dirty_1_16 : _GEN_5816; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6333 = 3'h3 == state ? dirty_1_17 : _GEN_5817; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6334 = 3'h3 == state ? dirty_1_18 : _GEN_5818; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6335 = 3'h3 == state ? dirty_1_19 : _GEN_5819; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6336 = 3'h3 == state ? dirty_1_20 : _GEN_5820; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6337 = 3'h3 == state ? dirty_1_21 : _GEN_5821; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6338 = 3'h3 == state ? dirty_1_22 : _GEN_5822; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6339 = 3'h3 == state ? dirty_1_23 : _GEN_5823; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6340 = 3'h3 == state ? dirty_1_24 : _GEN_5824; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6341 = 3'h3 == state ? dirty_1_25 : _GEN_5825; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6342 = 3'h3 == state ? dirty_1_26 : _GEN_5826; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6343 = 3'h3 == state ? dirty_1_27 : _GEN_5827; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6344 = 3'h3 == state ? dirty_1_28 : _GEN_5828; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6345 = 3'h3 == state ? dirty_1_29 : _GEN_5829; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6346 = 3'h3 == state ? dirty_1_30 : _GEN_5830; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6347 = 3'h3 == state ? dirty_1_31 : _GEN_5831; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6348 = 3'h3 == state ? dirty_1_32 : _GEN_5832; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6349 = 3'h3 == state ? dirty_1_33 : _GEN_5833; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6350 = 3'h3 == state ? dirty_1_34 : _GEN_5834; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6351 = 3'h3 == state ? dirty_1_35 : _GEN_5835; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6352 = 3'h3 == state ? dirty_1_36 : _GEN_5836; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6353 = 3'h3 == state ? dirty_1_37 : _GEN_5837; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6354 = 3'h3 == state ? dirty_1_38 : _GEN_5838; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6355 = 3'h3 == state ? dirty_1_39 : _GEN_5839; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6356 = 3'h3 == state ? dirty_1_40 : _GEN_5840; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6357 = 3'h3 == state ? dirty_1_41 : _GEN_5841; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6358 = 3'h3 == state ? dirty_1_42 : _GEN_5842; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6359 = 3'h3 == state ? dirty_1_43 : _GEN_5843; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6360 = 3'h3 == state ? dirty_1_44 : _GEN_5844; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6361 = 3'h3 == state ? dirty_1_45 : _GEN_5845; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6362 = 3'h3 == state ? dirty_1_46 : _GEN_5846; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6363 = 3'h3 == state ? dirty_1_47 : _GEN_5847; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6364 = 3'h3 == state ? dirty_1_48 : _GEN_5848; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6365 = 3'h3 == state ? dirty_1_49 : _GEN_5849; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6366 = 3'h3 == state ? dirty_1_50 : _GEN_5850; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6367 = 3'h3 == state ? dirty_1_51 : _GEN_5851; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6368 = 3'h3 == state ? dirty_1_52 : _GEN_5852; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6369 = 3'h3 == state ? dirty_1_53 : _GEN_5853; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6370 = 3'h3 == state ? dirty_1_54 : _GEN_5854; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6371 = 3'h3 == state ? dirty_1_55 : _GEN_5855; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6372 = 3'h3 == state ? dirty_1_56 : _GEN_5856; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6373 = 3'h3 == state ? dirty_1_57 : _GEN_5857; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6374 = 3'h3 == state ? dirty_1_58 : _GEN_5858; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6375 = 3'h3 == state ? dirty_1_59 : _GEN_5859; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6376 = 3'h3 == state ? dirty_1_60 : _GEN_5860; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6377 = 3'h3 == state ? dirty_1_61 : _GEN_5861; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6378 = 3'h3 == state ? dirty_1_62 : _GEN_5862; // @[d_cache.scala 81:18 27:26]
  wire  _GEN_6379 = 3'h3 == state ? dirty_1_63 : _GEN_5863; // @[d_cache.scala 81:18 27:26]
  wire [40:0] _GEN_6896 = 3'h2 == state ? {{9'd0}, write_back_addr} : _GEN_6251; // @[d_cache.scala 81:18 32:34]
  wire [40:0] _GEN_7413 = 3'h1 == state ? {{9'd0}, write_back_addr} : _GEN_6896; // @[d_cache.scala 81:18 32:34]
  wire [40:0] _GEN_7930 = 3'h0 == state ? {{9'd0}, write_back_addr} : _GEN_7413; // @[d_cache.scala 81:18 32:34]
  wire [63:0] _io_to_lsu_rdata_T = _GEN_456 >> shift_bit; // @[d_cache.scala 228:49]
  wire [63:0] _io_to_lsu_rdata_T_1 = _GEN_712 >> shift_bit; // @[d_cache.scala 235:49]
  wire [63:0] _GEN_7931 = way1_hit ? _io_to_lsu_rdata_T_1 : 64'h0; // @[d_cache.scala 234:33 235:33 242:33]
  wire [63:0] _GEN_7935 = way0_hit ? _io_to_lsu_rdata_T : _GEN_7931; // @[d_cache.scala 227:23 228:33]
  wire  _GEN_7937 = way0_hit | way1_hit; // @[d_cache.scala 227:23 230:34]
  wire  _GEN_7939 = way1_hit ? 1'h0 : 1'h1; // @[d_cache.scala 266:33 268:35 275:35]
  wire  _GEN_7940 = way0_hit ? 1'h0 : _GEN_7939; // @[d_cache.scala 259:23 261:35]
  wire  _T_34 = state == 3'h3; // @[d_cache.scala 281:21]
  wire [63:0] _GEN_8673 = {{32'd0}, io_from_lsu_araddr}; // @[d_cache.scala 289:48]
  wire [63:0] _io_to_axi_araddr_T = _GEN_8673 & 64'hfffffffffffffff8; // @[d_cache.scala 289:48]
  wire  _T_37 = state == 3'h6; // @[d_cache.scala 330:21]
  wire [31:0] _GEN_7943 = state == 3'h6 ? 32'h0 : io_from_lsu_araddr; // @[d_cache.scala 330:35 338:26 354:26]
  wire  _GEN_7944 = state == 3'h6 ? 1'h0 : io_from_lsu_rready; // @[d_cache.scala 330:35 339:26 355:26]
  wire [31:0] _GEN_7945 = state == 3'h6 ? write_back_addr : 32'h0; // @[d_cache.scala 330:35 340:26 356:26]
  wire [63:0] _GEN_7946 = state == 3'h6 ? write_back_data : 64'h0; // @[d_cache.scala 330:35 342:25 358:25]
  wire [7:0] _GEN_7947 = state == 3'h6 ? 8'hff : 8'h0; // @[d_cache.scala 330:35 343:25 359:25]
  wire  _GEN_7949 = state == 3'h5 | _T_37; // @[d_cache.scala 314:31 316:27]
  wire [31:0] _GEN_7950 = state == 3'h5 ? io_from_lsu_araddr : _GEN_7943; // @[d_cache.scala 314:31 322:26]
  wire  _GEN_7951 = state == 3'h5 ? io_from_lsu_rready : _GEN_7944; // @[d_cache.scala 314:31 323:26]
  wire [31:0] _GEN_7952 = state == 3'h5 ? 32'h0 : _GEN_7945; // @[d_cache.scala 314:31 324:26]
  wire  _GEN_7953 = state == 3'h5 ? 1'h0 : _T_37; // @[d_cache.scala 314:31 325:27]
  wire [63:0] _GEN_7954 = state == 3'h5 ? 64'h0 : _GEN_7946; // @[d_cache.scala 314:31 326:25]
  wire [7:0] _GEN_7955 = state == 3'h5 ? 8'h0 : _GEN_7947; // @[d_cache.scala 314:31 327:25]
  wire  _GEN_7957 = state == 3'h4 | _GEN_7949; // @[d_cache.scala 297:31 299:27]
  wire  _GEN_7958 = state == 3'h4 & io_from_axi_wready; // @[d_cache.scala 297:31 301:26]
  wire  _GEN_7959 = state == 3'h4 & io_from_axi_bvalid; // @[d_cache.scala 297:31 302:26]
  wire  _GEN_7960 = state == 3'h4 & io_from_axi_awready; // @[d_cache.scala 297:31 303:27]
  wire [31:0] _GEN_7961 = state == 3'h4 ? 32'h0 : _GEN_7950; // @[d_cache.scala 297:31 305:26]
  wire  _GEN_7962 = state == 3'h4 ? io_from_lsu_rready : _GEN_7951; // @[d_cache.scala 297:31 306:26]
  wire [31:0] _GEN_7963 = state == 3'h4 ? io_from_lsu_awaddr : _GEN_7952; // @[d_cache.scala 297:31 307:26]
  wire  _GEN_7964 = state == 3'h4 ? io_from_lsu_awvalid : _GEN_7953; // @[d_cache.scala 297:31 308:27]
  wire [63:0] _GEN_7965 = state == 3'h4 ? {{32'd0}, io_from_lsu_wdata} : _GEN_7954; // @[d_cache.scala 297:31 309:25]
  wire [7:0] _GEN_7966 = state == 3'h4 ? io_from_lsu_wstrb : _GEN_7955; // @[d_cache.scala 297:31 310:25]
  wire  _GEN_7967 = state == 3'h4 ? io_from_lsu_wvalid : _GEN_7953; // @[d_cache.scala 297:31 311:26]
  wire  _GEN_7968 = state == 3'h4 ? io_from_lsu_bready : _GEN_7953; // @[d_cache.scala 297:31 312:26]
  wire  _GEN_7970 = state == 3'h3 | _GEN_7957; // @[d_cache.scala 281:31 283:27]
  wire  _GEN_7971 = state == 3'h3 ? 1'h0 : _GEN_7958; // @[d_cache.scala 281:31 285:26]
  wire  _GEN_7972 = state == 3'h3 ? 1'h0 : _GEN_7959; // @[d_cache.scala 281:31 286:26]
  wire  _GEN_7973 = state == 3'h3 ? 1'h0 : _GEN_7960; // @[d_cache.scala 281:31 287:27]
  wire [63:0] _GEN_7975 = state == 3'h3 ? _io_to_axi_araddr_T : {{32'd0}, _GEN_7961}; // @[d_cache.scala 281:31 289:26]
  wire  _GEN_7976 = state == 3'h3 ? io_from_lsu_rready : _GEN_7962; // @[d_cache.scala 281:31 290:26]
  wire [31:0] _GEN_7977 = state == 3'h3 ? 32'h0 : _GEN_7963; // @[d_cache.scala 281:31 291:26]
  wire  _GEN_7978 = state == 3'h3 ? 1'h0 : _GEN_7964; // @[d_cache.scala 281:31 292:27]
  wire [63:0] _GEN_7979 = state == 3'h3 ? 64'h0 : _GEN_7965; // @[d_cache.scala 281:31 293:25]
  wire [7:0] _GEN_7980 = state == 3'h3 ? 8'h0 : _GEN_7966; // @[d_cache.scala 281:31 294:25]
  wire  _GEN_7981 = state == 3'h3 ? 1'h0 : _GEN_7967; // @[d_cache.scala 281:31 295:26]
  wire  _GEN_7982 = state == 3'h3 ? 1'h0 : _GEN_7968; // @[d_cache.scala 281:31 296:26]
  wire  _GEN_7983 = state == 3'h2 ? 1'h0 : _T_34; // @[d_cache.scala 249:33 250:27]
  wire [63:0] _GEN_7984 = state == 3'h2 ? {{32'd0}, io_from_lsu_araddr} : _GEN_7975; // @[d_cache.scala 249:33 251:26]
  wire  _GEN_7985 = state == 3'h2 ? 1'h0 : _GEN_7976; // @[d_cache.scala 249:33 252:26]
  wire [31:0] _GEN_7986 = state == 3'h2 ? 32'h0 : _GEN_7977; // @[d_cache.scala 249:33 253:26]
  wire  _GEN_7987 = state == 3'h2 ? 1'h0 : _GEN_7978; // @[d_cache.scala 249:33 254:27]
  wire [63:0] _GEN_7988 = state == 3'h2 ? 64'h0 : _GEN_7979; // @[d_cache.scala 249:33 255:25]
  wire [7:0] _GEN_7989 = state == 3'h2 ? 8'h0 : _GEN_7980; // @[d_cache.scala 249:33 256:25]
  wire  _GEN_7990 = state == 3'h2 ? 1'h0 : _GEN_7981; // @[d_cache.scala 249:33 257:26]
  wire  _GEN_7991 = state == 3'h2 ? 1'h0 : _GEN_7982; // @[d_cache.scala 249:33 258:26]
  wire  _GEN_7993 = state == 3'h2 ? _GEN_7940 : _GEN_7970; // @[d_cache.scala 249:33]
  wire  _GEN_7994 = state == 3'h2 ? _GEN_7937 : _GEN_7971; // @[d_cache.scala 249:33]
  wire  _GEN_7995 = state == 3'h2 ? _GEN_7937 : _GEN_7973; // @[d_cache.scala 249:33]
  wire  _GEN_7996 = state == 3'h2 ? _GEN_7937 : _GEN_7972; // @[d_cache.scala 249:33]
  wire  _GEN_7997 = state == 3'h1 ? 1'h0 : _GEN_7983; // @[d_cache.scala 217:33 218:27]
  wire [63:0] _GEN_7998 = state == 3'h1 ? {{32'd0}, io_from_lsu_araddr} : _GEN_7984; // @[d_cache.scala 217:33 219:26]
  wire  _GEN_7999 = state == 3'h1 ? io_from_lsu_rready : _GEN_7985; // @[d_cache.scala 217:33 220:26]
  wire [31:0] _GEN_8000 = state == 3'h1 ? 32'h0 : _GEN_7986; // @[d_cache.scala 217:33 221:26]
  wire  _GEN_8001 = state == 3'h1 ? 1'h0 : _GEN_7987; // @[d_cache.scala 217:33 222:27]
  wire [63:0] _GEN_8002 = state == 3'h1 ? 64'h0 : _GEN_7988; // @[d_cache.scala 217:33 223:25]
  wire [7:0] _GEN_8003 = state == 3'h1 ? 8'h0 : _GEN_7989; // @[d_cache.scala 217:33 224:25]
  wire  _GEN_8004 = state == 3'h1 ? 1'h0 : _GEN_7990; // @[d_cache.scala 217:33 225:26]
  wire  _GEN_8005 = state == 3'h1 ? io_from_lsu_bready : _GEN_7991; // @[d_cache.scala 217:33 226:26]
  wire [63:0] _GEN_8006 = state == 3'h1 ? _GEN_7935 : 64'h0; // @[d_cache.scala 217:33]
  wire  _GEN_8007 = state == 3'h1 | _GEN_7993; // @[d_cache.scala 217:33]
  wire  _GEN_8008 = state == 3'h1 & _GEN_7937; // @[d_cache.scala 217:33]
  wire  _GEN_8009 = state == 3'h1 ? 1'h0 : _GEN_7994; // @[d_cache.scala 217:33]
  wire  _GEN_8010 = state == 3'h1 ? 1'h0 : _GEN_7995; // @[d_cache.scala 217:33]
  wire  _GEN_8011 = state == 3'h1 ? 1'h0 : _GEN_7996; // @[d_cache.scala 217:33]
  wire [63:0] _GEN_8019 = state == 3'h0 ? {{32'd0}, io_from_lsu_araddr} : _GEN_7998; // @[d_cache.scala 201:23 209:26]
  wire [63:0] _GEN_8023 = state == 3'h0 ? 64'h0 : _GEN_8002; // @[d_cache.scala 201:23 213:25]
  wire [40:0] _GEN_8674 = reset ? 41'h0 : _GEN_7930; // @[d_cache.scala 32:{34,34}]
  wire  _GEN_8676 = ~_T_14 & _T_15; // @[d_cache.scala 93:27]
  assign io_to_lsu_arready = state == 3'h0 ? io_from_axi_arready : _GEN_8007; // @[d_cache.scala 201:23 203:27]
  assign io_to_lsu_rdata = state == 3'h0 ? 64'h0 : _GEN_8006; // @[d_cache.scala 201:23 202:25]
  assign io_to_lsu_rvalid = state == 3'h0 ? 1'h0 : _GEN_8008; // @[d_cache.scala 201:23 204:26]
  assign io_to_lsu_awready = state == 3'h0 ? io_from_axi_awready : _GEN_8010; // @[d_cache.scala 201:23 207:27]
  assign io_to_lsu_wready = state == 3'h0 ? 1'h0 : _GEN_8009; // @[d_cache.scala 201:23 205:26]
  assign io_to_lsu_bvalid = state == 3'h0 ? 1'h0 : _GEN_8011; // @[d_cache.scala 201:23 206:26]
  assign io_to_axi_araddr = _GEN_8019[31:0];
  assign io_to_axi_arvalid = state == 3'h0 ? 1'h0 : _GEN_7997; // @[d_cache.scala 201:23 208:27]
  assign io_to_axi_rready = state == 3'h0 ? io_from_lsu_rready : _GEN_7999; // @[d_cache.scala 201:23 210:26]
  assign io_to_axi_awaddr = state == 3'h0 ? 32'h0 : _GEN_8000; // @[d_cache.scala 201:23 211:26]
  assign io_to_axi_awvalid = state == 3'h0 ? 1'h0 : _GEN_8001; // @[d_cache.scala 201:23 212:27]
  assign io_to_axi_wdata = _GEN_8023[31:0];
  assign io_to_axi_wstrb = state == 3'h0 ? 8'h0 : _GEN_8003; // @[d_cache.scala 201:23 214:25]
  assign io_to_axi_wvalid = state == 3'h0 ? 1'h0 : _GEN_8004; // @[d_cache.scala 201:23 215:26]
  assign io_to_axi_bready = state == 3'h0 ? io_from_lsu_bready : _GEN_8005; // @[d_cache.scala 201:23 216:26]
  always @(posedge clock) begin
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_0 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_0 <= _GEN_1100;
        end else begin
          ram_0_0 <= _GEN_5866;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_1 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_1 <= _GEN_1101;
        end else begin
          ram_0_1 <= _GEN_5867;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_2 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_2 <= _GEN_1102;
        end else begin
          ram_0_2 <= _GEN_5868;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_3 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_3 <= _GEN_1103;
        end else begin
          ram_0_3 <= _GEN_5869;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_4 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_4 <= _GEN_1104;
        end else begin
          ram_0_4 <= _GEN_5870;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_5 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_5 <= _GEN_1105;
        end else begin
          ram_0_5 <= _GEN_5871;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_6 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_6 <= _GEN_1106;
        end else begin
          ram_0_6 <= _GEN_5872;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_7 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_7 <= _GEN_1107;
        end else begin
          ram_0_7 <= _GEN_5873;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_8 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_8 <= _GEN_1108;
        end else begin
          ram_0_8 <= _GEN_5874;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_9 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_9 <= _GEN_1109;
        end else begin
          ram_0_9 <= _GEN_5875;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_10 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_10 <= _GEN_1110;
        end else begin
          ram_0_10 <= _GEN_5876;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_11 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_11 <= _GEN_1111;
        end else begin
          ram_0_11 <= _GEN_5877;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_12 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_12 <= _GEN_1112;
        end else begin
          ram_0_12 <= _GEN_5878;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_13 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_13 <= _GEN_1113;
        end else begin
          ram_0_13 <= _GEN_5879;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_14 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_14 <= _GEN_1114;
        end else begin
          ram_0_14 <= _GEN_5880;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_15 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_15 <= _GEN_1115;
        end else begin
          ram_0_15 <= _GEN_5881;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_16 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_16 <= _GEN_1116;
        end else begin
          ram_0_16 <= _GEN_5882;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_17 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_17 <= _GEN_1117;
        end else begin
          ram_0_17 <= _GEN_5883;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_18 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_18 <= _GEN_1118;
        end else begin
          ram_0_18 <= _GEN_5884;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_19 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_19 <= _GEN_1119;
        end else begin
          ram_0_19 <= _GEN_5885;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_20 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_20 <= _GEN_1120;
        end else begin
          ram_0_20 <= _GEN_5886;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_21 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_21 <= _GEN_1121;
        end else begin
          ram_0_21 <= _GEN_5887;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_22 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_22 <= _GEN_1122;
        end else begin
          ram_0_22 <= _GEN_5888;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_23 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_23 <= _GEN_1123;
        end else begin
          ram_0_23 <= _GEN_5889;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_24 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_24 <= _GEN_1124;
        end else begin
          ram_0_24 <= _GEN_5890;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_25 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_25 <= _GEN_1125;
        end else begin
          ram_0_25 <= _GEN_5891;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_26 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_26 <= _GEN_1126;
        end else begin
          ram_0_26 <= _GEN_5892;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_27 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_27 <= _GEN_1127;
        end else begin
          ram_0_27 <= _GEN_5893;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_28 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_28 <= _GEN_1128;
        end else begin
          ram_0_28 <= _GEN_5894;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_29 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_29 <= _GEN_1129;
        end else begin
          ram_0_29 <= _GEN_5895;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_30 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_30 <= _GEN_1130;
        end else begin
          ram_0_30 <= _GEN_5896;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_31 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_31 <= _GEN_1131;
        end else begin
          ram_0_31 <= _GEN_5897;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_32 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_32 <= _GEN_1132;
        end else begin
          ram_0_32 <= _GEN_5898;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_33 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_33 <= _GEN_1133;
        end else begin
          ram_0_33 <= _GEN_5899;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_34 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_34 <= _GEN_1134;
        end else begin
          ram_0_34 <= _GEN_5900;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_35 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_35 <= _GEN_1135;
        end else begin
          ram_0_35 <= _GEN_5901;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_36 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_36 <= _GEN_1136;
        end else begin
          ram_0_36 <= _GEN_5902;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_37 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_37 <= _GEN_1137;
        end else begin
          ram_0_37 <= _GEN_5903;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_38 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_38 <= _GEN_1138;
        end else begin
          ram_0_38 <= _GEN_5904;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_39 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_39 <= _GEN_1139;
        end else begin
          ram_0_39 <= _GEN_5905;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_40 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_40 <= _GEN_1140;
        end else begin
          ram_0_40 <= _GEN_5906;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_41 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_41 <= _GEN_1141;
        end else begin
          ram_0_41 <= _GEN_5907;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_42 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_42 <= _GEN_1142;
        end else begin
          ram_0_42 <= _GEN_5908;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_43 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_43 <= _GEN_1143;
        end else begin
          ram_0_43 <= _GEN_5909;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_44 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_44 <= _GEN_1144;
        end else begin
          ram_0_44 <= _GEN_5910;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_45 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_45 <= _GEN_1145;
        end else begin
          ram_0_45 <= _GEN_5911;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_46 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_46 <= _GEN_1146;
        end else begin
          ram_0_46 <= _GEN_5912;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_47 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_47 <= _GEN_1147;
        end else begin
          ram_0_47 <= _GEN_5913;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_48 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_48 <= _GEN_1148;
        end else begin
          ram_0_48 <= _GEN_5914;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_49 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_49 <= _GEN_1149;
        end else begin
          ram_0_49 <= _GEN_5915;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_50 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_50 <= _GEN_1150;
        end else begin
          ram_0_50 <= _GEN_5916;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_51 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_51 <= _GEN_1151;
        end else begin
          ram_0_51 <= _GEN_5917;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_52 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_52 <= _GEN_1152;
        end else begin
          ram_0_52 <= _GEN_5918;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_53 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_53 <= _GEN_1153;
        end else begin
          ram_0_53 <= _GEN_5919;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_54 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_54 <= _GEN_1154;
        end else begin
          ram_0_54 <= _GEN_5920;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_55 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_55 <= _GEN_1155;
        end else begin
          ram_0_55 <= _GEN_5921;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_56 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_56 <= _GEN_1156;
        end else begin
          ram_0_56 <= _GEN_5922;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_57 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_57 <= _GEN_1157;
        end else begin
          ram_0_57 <= _GEN_5923;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_58 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_58 <= _GEN_1158;
        end else begin
          ram_0_58 <= _GEN_5924;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_59 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_59 <= _GEN_1159;
        end else begin
          ram_0_59 <= _GEN_5925;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_60 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_60 <= _GEN_1160;
        end else begin
          ram_0_60 <= _GEN_5926;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_61 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_61 <= _GEN_1161;
        end else begin
          ram_0_61 <= _GEN_5927;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_62 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_62 <= _GEN_1162;
        end else begin
          ram_0_62 <= _GEN_5928;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_63 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_63 <= _GEN_1163;
        end else begin
          ram_0_63 <= _GEN_5929;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_0 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_0 <= _GEN_1293;
        end else begin
          ram_1_0 <= _GEN_6058;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_1 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_1 <= _GEN_1294;
        end else begin
          ram_1_1 <= _GEN_6059;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_2 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_2 <= _GEN_1295;
        end else begin
          ram_1_2 <= _GEN_6060;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_3 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_3 <= _GEN_1296;
        end else begin
          ram_1_3 <= _GEN_6061;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_4 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_4 <= _GEN_1297;
        end else begin
          ram_1_4 <= _GEN_6062;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_5 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_5 <= _GEN_1298;
        end else begin
          ram_1_5 <= _GEN_6063;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_6 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_6 <= _GEN_1299;
        end else begin
          ram_1_6 <= _GEN_6064;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_7 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_7 <= _GEN_1300;
        end else begin
          ram_1_7 <= _GEN_6065;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_8 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_8 <= _GEN_1301;
        end else begin
          ram_1_8 <= _GEN_6066;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_9 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_9 <= _GEN_1302;
        end else begin
          ram_1_9 <= _GEN_6067;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_10 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_10 <= _GEN_1303;
        end else begin
          ram_1_10 <= _GEN_6068;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_11 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_11 <= _GEN_1304;
        end else begin
          ram_1_11 <= _GEN_6069;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_12 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_12 <= _GEN_1305;
        end else begin
          ram_1_12 <= _GEN_6070;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_13 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_13 <= _GEN_1306;
        end else begin
          ram_1_13 <= _GEN_6071;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_14 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_14 <= _GEN_1307;
        end else begin
          ram_1_14 <= _GEN_6072;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_15 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_15 <= _GEN_1308;
        end else begin
          ram_1_15 <= _GEN_6073;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_16 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_16 <= _GEN_1309;
        end else begin
          ram_1_16 <= _GEN_6074;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_17 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_17 <= _GEN_1310;
        end else begin
          ram_1_17 <= _GEN_6075;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_18 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_18 <= _GEN_1311;
        end else begin
          ram_1_18 <= _GEN_6076;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_19 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_19 <= _GEN_1312;
        end else begin
          ram_1_19 <= _GEN_6077;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_20 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_20 <= _GEN_1313;
        end else begin
          ram_1_20 <= _GEN_6078;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_21 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_21 <= _GEN_1314;
        end else begin
          ram_1_21 <= _GEN_6079;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_22 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_22 <= _GEN_1315;
        end else begin
          ram_1_22 <= _GEN_6080;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_23 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_23 <= _GEN_1316;
        end else begin
          ram_1_23 <= _GEN_6081;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_24 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_24 <= _GEN_1317;
        end else begin
          ram_1_24 <= _GEN_6082;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_25 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_25 <= _GEN_1318;
        end else begin
          ram_1_25 <= _GEN_6083;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_26 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_26 <= _GEN_1319;
        end else begin
          ram_1_26 <= _GEN_6084;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_27 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_27 <= _GEN_1320;
        end else begin
          ram_1_27 <= _GEN_6085;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_28 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_28 <= _GEN_1321;
        end else begin
          ram_1_28 <= _GEN_6086;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_29 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_29 <= _GEN_1322;
        end else begin
          ram_1_29 <= _GEN_6087;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_30 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_30 <= _GEN_1323;
        end else begin
          ram_1_30 <= _GEN_6088;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_31 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_31 <= _GEN_1324;
        end else begin
          ram_1_31 <= _GEN_6089;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_32 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_32 <= _GEN_1325;
        end else begin
          ram_1_32 <= _GEN_6090;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_33 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_33 <= _GEN_1326;
        end else begin
          ram_1_33 <= _GEN_6091;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_34 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_34 <= _GEN_1327;
        end else begin
          ram_1_34 <= _GEN_6092;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_35 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_35 <= _GEN_1328;
        end else begin
          ram_1_35 <= _GEN_6093;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_36 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_36 <= _GEN_1329;
        end else begin
          ram_1_36 <= _GEN_6094;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_37 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_37 <= _GEN_1330;
        end else begin
          ram_1_37 <= _GEN_6095;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_38 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_38 <= _GEN_1331;
        end else begin
          ram_1_38 <= _GEN_6096;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_39 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_39 <= _GEN_1332;
        end else begin
          ram_1_39 <= _GEN_6097;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_40 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_40 <= _GEN_1333;
        end else begin
          ram_1_40 <= _GEN_6098;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_41 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_41 <= _GEN_1334;
        end else begin
          ram_1_41 <= _GEN_6099;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_42 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_42 <= _GEN_1335;
        end else begin
          ram_1_42 <= _GEN_6100;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_43 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_43 <= _GEN_1336;
        end else begin
          ram_1_43 <= _GEN_6101;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_44 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_44 <= _GEN_1337;
        end else begin
          ram_1_44 <= _GEN_6102;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_45 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_45 <= _GEN_1338;
        end else begin
          ram_1_45 <= _GEN_6103;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_46 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_46 <= _GEN_1339;
        end else begin
          ram_1_46 <= _GEN_6104;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_47 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_47 <= _GEN_1340;
        end else begin
          ram_1_47 <= _GEN_6105;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_48 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_48 <= _GEN_1341;
        end else begin
          ram_1_48 <= _GEN_6106;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_49 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_49 <= _GEN_1342;
        end else begin
          ram_1_49 <= _GEN_6107;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_50 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_50 <= _GEN_1343;
        end else begin
          ram_1_50 <= _GEN_6108;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_51 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_51 <= _GEN_1344;
        end else begin
          ram_1_51 <= _GEN_6109;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_52 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_52 <= _GEN_1345;
        end else begin
          ram_1_52 <= _GEN_6110;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_53 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_53 <= _GEN_1346;
        end else begin
          ram_1_53 <= _GEN_6111;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_54 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_54 <= _GEN_1347;
        end else begin
          ram_1_54 <= _GEN_6112;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_55 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_55 <= _GEN_1348;
        end else begin
          ram_1_55 <= _GEN_6113;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_56 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_56 <= _GEN_1349;
        end else begin
          ram_1_56 <= _GEN_6114;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_57 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_57 <= _GEN_1350;
        end else begin
          ram_1_57 <= _GEN_6115;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_58 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_58 <= _GEN_1351;
        end else begin
          ram_1_58 <= _GEN_6116;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_59 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_59 <= _GEN_1352;
        end else begin
          ram_1_59 <= _GEN_6117;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_60 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_60 <= _GEN_1353;
        end else begin
          ram_1_60 <= _GEN_6118;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_61 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_61 <= _GEN_1354;
        end else begin
          ram_1_61 <= _GEN_6119;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_62 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_62 <= _GEN_1355;
        end else begin
          ram_1_62 <= _GEN_6120;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_63 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_1_63 <= _GEN_1356;
        end else begin
          ram_1_63 <= _GEN_6121;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_0 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_0 <= _GEN_5930;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_1 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_1 <= _GEN_5931;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_2 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_2 <= _GEN_5932;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_3 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_3 <= _GEN_5933;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_4 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_4 <= _GEN_5934;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_5 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_5 <= _GEN_5935;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_6 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_6 <= _GEN_5936;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_7 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_7 <= _GEN_5937;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_8 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_8 <= _GEN_5938;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_9 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_9 <= _GEN_5939;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_10 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_10 <= _GEN_5940;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_11 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_11 <= _GEN_5941;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_12 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_12 <= _GEN_5942;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_13 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_13 <= _GEN_5943;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_14 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_14 <= _GEN_5944;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_15 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_15 <= _GEN_5945;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_16 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_16 <= _GEN_5946;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_17 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_17 <= _GEN_5947;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_18 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_18 <= _GEN_5948;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_19 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_19 <= _GEN_5949;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_20 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_20 <= _GEN_5950;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_21 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_21 <= _GEN_5951;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_22 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_22 <= _GEN_5952;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_23 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_23 <= _GEN_5953;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_24 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_24 <= _GEN_5954;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_25 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_25 <= _GEN_5955;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_26 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_26 <= _GEN_5956;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_27 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_27 <= _GEN_5957;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_28 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_28 <= _GEN_5958;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_29 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_29 <= _GEN_5959;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_30 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_30 <= _GEN_5960;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_31 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_31 <= _GEN_5961;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_32 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_32 <= _GEN_5962;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_33 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_33 <= _GEN_5963;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_34 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_34 <= _GEN_5964;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_35 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_35 <= _GEN_5965;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_36 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_36 <= _GEN_5966;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_37 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_37 <= _GEN_5967;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_38 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_38 <= _GEN_5968;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_39 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_39 <= _GEN_5969;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_40 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_40 <= _GEN_5970;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_41 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_41 <= _GEN_5971;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_42 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_42 <= _GEN_5972;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_43 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_43 <= _GEN_5973;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_44 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_44 <= _GEN_5974;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_45 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_45 <= _GEN_5975;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_46 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_46 <= _GEN_5976;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_47 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_47 <= _GEN_5977;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_48 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_48 <= _GEN_5978;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_49 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_49 <= _GEN_5979;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_50 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_50 <= _GEN_5980;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_51 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_51 <= _GEN_5981;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_52 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_52 <= _GEN_5982;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_53 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_53 <= _GEN_5983;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_54 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_54 <= _GEN_5984;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_55 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_55 <= _GEN_5985;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_56 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_56 <= _GEN_5986;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_57 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_57 <= _GEN_5987;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_58 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_58 <= _GEN_5988;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_59 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_59 <= _GEN_5989;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_60 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_60 <= _GEN_5990;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_61 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_61 <= _GEN_5991;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_62 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_62 <= _GEN_5992;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_63 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_63 <= _GEN_5993;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_0 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_0 <= _GEN_6122;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_1 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_1 <= _GEN_6123;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_2 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_2 <= _GEN_6124;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_3 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_3 <= _GEN_6125;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_4 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_4 <= _GEN_6126;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_5 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_5 <= _GEN_6127;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_6 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_6 <= _GEN_6128;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_7 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_7 <= _GEN_6129;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_8 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_8 <= _GEN_6130;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_9 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_9 <= _GEN_6131;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_10 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_10 <= _GEN_6132;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_11 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_11 <= _GEN_6133;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_12 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_12 <= _GEN_6134;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_13 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_13 <= _GEN_6135;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_14 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_14 <= _GEN_6136;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_15 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_15 <= _GEN_6137;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_16 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_16 <= _GEN_6138;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_17 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_17 <= _GEN_6139;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_18 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_18 <= _GEN_6140;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_19 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_19 <= _GEN_6141;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_20 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_20 <= _GEN_6142;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_21 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_21 <= _GEN_6143;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_22 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_22 <= _GEN_6144;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_23 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_23 <= _GEN_6145;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_24 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_24 <= _GEN_6146;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_25 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_25 <= _GEN_6147;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_26 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_26 <= _GEN_6148;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_27 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_27 <= _GEN_6149;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_28 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_28 <= _GEN_6150;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_29 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_29 <= _GEN_6151;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_30 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_30 <= _GEN_6152;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_31 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_31 <= _GEN_6153;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_32 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_32 <= _GEN_6154;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_33 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_33 <= _GEN_6155;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_34 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_34 <= _GEN_6156;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_35 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_35 <= _GEN_6157;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_36 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_36 <= _GEN_6158;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_37 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_37 <= _GEN_6159;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_38 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_38 <= _GEN_6160;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_39 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_39 <= _GEN_6161;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_40 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_40 <= _GEN_6162;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_41 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_41 <= _GEN_6163;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_42 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_42 <= _GEN_6164;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_43 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_43 <= _GEN_6165;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_44 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_44 <= _GEN_6166;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_45 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_45 <= _GEN_6167;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_46 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_46 <= _GEN_6168;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_47 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_47 <= _GEN_6169;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_48 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_48 <= _GEN_6170;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_49 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_49 <= _GEN_6171;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_50 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_50 <= _GEN_6172;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_51 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_51 <= _GEN_6173;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_52 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_52 <= _GEN_6174;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_53 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_53 <= _GEN_6175;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_54 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_54 <= _GEN_6176;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_55 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_55 <= _GEN_6177;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_56 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_56 <= _GEN_6178;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_57 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_57 <= _GEN_6179;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_58 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_58 <= _GEN_6180;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_59 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_59 <= _GEN_6181;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_60 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_60 <= _GEN_6182;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_61 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_61 <= _GEN_6183;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_62 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_62 <= _GEN_6184;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_63 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_1_63 <= _GEN_6185;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_0 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_0 <= _GEN_1164;
        end else begin
          valid_0_0 <= _GEN_5994;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_1 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_1 <= _GEN_1165;
        end else begin
          valid_0_1 <= _GEN_5995;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_2 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_2 <= _GEN_1166;
        end else begin
          valid_0_2 <= _GEN_5996;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_3 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_3 <= _GEN_1167;
        end else begin
          valid_0_3 <= _GEN_5997;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_4 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_4 <= _GEN_1168;
        end else begin
          valid_0_4 <= _GEN_5998;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_5 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_5 <= _GEN_1169;
        end else begin
          valid_0_5 <= _GEN_5999;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_6 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_6 <= _GEN_1170;
        end else begin
          valid_0_6 <= _GEN_6000;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_7 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_7 <= _GEN_1171;
        end else begin
          valid_0_7 <= _GEN_6001;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_8 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_8 <= _GEN_1172;
        end else begin
          valid_0_8 <= _GEN_6002;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_9 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_9 <= _GEN_1173;
        end else begin
          valid_0_9 <= _GEN_6003;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_10 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_10 <= _GEN_1174;
        end else begin
          valid_0_10 <= _GEN_6004;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_11 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_11 <= _GEN_1175;
        end else begin
          valid_0_11 <= _GEN_6005;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_12 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_12 <= _GEN_1176;
        end else begin
          valid_0_12 <= _GEN_6006;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_13 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_13 <= _GEN_1177;
        end else begin
          valid_0_13 <= _GEN_6007;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_14 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_14 <= _GEN_1178;
        end else begin
          valid_0_14 <= _GEN_6008;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_15 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_15 <= _GEN_1179;
        end else begin
          valid_0_15 <= _GEN_6009;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_16 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_16 <= _GEN_1180;
        end else begin
          valid_0_16 <= _GEN_6010;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_17 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_17 <= _GEN_1181;
        end else begin
          valid_0_17 <= _GEN_6011;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_18 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_18 <= _GEN_1182;
        end else begin
          valid_0_18 <= _GEN_6012;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_19 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_19 <= _GEN_1183;
        end else begin
          valid_0_19 <= _GEN_6013;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_20 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_20 <= _GEN_1184;
        end else begin
          valid_0_20 <= _GEN_6014;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_21 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_21 <= _GEN_1185;
        end else begin
          valid_0_21 <= _GEN_6015;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_22 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_22 <= _GEN_1186;
        end else begin
          valid_0_22 <= _GEN_6016;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_23 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_23 <= _GEN_1187;
        end else begin
          valid_0_23 <= _GEN_6017;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_24 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_24 <= _GEN_1188;
        end else begin
          valid_0_24 <= _GEN_6018;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_25 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_25 <= _GEN_1189;
        end else begin
          valid_0_25 <= _GEN_6019;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_26 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_26 <= _GEN_1190;
        end else begin
          valid_0_26 <= _GEN_6020;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_27 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_27 <= _GEN_1191;
        end else begin
          valid_0_27 <= _GEN_6021;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_28 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_28 <= _GEN_1192;
        end else begin
          valid_0_28 <= _GEN_6022;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_29 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_29 <= _GEN_1193;
        end else begin
          valid_0_29 <= _GEN_6023;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_30 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_30 <= _GEN_1194;
        end else begin
          valid_0_30 <= _GEN_6024;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_31 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_31 <= _GEN_1195;
        end else begin
          valid_0_31 <= _GEN_6025;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_32 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_32 <= _GEN_1196;
        end else begin
          valid_0_32 <= _GEN_6026;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_33 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_33 <= _GEN_1197;
        end else begin
          valid_0_33 <= _GEN_6027;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_34 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_34 <= _GEN_1198;
        end else begin
          valid_0_34 <= _GEN_6028;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_35 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_35 <= _GEN_1199;
        end else begin
          valid_0_35 <= _GEN_6029;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_36 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_36 <= _GEN_1200;
        end else begin
          valid_0_36 <= _GEN_6030;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_37 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_37 <= _GEN_1201;
        end else begin
          valid_0_37 <= _GEN_6031;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_38 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_38 <= _GEN_1202;
        end else begin
          valid_0_38 <= _GEN_6032;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_39 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_39 <= _GEN_1203;
        end else begin
          valid_0_39 <= _GEN_6033;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_40 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_40 <= _GEN_1204;
        end else begin
          valid_0_40 <= _GEN_6034;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_41 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_41 <= _GEN_1205;
        end else begin
          valid_0_41 <= _GEN_6035;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_42 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_42 <= _GEN_1206;
        end else begin
          valid_0_42 <= _GEN_6036;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_43 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_43 <= _GEN_1207;
        end else begin
          valid_0_43 <= _GEN_6037;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_44 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_44 <= _GEN_1208;
        end else begin
          valid_0_44 <= _GEN_6038;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_45 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_45 <= _GEN_1209;
        end else begin
          valid_0_45 <= _GEN_6039;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_46 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_46 <= _GEN_1210;
        end else begin
          valid_0_46 <= _GEN_6040;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_47 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_47 <= _GEN_1211;
        end else begin
          valid_0_47 <= _GEN_6041;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_48 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_48 <= _GEN_1212;
        end else begin
          valid_0_48 <= _GEN_6042;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_49 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_49 <= _GEN_1213;
        end else begin
          valid_0_49 <= _GEN_6043;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_50 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_50 <= _GEN_1214;
        end else begin
          valid_0_50 <= _GEN_6044;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_51 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_51 <= _GEN_1215;
        end else begin
          valid_0_51 <= _GEN_6045;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_52 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_52 <= _GEN_1216;
        end else begin
          valid_0_52 <= _GEN_6046;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_53 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_53 <= _GEN_1217;
        end else begin
          valid_0_53 <= _GEN_6047;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_54 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_54 <= _GEN_1218;
        end else begin
          valid_0_54 <= _GEN_6048;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_55 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_55 <= _GEN_1219;
        end else begin
          valid_0_55 <= _GEN_6049;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_56 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_56 <= _GEN_1220;
        end else begin
          valid_0_56 <= _GEN_6050;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_57 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_57 <= _GEN_1221;
        end else begin
          valid_0_57 <= _GEN_6051;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_58 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_58 <= _GEN_1222;
        end else begin
          valid_0_58 <= _GEN_6052;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_59 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_59 <= _GEN_1223;
        end else begin
          valid_0_59 <= _GEN_6053;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_60 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_60 <= _GEN_1224;
        end else begin
          valid_0_60 <= _GEN_6054;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_61 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_61 <= _GEN_1225;
        end else begin
          valid_0_61 <= _GEN_6055;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_62 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_62 <= _GEN_1226;
        end else begin
          valid_0_62 <= _GEN_6056;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_63 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_63 <= _GEN_1227;
        end else begin
          valid_0_63 <= _GEN_6057;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_0 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_0 <= _GEN_1357;
        end else begin
          valid_1_0 <= _GEN_6186;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_1 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_1 <= _GEN_1358;
        end else begin
          valid_1_1 <= _GEN_6187;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_2 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_2 <= _GEN_1359;
        end else begin
          valid_1_2 <= _GEN_6188;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_3 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_3 <= _GEN_1360;
        end else begin
          valid_1_3 <= _GEN_6189;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_4 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_4 <= _GEN_1361;
        end else begin
          valid_1_4 <= _GEN_6190;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_5 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_5 <= _GEN_1362;
        end else begin
          valid_1_5 <= _GEN_6191;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_6 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_6 <= _GEN_1363;
        end else begin
          valid_1_6 <= _GEN_6192;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_7 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_7 <= _GEN_1364;
        end else begin
          valid_1_7 <= _GEN_6193;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_8 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_8 <= _GEN_1365;
        end else begin
          valid_1_8 <= _GEN_6194;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_9 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_9 <= _GEN_1366;
        end else begin
          valid_1_9 <= _GEN_6195;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_10 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_10 <= _GEN_1367;
        end else begin
          valid_1_10 <= _GEN_6196;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_11 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_11 <= _GEN_1368;
        end else begin
          valid_1_11 <= _GEN_6197;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_12 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_12 <= _GEN_1369;
        end else begin
          valid_1_12 <= _GEN_6198;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_13 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_13 <= _GEN_1370;
        end else begin
          valid_1_13 <= _GEN_6199;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_14 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_14 <= _GEN_1371;
        end else begin
          valid_1_14 <= _GEN_6200;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_15 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_15 <= _GEN_1372;
        end else begin
          valid_1_15 <= _GEN_6201;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_16 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_16 <= _GEN_1373;
        end else begin
          valid_1_16 <= _GEN_6202;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_17 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_17 <= _GEN_1374;
        end else begin
          valid_1_17 <= _GEN_6203;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_18 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_18 <= _GEN_1375;
        end else begin
          valid_1_18 <= _GEN_6204;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_19 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_19 <= _GEN_1376;
        end else begin
          valid_1_19 <= _GEN_6205;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_20 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_20 <= _GEN_1377;
        end else begin
          valid_1_20 <= _GEN_6206;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_21 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_21 <= _GEN_1378;
        end else begin
          valid_1_21 <= _GEN_6207;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_22 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_22 <= _GEN_1379;
        end else begin
          valid_1_22 <= _GEN_6208;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_23 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_23 <= _GEN_1380;
        end else begin
          valid_1_23 <= _GEN_6209;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_24 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_24 <= _GEN_1381;
        end else begin
          valid_1_24 <= _GEN_6210;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_25 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_25 <= _GEN_1382;
        end else begin
          valid_1_25 <= _GEN_6211;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_26 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_26 <= _GEN_1383;
        end else begin
          valid_1_26 <= _GEN_6212;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_27 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_27 <= _GEN_1384;
        end else begin
          valid_1_27 <= _GEN_6213;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_28 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_28 <= _GEN_1385;
        end else begin
          valid_1_28 <= _GEN_6214;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_29 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_29 <= _GEN_1386;
        end else begin
          valid_1_29 <= _GEN_6215;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_30 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_30 <= _GEN_1387;
        end else begin
          valid_1_30 <= _GEN_6216;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_31 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_31 <= _GEN_1388;
        end else begin
          valid_1_31 <= _GEN_6217;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_32 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_32 <= _GEN_1389;
        end else begin
          valid_1_32 <= _GEN_6218;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_33 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_33 <= _GEN_1390;
        end else begin
          valid_1_33 <= _GEN_6219;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_34 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_34 <= _GEN_1391;
        end else begin
          valid_1_34 <= _GEN_6220;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_35 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_35 <= _GEN_1392;
        end else begin
          valid_1_35 <= _GEN_6221;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_36 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_36 <= _GEN_1393;
        end else begin
          valid_1_36 <= _GEN_6222;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_37 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_37 <= _GEN_1394;
        end else begin
          valid_1_37 <= _GEN_6223;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_38 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_38 <= _GEN_1395;
        end else begin
          valid_1_38 <= _GEN_6224;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_39 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_39 <= _GEN_1396;
        end else begin
          valid_1_39 <= _GEN_6225;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_40 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_40 <= _GEN_1397;
        end else begin
          valid_1_40 <= _GEN_6226;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_41 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_41 <= _GEN_1398;
        end else begin
          valid_1_41 <= _GEN_6227;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_42 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_42 <= _GEN_1399;
        end else begin
          valid_1_42 <= _GEN_6228;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_43 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_43 <= _GEN_1400;
        end else begin
          valid_1_43 <= _GEN_6229;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_44 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_44 <= _GEN_1401;
        end else begin
          valid_1_44 <= _GEN_6230;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_45 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_45 <= _GEN_1402;
        end else begin
          valid_1_45 <= _GEN_6231;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_46 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_46 <= _GEN_1403;
        end else begin
          valid_1_46 <= _GEN_6232;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_47 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_47 <= _GEN_1404;
        end else begin
          valid_1_47 <= _GEN_6233;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_48 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_48 <= _GEN_1405;
        end else begin
          valid_1_48 <= _GEN_6234;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_49 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_49 <= _GEN_1406;
        end else begin
          valid_1_49 <= _GEN_6235;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_50 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_50 <= _GEN_1407;
        end else begin
          valid_1_50 <= _GEN_6236;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_51 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_51 <= _GEN_1408;
        end else begin
          valid_1_51 <= _GEN_6237;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_52 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_52 <= _GEN_1409;
        end else begin
          valid_1_52 <= _GEN_6238;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_53 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_53 <= _GEN_1410;
        end else begin
          valid_1_53 <= _GEN_6239;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_54 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_54 <= _GEN_1411;
        end else begin
          valid_1_54 <= _GEN_6240;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_55 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_55 <= _GEN_1412;
        end else begin
          valid_1_55 <= _GEN_6241;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_56 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_56 <= _GEN_1413;
        end else begin
          valid_1_56 <= _GEN_6242;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_57 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_57 <= _GEN_1414;
        end else begin
          valid_1_57 <= _GEN_6243;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_58 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_58 <= _GEN_1415;
        end else begin
          valid_1_58 <= _GEN_6244;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_59 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_59 <= _GEN_1416;
        end else begin
          valid_1_59 <= _GEN_6245;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_60 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_60 <= _GEN_1417;
        end else begin
          valid_1_60 <= _GEN_6246;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_61 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_61 <= _GEN_1418;
        end else begin
          valid_1_61 <= _GEN_6247;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_62 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_62 <= _GEN_1419;
        end else begin
          valid_1_62 <= _GEN_6248;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_63 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_1_63 <= _GEN_1420;
        end else begin
          valid_1_63 <= _GEN_6249;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_0 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_0 <= _GEN_1228;
        end else begin
          dirty_0_0 <= _GEN_6252;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_1 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_1 <= _GEN_1229;
        end else begin
          dirty_0_1 <= _GEN_6253;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_2 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_2 <= _GEN_1230;
        end else begin
          dirty_0_2 <= _GEN_6254;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_3 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_3 <= _GEN_1231;
        end else begin
          dirty_0_3 <= _GEN_6255;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_4 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_4 <= _GEN_1232;
        end else begin
          dirty_0_4 <= _GEN_6256;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_5 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_5 <= _GEN_1233;
        end else begin
          dirty_0_5 <= _GEN_6257;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_6 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_6 <= _GEN_1234;
        end else begin
          dirty_0_6 <= _GEN_6258;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_7 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_7 <= _GEN_1235;
        end else begin
          dirty_0_7 <= _GEN_6259;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_8 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_8 <= _GEN_1236;
        end else begin
          dirty_0_8 <= _GEN_6260;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_9 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_9 <= _GEN_1237;
        end else begin
          dirty_0_9 <= _GEN_6261;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_10 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_10 <= _GEN_1238;
        end else begin
          dirty_0_10 <= _GEN_6262;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_11 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_11 <= _GEN_1239;
        end else begin
          dirty_0_11 <= _GEN_6263;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_12 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_12 <= _GEN_1240;
        end else begin
          dirty_0_12 <= _GEN_6264;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_13 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_13 <= _GEN_1241;
        end else begin
          dirty_0_13 <= _GEN_6265;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_14 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_14 <= _GEN_1242;
        end else begin
          dirty_0_14 <= _GEN_6266;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_15 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_15 <= _GEN_1243;
        end else begin
          dirty_0_15 <= _GEN_6267;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_16 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_16 <= _GEN_1244;
        end else begin
          dirty_0_16 <= _GEN_6268;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_17 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_17 <= _GEN_1245;
        end else begin
          dirty_0_17 <= _GEN_6269;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_18 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_18 <= _GEN_1246;
        end else begin
          dirty_0_18 <= _GEN_6270;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_19 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_19 <= _GEN_1247;
        end else begin
          dirty_0_19 <= _GEN_6271;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_20 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_20 <= _GEN_1248;
        end else begin
          dirty_0_20 <= _GEN_6272;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_21 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_21 <= _GEN_1249;
        end else begin
          dirty_0_21 <= _GEN_6273;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_22 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_22 <= _GEN_1250;
        end else begin
          dirty_0_22 <= _GEN_6274;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_23 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_23 <= _GEN_1251;
        end else begin
          dirty_0_23 <= _GEN_6275;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_24 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_24 <= _GEN_1252;
        end else begin
          dirty_0_24 <= _GEN_6276;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_25 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_25 <= _GEN_1253;
        end else begin
          dirty_0_25 <= _GEN_6277;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_26 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_26 <= _GEN_1254;
        end else begin
          dirty_0_26 <= _GEN_6278;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_27 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_27 <= _GEN_1255;
        end else begin
          dirty_0_27 <= _GEN_6279;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_28 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_28 <= _GEN_1256;
        end else begin
          dirty_0_28 <= _GEN_6280;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_29 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_29 <= _GEN_1257;
        end else begin
          dirty_0_29 <= _GEN_6281;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_30 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_30 <= _GEN_1258;
        end else begin
          dirty_0_30 <= _GEN_6282;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_31 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_31 <= _GEN_1259;
        end else begin
          dirty_0_31 <= _GEN_6283;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_32 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_32 <= _GEN_1260;
        end else begin
          dirty_0_32 <= _GEN_6284;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_33 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_33 <= _GEN_1261;
        end else begin
          dirty_0_33 <= _GEN_6285;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_34 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_34 <= _GEN_1262;
        end else begin
          dirty_0_34 <= _GEN_6286;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_35 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_35 <= _GEN_1263;
        end else begin
          dirty_0_35 <= _GEN_6287;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_36 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_36 <= _GEN_1264;
        end else begin
          dirty_0_36 <= _GEN_6288;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_37 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_37 <= _GEN_1265;
        end else begin
          dirty_0_37 <= _GEN_6289;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_38 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_38 <= _GEN_1266;
        end else begin
          dirty_0_38 <= _GEN_6290;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_39 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_39 <= _GEN_1267;
        end else begin
          dirty_0_39 <= _GEN_6291;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_40 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_40 <= _GEN_1268;
        end else begin
          dirty_0_40 <= _GEN_6292;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_41 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_41 <= _GEN_1269;
        end else begin
          dirty_0_41 <= _GEN_6293;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_42 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_42 <= _GEN_1270;
        end else begin
          dirty_0_42 <= _GEN_6294;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_43 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_43 <= _GEN_1271;
        end else begin
          dirty_0_43 <= _GEN_6295;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_44 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_44 <= _GEN_1272;
        end else begin
          dirty_0_44 <= _GEN_6296;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_45 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_45 <= _GEN_1273;
        end else begin
          dirty_0_45 <= _GEN_6297;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_46 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_46 <= _GEN_1274;
        end else begin
          dirty_0_46 <= _GEN_6298;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_47 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_47 <= _GEN_1275;
        end else begin
          dirty_0_47 <= _GEN_6299;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_48 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_48 <= _GEN_1276;
        end else begin
          dirty_0_48 <= _GEN_6300;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_49 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_49 <= _GEN_1277;
        end else begin
          dirty_0_49 <= _GEN_6301;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_50 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_50 <= _GEN_1278;
        end else begin
          dirty_0_50 <= _GEN_6302;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_51 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_51 <= _GEN_1279;
        end else begin
          dirty_0_51 <= _GEN_6303;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_52 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_52 <= _GEN_1280;
        end else begin
          dirty_0_52 <= _GEN_6304;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_53 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_53 <= _GEN_1281;
        end else begin
          dirty_0_53 <= _GEN_6305;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_54 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_54 <= _GEN_1282;
        end else begin
          dirty_0_54 <= _GEN_6306;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_55 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_55 <= _GEN_1283;
        end else begin
          dirty_0_55 <= _GEN_6307;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_56 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_56 <= _GEN_1284;
        end else begin
          dirty_0_56 <= _GEN_6308;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_57 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_57 <= _GEN_1285;
        end else begin
          dirty_0_57 <= _GEN_6309;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_58 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_58 <= _GEN_1286;
        end else begin
          dirty_0_58 <= _GEN_6310;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_59 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_59 <= _GEN_1287;
        end else begin
          dirty_0_59 <= _GEN_6311;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_60 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_60 <= _GEN_1288;
        end else begin
          dirty_0_60 <= _GEN_6312;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_61 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_61 <= _GEN_1289;
        end else begin
          dirty_0_61 <= _GEN_6313;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_62 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_62 <= _GEN_1290;
        end else begin
          dirty_0_62 <= _GEN_6314;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_63 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_63 <= _GEN_1291;
        end else begin
          dirty_0_63 <= _GEN_6315;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_0 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_0 <= _GEN_1421;
        end else begin
          dirty_1_0 <= _GEN_6316;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_1 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_1 <= _GEN_1422;
        end else begin
          dirty_1_1 <= _GEN_6317;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_2 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_2 <= _GEN_1423;
        end else begin
          dirty_1_2 <= _GEN_6318;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_3 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_3 <= _GEN_1424;
        end else begin
          dirty_1_3 <= _GEN_6319;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_4 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_4 <= _GEN_1425;
        end else begin
          dirty_1_4 <= _GEN_6320;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_5 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_5 <= _GEN_1426;
        end else begin
          dirty_1_5 <= _GEN_6321;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_6 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_6 <= _GEN_1427;
        end else begin
          dirty_1_6 <= _GEN_6322;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_7 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_7 <= _GEN_1428;
        end else begin
          dirty_1_7 <= _GEN_6323;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_8 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_8 <= _GEN_1429;
        end else begin
          dirty_1_8 <= _GEN_6324;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_9 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_9 <= _GEN_1430;
        end else begin
          dirty_1_9 <= _GEN_6325;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_10 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_10 <= _GEN_1431;
        end else begin
          dirty_1_10 <= _GEN_6326;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_11 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_11 <= _GEN_1432;
        end else begin
          dirty_1_11 <= _GEN_6327;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_12 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_12 <= _GEN_1433;
        end else begin
          dirty_1_12 <= _GEN_6328;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_13 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_13 <= _GEN_1434;
        end else begin
          dirty_1_13 <= _GEN_6329;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_14 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_14 <= _GEN_1435;
        end else begin
          dirty_1_14 <= _GEN_6330;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_15 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_15 <= _GEN_1436;
        end else begin
          dirty_1_15 <= _GEN_6331;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_16 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_16 <= _GEN_1437;
        end else begin
          dirty_1_16 <= _GEN_6332;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_17 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_17 <= _GEN_1438;
        end else begin
          dirty_1_17 <= _GEN_6333;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_18 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_18 <= _GEN_1439;
        end else begin
          dirty_1_18 <= _GEN_6334;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_19 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_19 <= _GEN_1440;
        end else begin
          dirty_1_19 <= _GEN_6335;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_20 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_20 <= _GEN_1441;
        end else begin
          dirty_1_20 <= _GEN_6336;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_21 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_21 <= _GEN_1442;
        end else begin
          dirty_1_21 <= _GEN_6337;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_22 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_22 <= _GEN_1443;
        end else begin
          dirty_1_22 <= _GEN_6338;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_23 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_23 <= _GEN_1444;
        end else begin
          dirty_1_23 <= _GEN_6339;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_24 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_24 <= _GEN_1445;
        end else begin
          dirty_1_24 <= _GEN_6340;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_25 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_25 <= _GEN_1446;
        end else begin
          dirty_1_25 <= _GEN_6341;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_26 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_26 <= _GEN_1447;
        end else begin
          dirty_1_26 <= _GEN_6342;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_27 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_27 <= _GEN_1448;
        end else begin
          dirty_1_27 <= _GEN_6343;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_28 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_28 <= _GEN_1449;
        end else begin
          dirty_1_28 <= _GEN_6344;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_29 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_29 <= _GEN_1450;
        end else begin
          dirty_1_29 <= _GEN_6345;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_30 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_30 <= _GEN_1451;
        end else begin
          dirty_1_30 <= _GEN_6346;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_31 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_31 <= _GEN_1452;
        end else begin
          dirty_1_31 <= _GEN_6347;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_32 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_32 <= _GEN_1453;
        end else begin
          dirty_1_32 <= _GEN_6348;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_33 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_33 <= _GEN_1454;
        end else begin
          dirty_1_33 <= _GEN_6349;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_34 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_34 <= _GEN_1455;
        end else begin
          dirty_1_34 <= _GEN_6350;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_35 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_35 <= _GEN_1456;
        end else begin
          dirty_1_35 <= _GEN_6351;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_36 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_36 <= _GEN_1457;
        end else begin
          dirty_1_36 <= _GEN_6352;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_37 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_37 <= _GEN_1458;
        end else begin
          dirty_1_37 <= _GEN_6353;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_38 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_38 <= _GEN_1459;
        end else begin
          dirty_1_38 <= _GEN_6354;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_39 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_39 <= _GEN_1460;
        end else begin
          dirty_1_39 <= _GEN_6355;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_40 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_40 <= _GEN_1461;
        end else begin
          dirty_1_40 <= _GEN_6356;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_41 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_41 <= _GEN_1462;
        end else begin
          dirty_1_41 <= _GEN_6357;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_42 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_42 <= _GEN_1463;
        end else begin
          dirty_1_42 <= _GEN_6358;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_43 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_43 <= _GEN_1464;
        end else begin
          dirty_1_43 <= _GEN_6359;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_44 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_44 <= _GEN_1465;
        end else begin
          dirty_1_44 <= _GEN_6360;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_45 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_45 <= _GEN_1466;
        end else begin
          dirty_1_45 <= _GEN_6361;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_46 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_46 <= _GEN_1467;
        end else begin
          dirty_1_46 <= _GEN_6362;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_47 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_47 <= _GEN_1468;
        end else begin
          dirty_1_47 <= _GEN_6363;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_48 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_48 <= _GEN_1469;
        end else begin
          dirty_1_48 <= _GEN_6364;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_49 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_49 <= _GEN_1470;
        end else begin
          dirty_1_49 <= _GEN_6365;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_50 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_50 <= _GEN_1471;
        end else begin
          dirty_1_50 <= _GEN_6366;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_51 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_51 <= _GEN_1472;
        end else begin
          dirty_1_51 <= _GEN_6367;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_52 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_52 <= _GEN_1473;
        end else begin
          dirty_1_52 <= _GEN_6368;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_53 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_53 <= _GEN_1474;
        end else begin
          dirty_1_53 <= _GEN_6369;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_54 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_54 <= _GEN_1475;
        end else begin
          dirty_1_54 <= _GEN_6370;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_55 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_55 <= _GEN_1476;
        end else begin
          dirty_1_55 <= _GEN_6371;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_56 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_56 <= _GEN_1477;
        end else begin
          dirty_1_56 <= _GEN_6372;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_57 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_57 <= _GEN_1478;
        end else begin
          dirty_1_57 <= _GEN_6373;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_58 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_58 <= _GEN_1479;
        end else begin
          dirty_1_58 <= _GEN_6374;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_59 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_59 <= _GEN_1480;
        end else begin
          dirty_1_59 <= _GEN_6375;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_60 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_60 <= _GEN_1481;
        end else begin
          dirty_1_60 <= _GEN_6376;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_61 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_61 <= _GEN_1482;
        end else begin
          dirty_1_61 <= _GEN_6377;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_62 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_62 <= _GEN_1483;
        end else begin
          dirty_1_62 <= _GEN_6378;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_63 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_1_63 <= _GEN_1484;
        end else begin
          dirty_1_63 <= _GEN_6379;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:27]
      way0_hit <= 1'h0; // @[d_cache.scala 28:27]
    end else begin
      way0_hit <= _T_4;
    end
    if (reset) begin // @[d_cache.scala 29:27]
      way1_hit <= 1'h0; // @[d_cache.scala 29:27]
    end else begin
      way1_hit <= _T_7;
    end
    if (reset) begin // @[d_cache.scala 31:34]
      write_back_data <= 64'h0; // @[d_cache.scala 31:34]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          write_back_data <= _GEN_6250;
        end
      end
    end
    write_back_addr <= _GEN_8674[31:0]; // @[d_cache.scala 32:{34,34}]
    if (reset) begin // @[d_cache.scala 35:28]
      unuse_way <= 2'h0; // @[d_cache.scala 35:28]
    end else if (~_GEN_127) begin // @[d_cache.scala 68:31]
      unuse_way <= 2'h1; // @[d_cache.scala 69:19]
    end else if (~_GEN_256) begin // @[d_cache.scala 70:37]
      unuse_way <= 2'h2; // @[d_cache.scala 71:19]
    end else begin
      unuse_way <= 2'h0; // @[d_cache.scala 73:19]
    end
    if (reset) begin // @[d_cache.scala 36:31]
      receive_data <= 64'h0; // @[d_cache.scala 36:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          receive_data <= _GEN_5865;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:24]
      quene <= 1'h0; // @[d_cache.scala 37:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          quene <= _GEN_1292;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 76:24]
      state <= 3'h0; // @[d_cache.scala 76:24]
    end else if (3'h0 == state) begin // @[d_cache.scala 81:18]
      if (io_from_lsu_arvalid) begin // @[d_cache.scala 83:38]
        state <= 3'h1; // @[d_cache.scala 84:23]
      end else if (io_from_lsu_awvalid) begin // @[d_cache.scala 85:44]
        state <= 3'h2; // @[d_cache.scala 86:23]
      end
    end else if (3'h1 == state) begin // @[d_cache.scala 81:18]
      if (way0_hit) begin // @[d_cache.scala 91:27]
        state <= _GEN_326;
      end else begin
        state <= _GEN_391;
      end
    end else if (3'h2 == state) begin // @[d_cache.scala 81:18]
      state <= _GEN_1099;
    end else begin
      state <= _GEN_5864;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"read addr : %x  write addr : %x\n",io_from_lsu_araddr,io_from_lsu_awaddr); // @[d_cache.scala 15:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"d_cache state:%d\n",state); // @[d_cache.scala 77:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"receive data:%x\n",receive_data); // @[d_cache.scala 79:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_14 & _T_15 & way0_hit & io_from_lsu_rready & _T_1) begin
          $fwrite(32'h80000002,"dirty_0:%d\n",6'h3f == index ? dirty_0_63 : _GEN_324); // @[d_cache.scala 93:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_8676 & ~way0_hit & way1_hit & io_from_lsu_rready & _T_1) begin
          $fwrite(32'h80000002,"dirty_1:%d\n",6'h3f == index ? dirty_1_63 : _GEN_389); // @[d_cache.scala 99:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"cacheline0:%x   cacheline1:%x\n",_GEN_456,_GEN_712); // @[d_cache.scala 364:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ram_0_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ram_0_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ram_0_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ram_0_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ram_0_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ram_0_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ram_0_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ram_0_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  ram_0_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  ram_0_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  ram_0_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  ram_0_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  ram_0_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  ram_0_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  ram_0_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  ram_0_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  ram_0_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  ram_0_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  ram_0_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  ram_0_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  ram_0_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  ram_0_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  ram_0_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  ram_0_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  ram_0_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  ram_0_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  ram_0_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  ram_0_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  ram_0_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  ram_0_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  ram_0_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  ram_0_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  ram_0_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  ram_0_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  ram_0_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  ram_0_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  ram_0_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  ram_0_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  ram_0_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  ram_0_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  ram_0_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  ram_0_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  ram_0_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  ram_0_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  ram_0_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  ram_0_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  ram_0_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  ram_0_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  ram_0_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  ram_0_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  ram_0_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  ram_0_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  ram_0_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  ram_0_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  ram_0_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  ram_0_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  ram_0_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  ram_0_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  ram_0_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  ram_0_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  ram_0_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  ram_0_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  ram_0_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  ram_0_63 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  ram_1_0 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  ram_1_1 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  ram_1_2 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  ram_1_3 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  ram_1_4 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  ram_1_5 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  ram_1_6 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  ram_1_7 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  ram_1_8 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  ram_1_9 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  ram_1_10 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  ram_1_11 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  ram_1_12 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  ram_1_13 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  ram_1_14 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  ram_1_15 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  ram_1_16 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  ram_1_17 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  ram_1_18 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  ram_1_19 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  ram_1_20 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  ram_1_21 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  ram_1_22 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  ram_1_23 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  ram_1_24 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  ram_1_25 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  ram_1_26 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  ram_1_27 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  ram_1_28 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  ram_1_29 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  ram_1_30 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  ram_1_31 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  ram_1_32 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  ram_1_33 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  ram_1_34 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  ram_1_35 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  ram_1_36 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  ram_1_37 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  ram_1_38 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  ram_1_39 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  ram_1_40 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  ram_1_41 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  ram_1_42 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  ram_1_43 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  ram_1_44 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  ram_1_45 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  ram_1_46 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  ram_1_47 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  ram_1_48 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  ram_1_49 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  ram_1_50 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  ram_1_51 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  ram_1_52 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  ram_1_53 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  ram_1_54 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  ram_1_55 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  ram_1_56 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  ram_1_57 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  ram_1_58 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  ram_1_59 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  ram_1_60 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  ram_1_61 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  ram_1_62 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  ram_1_63 = _RAND_127[63:0];
  _RAND_128 = {1{`RANDOM}};
  tag_0_0 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  tag_0_1 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  tag_0_2 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  tag_0_3 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  tag_0_4 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  tag_0_5 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  tag_0_6 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  tag_0_7 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  tag_0_8 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  tag_0_9 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  tag_0_10 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  tag_0_11 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  tag_0_12 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  tag_0_13 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  tag_0_14 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  tag_0_15 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  tag_0_16 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  tag_0_17 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  tag_0_18 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  tag_0_19 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  tag_0_20 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  tag_0_21 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  tag_0_22 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  tag_0_23 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  tag_0_24 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  tag_0_25 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  tag_0_26 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  tag_0_27 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  tag_0_28 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  tag_0_29 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  tag_0_30 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  tag_0_31 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  tag_0_32 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  tag_0_33 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  tag_0_34 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  tag_0_35 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  tag_0_36 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  tag_0_37 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  tag_0_38 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  tag_0_39 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  tag_0_40 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  tag_0_41 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  tag_0_42 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  tag_0_43 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  tag_0_44 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  tag_0_45 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  tag_0_46 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  tag_0_47 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  tag_0_48 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  tag_0_49 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  tag_0_50 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  tag_0_51 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  tag_0_52 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  tag_0_53 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  tag_0_54 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  tag_0_55 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  tag_0_56 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  tag_0_57 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  tag_0_58 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  tag_0_59 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  tag_0_60 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  tag_0_61 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  tag_0_62 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  tag_0_63 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  tag_1_0 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  tag_1_1 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  tag_1_2 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  tag_1_3 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  tag_1_4 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  tag_1_5 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  tag_1_6 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  tag_1_7 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  tag_1_8 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  tag_1_9 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  tag_1_10 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  tag_1_11 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  tag_1_12 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  tag_1_13 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  tag_1_14 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  tag_1_15 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  tag_1_16 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  tag_1_17 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  tag_1_18 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  tag_1_19 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  tag_1_20 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  tag_1_21 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  tag_1_22 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  tag_1_23 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  tag_1_24 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  tag_1_25 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  tag_1_26 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  tag_1_27 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  tag_1_28 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  tag_1_29 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  tag_1_30 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  tag_1_31 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  tag_1_32 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  tag_1_33 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  tag_1_34 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  tag_1_35 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  tag_1_36 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  tag_1_37 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  tag_1_38 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  tag_1_39 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  tag_1_40 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  tag_1_41 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  tag_1_42 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  tag_1_43 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  tag_1_44 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  tag_1_45 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  tag_1_46 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  tag_1_47 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  tag_1_48 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  tag_1_49 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  tag_1_50 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  tag_1_51 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  tag_1_52 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  tag_1_53 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  tag_1_54 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  tag_1_55 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  tag_1_56 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  tag_1_57 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  tag_1_58 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  tag_1_59 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  tag_1_60 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  tag_1_61 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  tag_1_62 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  tag_1_63 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  valid_0_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_0_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_0_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_0_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_0_4 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_0_5 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_0_6 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_0_7 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_0_8 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_0_9 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_0_10 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_0_11 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_0_12 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_0_13 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_0_14 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_0_15 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_0_16 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_0_17 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_0_18 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_0_19 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_0_20 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_0_21 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_0_22 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_0_23 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_0_24 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_0_25 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_0_26 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_0_27 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_0_28 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_0_29 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_0_30 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_0_31 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_0_32 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_0_33 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_0_34 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_0_35 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_0_36 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_0_37 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_0_38 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_0_39 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_0_40 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_0_41 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_0_42 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_0_43 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_0_44 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_0_45 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_0_46 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_0_47 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_0_48 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_0_49 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_0_50 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_0_51 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_0_52 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_0_53 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_0_54 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_0_55 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_0_56 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_0_57 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_0_58 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_0_59 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_0_60 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_0_61 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_0_62 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_0_63 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_1_0 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_1_1 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_1_2 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_1_3 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_1_4 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_1_5 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_1_6 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_1_7 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_1_8 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_1_9 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_1_10 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_1_11 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_1_12 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_1_13 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_1_14 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_1_15 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_1_16 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_1_17 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_1_18 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_1_19 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_1_20 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_1_21 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_1_22 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_1_23 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_1_24 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_1_25 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_1_26 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_1_27 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_1_28 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_1_29 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_1_30 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_1_31 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_1_32 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_1_33 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_1_34 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_1_35 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_1_36 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_1_37 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_1_38 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_1_39 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_1_40 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_1_41 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_1_42 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_1_43 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_1_44 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_1_45 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_1_46 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_1_47 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_1_48 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_1_49 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_1_50 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_1_51 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_1_52 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_1_53 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_1_54 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_1_55 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_1_56 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_1_57 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_1_58 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_1_59 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_1_60 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_1_61 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_1_62 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_1_63 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  dirty_0_0 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  dirty_0_1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  dirty_0_2 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  dirty_0_3 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  dirty_0_4 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  dirty_0_5 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  dirty_0_6 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  dirty_0_7 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  dirty_0_8 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  dirty_0_9 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  dirty_0_10 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  dirty_0_11 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  dirty_0_12 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  dirty_0_13 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  dirty_0_14 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  dirty_0_15 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  dirty_0_16 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  dirty_0_17 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  dirty_0_18 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  dirty_0_19 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  dirty_0_20 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  dirty_0_21 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  dirty_0_22 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  dirty_0_23 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  dirty_0_24 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  dirty_0_25 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  dirty_0_26 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  dirty_0_27 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  dirty_0_28 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  dirty_0_29 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  dirty_0_30 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  dirty_0_31 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  dirty_0_32 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  dirty_0_33 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  dirty_0_34 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  dirty_0_35 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  dirty_0_36 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  dirty_0_37 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  dirty_0_38 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  dirty_0_39 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  dirty_0_40 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  dirty_0_41 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  dirty_0_42 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  dirty_0_43 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  dirty_0_44 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  dirty_0_45 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  dirty_0_46 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  dirty_0_47 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  dirty_0_48 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  dirty_0_49 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  dirty_0_50 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  dirty_0_51 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  dirty_0_52 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  dirty_0_53 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  dirty_0_54 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  dirty_0_55 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  dirty_0_56 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  dirty_0_57 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  dirty_0_58 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  dirty_0_59 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  dirty_0_60 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  dirty_0_61 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  dirty_0_62 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  dirty_0_63 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  dirty_1_0 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  dirty_1_1 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  dirty_1_2 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  dirty_1_3 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  dirty_1_4 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  dirty_1_5 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  dirty_1_6 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  dirty_1_7 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  dirty_1_8 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  dirty_1_9 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  dirty_1_10 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  dirty_1_11 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  dirty_1_12 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  dirty_1_13 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  dirty_1_14 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  dirty_1_15 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  dirty_1_16 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  dirty_1_17 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  dirty_1_18 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  dirty_1_19 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  dirty_1_20 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  dirty_1_21 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  dirty_1_22 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  dirty_1_23 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  dirty_1_24 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  dirty_1_25 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  dirty_1_26 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  dirty_1_27 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  dirty_1_28 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  dirty_1_29 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  dirty_1_30 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  dirty_1_31 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  dirty_1_32 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  dirty_1_33 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  dirty_1_34 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  dirty_1_35 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  dirty_1_36 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  dirty_1_37 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  dirty_1_38 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  dirty_1_39 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  dirty_1_40 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  dirty_1_41 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  dirty_1_42 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  dirty_1_43 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  dirty_1_44 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  dirty_1_45 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  dirty_1_46 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  dirty_1_47 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  dirty_1_48 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  dirty_1_49 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  dirty_1_50 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  dirty_1_51 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  dirty_1_52 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  dirty_1_53 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  dirty_1_54 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  dirty_1_55 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  dirty_1_56 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  dirty_1_57 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  dirty_1_58 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  dirty_1_59 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  dirty_1_60 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  dirty_1_61 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  dirty_1_62 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  dirty_1_63 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  way0_hit = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  way1_hit = _RAND_513[0:0];
  _RAND_514 = {2{`RANDOM}};
  write_back_data = _RAND_514[63:0];
  _RAND_515 = {1{`RANDOM}};
  write_back_addr = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  unuse_way = _RAND_516[1:0];
  _RAND_517 = {2{`RANDOM}};
  receive_data = _RAND_517[63:0];
  _RAND_518 = {1{`RANDOM}};
  quene = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  state = _RAND_519[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IDU(
  input  [31:0] io_inst,
  output [31:0] io_inst_now,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2,
  output [4:0]  io_rd,
  output [63:0] io_imm,
  output        io_ctrl_sign_reg_write,
  output        io_ctrl_sign_csr_write,
  output        io_ctrl_sign_src2_is_imm,
  output        io_ctrl_sign_src1_is_pc,
  output        io_ctrl_sign_Writemem_en,
  output        io_ctrl_sign_Readmem_en,
  output [7:0]  io_ctrl_sign_Wmask
);
  wire [4:0] rd = io_inst[11:7]; // @[IDU.scala 150:15]
  wire [31:0] _inst_type_T = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_1 = 32'h13 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_2 = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_3 = 32'h17 == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_5 = 32'h37 == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_7 = 32'h6f == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_9 = 32'h67 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_11 = 32'h3023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_13 = 32'h3013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_15 = 32'h2003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_16 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_17 = 32'h3b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_19 = 32'h40000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_21 = 32'h1063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_23 = 32'h63 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_25 = 32'h3003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_27 = 32'h1b == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_29 = 32'h33 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_30 = io_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_31 = 32'h40005013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_33 = 32'h4003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_35 = 32'h1023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_37 = 32'h23 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_39 = 32'h6033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_41 = 32'h4013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_43 = 32'h7033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_45 = 32'h7013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_47 = 32'h4000003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_49 = 32'h103b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_51 = 32'h1013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_53 = 32'h5013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_55 = 32'h101b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_57 = 32'h4000501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_59 = 32'h501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_61 = 32'h4000503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_63 = 32'h503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_65 = 32'h3033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_67 = 32'h2033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_69 = 32'h5063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_71 = 32'h4063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_73 = 32'h6063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_75 = 32'h2023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_77 = 32'h1003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_79 = 32'h5003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_81 = 32'h2000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_83 = 32'h200003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_85 = 32'h200403b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_87 = 32'h200603b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_89 = 32'h4033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_91 = 32'h6013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_93 = 32'h2005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_95 = 32'h2004033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_97 = 32'h200503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_99 = 32'h200703b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_101 = 32'h2007033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_103 = 32'h2006033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_105 = 32'h1033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_107 = 32'h5033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_109 = 32'h40005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_111 = 32'h2013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_113 = 32'h6003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_115 = 32'h3 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_117 = 32'h7063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_119 = 32'h73 == io_inst; // @[Lookup.scala 31:38]
  wire  _inst_type_T_121 = 32'h1073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_123 = 32'h2073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_125 = 32'h3073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [6:0] _inst_type_T_126 = _inst_type_T_125 ? 7'h40 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_127 = _inst_type_T_123 ? 7'h40 : _inst_type_T_126; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_128 = _inst_type_T_121 ? 7'h40 : _inst_type_T_127; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_129 = _inst_type_T_119 ? 7'h40 : _inst_type_T_128; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_130 = _inst_type_T_117 ? 7'h45 : _inst_type_T_129; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_131 = _inst_type_T_115 ? 7'h40 : _inst_type_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_132 = _inst_type_T_113 ? 7'h40 : _inst_type_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_133 = _inst_type_T_111 ? 7'h40 : _inst_type_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_134 = _inst_type_T_109 ? 7'h41 : _inst_type_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_135 = _inst_type_T_107 ? 7'h41 : _inst_type_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_136 = _inst_type_T_105 ? 7'h41 : _inst_type_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_137 = _inst_type_T_103 ? 7'h41 : _inst_type_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_138 = _inst_type_T_101 ? 7'h41 : _inst_type_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_139 = _inst_type_T_99 ? 7'h41 : _inst_type_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_140 = _inst_type_T_97 ? 7'h41 : _inst_type_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_141 = _inst_type_T_95 ? 7'h41 : _inst_type_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_142 = _inst_type_T_93 ? 7'h41 : _inst_type_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_143 = _inst_type_T_91 ? 7'h40 : _inst_type_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_144 = _inst_type_T_89 ? 7'h41 : _inst_type_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_145 = _inst_type_T_87 ? 7'h41 : _inst_type_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_146 = _inst_type_T_85 ? 7'h41 : _inst_type_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_147 = _inst_type_T_83 ? 7'h41 : _inst_type_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_148 = _inst_type_T_81 ? 7'h41 : _inst_type_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_149 = _inst_type_T_79 ? 7'h40 : _inst_type_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_150 = _inst_type_T_77 ? 7'h40 : _inst_type_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_151 = _inst_type_T_75 ? 7'h44 : _inst_type_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_152 = _inst_type_T_73 ? 7'h45 : _inst_type_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_153 = _inst_type_T_71 ? 7'h45 : _inst_type_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_154 = _inst_type_T_69 ? 7'h45 : _inst_type_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_155 = _inst_type_T_67 ? 7'h41 : _inst_type_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_156 = _inst_type_T_65 ? 7'h41 : _inst_type_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_157 = _inst_type_T_63 ? 7'h41 : _inst_type_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_158 = _inst_type_T_61 ? 7'h41 : _inst_type_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_159 = _inst_type_T_59 ? 7'h40 : _inst_type_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_160 = _inst_type_T_57 ? 7'h40 : _inst_type_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_161 = _inst_type_T_55 ? 7'h40 : _inst_type_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_162 = _inst_type_T_53 ? 7'h40 : _inst_type_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_163 = _inst_type_T_51 ? 7'h40 : _inst_type_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_164 = _inst_type_T_49 ? 7'h41 : _inst_type_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_165 = _inst_type_T_47 ? 7'h41 : _inst_type_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_166 = _inst_type_T_45 ? 7'h40 : _inst_type_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_167 = _inst_type_T_43 ? 7'h41 : _inst_type_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_168 = _inst_type_T_41 ? 7'h40 : _inst_type_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_169 = _inst_type_T_39 ? 7'h41 : _inst_type_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_170 = _inst_type_T_37 ? 7'h44 : _inst_type_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_171 = _inst_type_T_35 ? 7'h44 : _inst_type_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_172 = _inst_type_T_33 ? 7'h40 : _inst_type_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_173 = _inst_type_T_31 ? 7'h40 : _inst_type_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_174 = _inst_type_T_29 ? 7'h41 : _inst_type_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_175 = _inst_type_T_27 ? 7'h40 : _inst_type_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_176 = _inst_type_T_25 ? 7'h40 : _inst_type_T_175; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_177 = _inst_type_T_23 ? 7'h45 : _inst_type_T_176; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_178 = _inst_type_T_21 ? 7'h45 : _inst_type_T_177; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_179 = _inst_type_T_19 ? 7'h41 : _inst_type_T_178; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_180 = _inst_type_T_17 ? 7'h41 : _inst_type_T_179; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_181 = _inst_type_T_15 ? 7'h40 : _inst_type_T_180; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_182 = _inst_type_T_13 ? 7'h40 : _inst_type_T_181; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_183 = _inst_type_T_11 ? 7'h44 : _inst_type_T_182; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_184 = _inst_type_T_9 ? 7'h40 : _inst_type_T_183; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_185 = _inst_type_T_7 ? 7'h43 : _inst_type_T_184; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_186 = _inst_type_T_5 ? 7'h42 : _inst_type_T_185; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_187 = _inst_type_T_3 ? 7'h42 : _inst_type_T_186; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_188 = _inst_type_T_1 ? 7'h40 : _inst_type_T_187; // @[Lookup.scala 34:39]
  wire [11:0] imm_imm = io_inst[31:20]; // @[IDU.scala 24:23]
  wire [51:0] _imm_T_2 = imm_imm[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_3 = {_imm_T_2,imm_imm}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_1 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21]}; // @[Cat.scala 31:58]
  wire [42:0] _imm_T_6 = imm_imm_1[19] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_7 = {_imm_T_6,io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_2 = io_inst[31:12]; // @[IDU.scala 28:23]
  wire [31:0] _imm_T_10 = imm_imm_2[19] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_12 = {_imm_T_10,imm_imm_2,12'h0}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_3 = {io_inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [51:0] _imm_T_15 = imm_imm_3[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_16 = {_imm_T_15,io_inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_4 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8]}; // @[Cat.scala 31:58]
  wire [50:0] _imm_T_19 = imm_imm_4[11] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_20 = {_imm_T_19,io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] inst_type = {{25'd0}, _inst_type_T_188}; // @[IDU.scala 133:25 152:15]
  wire [63:0] _imm_T_22 = 32'h40 == inst_type ? _imm_T_3 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_24 = 32'h43 == inst_type ? _imm_T_7 : _imm_T_22; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_26 = 32'h42 == inst_type ? _imm_T_12 : _imm_T_24; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_28 = 32'h44 == inst_type ? _imm_T_16 : _imm_T_26; // @[Mux.scala 81:58]
  wire  _inst_now_T_3 = 32'h100073 == io_inst; // @[Lookup.scala 31:38]
  wire  _inst_now_T_123 = 32'h30200073 == io_inst; // @[Lookup.scala 31:38]
  wire [6:0] _inst_now_T_130 = _inst_type_T_125 ? 7'h47 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_131 = _inst_type_T_123 ? 7'h46 : _inst_now_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_132 = _inst_type_T_121 ? 7'h3f : _inst_now_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_133 = _inst_now_T_123 ? 7'h3e : _inst_now_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_134 = _inst_type_T_119 ? 7'h3d : _inst_now_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_135 = _inst_type_T_117 ? 7'h3c : _inst_now_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_136 = _inst_type_T_115 ? 7'h3b : _inst_now_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_137 = _inst_type_T_113 ? 7'h3a : _inst_now_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_138 = _inst_type_T_111 ? 7'h36 : _inst_now_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_139 = _inst_type_T_109 ? 7'h39 : _inst_now_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_140 = _inst_type_T_107 ? 7'h38 : _inst_now_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_141 = _inst_type_T_105 ? 7'h37 : _inst_now_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_142 = _inst_type_T_103 ? 7'h34 : _inst_now_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_143 = _inst_type_T_101 ? 7'h33 : _inst_now_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_144 = _inst_type_T_99 ? 7'h32 : _inst_now_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_145 = _inst_type_T_97 ? 7'h35 : _inst_now_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_146 = _inst_type_T_95 ? 7'h31 : _inst_now_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_147 = _inst_type_T_93 ? 7'h30 : _inst_now_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_148 = _inst_type_T_91 ? 7'h2f : _inst_now_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_149 = _inst_type_T_89 ? 7'h2e : _inst_now_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_150 = _inst_type_T_87 ? 7'h14 : _inst_now_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_151 = _inst_type_T_85 ? 7'h13 : _inst_now_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_152 = _inst_type_T_83 ? 7'h12 : _inst_now_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_153 = _inst_type_T_81 ? 7'h11 : _inst_now_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_154 = _inst_type_T_79 ? 7'h25 : _inst_now_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_155 = _inst_type_T_77 ? 7'h24 : _inst_now_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_156 = _inst_type_T_75 ? 7'h27 : _inst_now_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_157 = _inst_type_T_73 ? 7'h2d : _inst_now_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_158 = _inst_type_T_71 ? 7'h2c : _inst_now_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_159 = _inst_type_T_69 ? 7'h2b : _inst_now_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_160 = _inst_type_T_67 ? 7'h1f : _inst_now_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_161 = _inst_type_T_65 ? 7'h1e : _inst_now_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_162 = _inst_type_T_63 ? 7'h1d : _inst_now_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_163 = _inst_type_T_61 ? 7'h1c : _inst_now_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_164 = _inst_type_T_59 ? 7'h1b : _inst_now_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_165 = _inst_type_T_57 ? 7'h1a : _inst_now_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_166 = _inst_type_T_55 ? 7'h19 : _inst_now_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_167 = _inst_type_T_53 ? 7'h18 : _inst_now_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_168 = _inst_type_T_51 ? 7'h17 : _inst_now_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_169 = _inst_type_T_49 ? 7'h16 : _inst_now_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_170 = _inst_type_T_47 ? 7'hd : _inst_now_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_171 = _inst_type_T_45 ? 7'h9 : _inst_now_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_172 = _inst_type_T_43 ? 7'h8 : _inst_now_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_173 = _inst_type_T_41 ? 7'ha : _inst_now_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_174 = _inst_type_T_39 ? 7'hb : _inst_now_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_175 = _inst_type_T_37 ? 7'h28 : _inst_now_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_176 = _inst_type_T_35 ? 7'h26 : _inst_now_T_175; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_177 = _inst_type_T_33 ? 7'h23 : _inst_now_T_176; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_178 = _inst_type_T_31 ? 7'h15 : _inst_now_T_177; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_179 = _inst_type_T_29 ? 7'hf : _inst_now_T_178; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_180 = _inst_type_T_27 ? 7'h10 : _inst_now_T_179; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_181 = _inst_type_T_25 ? 7'h22 : _inst_now_T_180; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_182 = _inst_type_T_23 ? 7'h29 : _inst_now_T_181; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_183 = _inst_type_T_21 ? 7'h2a : _inst_now_T_182; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_184 = _inst_type_T_19 ? 7'he : _inst_now_T_183; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_185 = _inst_type_T_17 ? 7'hc : _inst_now_T_184; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_186 = _inst_type_T_15 ? 7'h21 : _inst_now_T_185; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_187 = _inst_type_T_13 ? 7'h20 : _inst_now_T_186; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_188 = _inst_type_T_11 ? 7'h7 : _inst_now_T_187; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_189 = _inst_type_T_9 ? 7'h6 : _inst_now_T_188; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_190 = _inst_type_T_7 ? 7'h5 : _inst_now_T_189; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_191 = _inst_type_T_5 ? 7'h4 : _inst_now_T_190; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_192 = _inst_type_T_3 ? 7'h3 : _inst_now_T_191; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_193 = _inst_now_T_3 ? 7'h2 : _inst_now_T_192; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_194 = _inst_type_T_1 ? 7'h1 : _inst_now_T_193; // @[Lookup.scala 34:39]
  wire  _reg_write_T_26 = _inst_now_T_123 ? 1'h0 : 1'h1; // @[Lookup.scala 34:39]
  wire  _reg_write_T_27 = _inst_type_T_119 ? 1'h0 : _reg_write_T_26; // @[Lookup.scala 34:39]
  wire  _reg_write_T_28 = _inst_type_T_117 ? 1'h0 : _reg_write_T_27; // @[Lookup.scala 34:39]
  wire  _reg_write_T_29 = _inst_type_T_73 ? 1'h0 : _reg_write_T_28; // @[Lookup.scala 34:39]
  wire  _reg_write_T_30 = _inst_type_T_71 ? 1'h0 : _reg_write_T_29; // @[Lookup.scala 34:39]
  wire  _reg_write_T_31 = _inst_type_T_69 ? 1'h0 : _reg_write_T_30; // @[Lookup.scala 34:39]
  wire  _reg_write_T_32 = _inst_type_T_23 ? 1'h0 : _reg_write_T_31; // @[Lookup.scala 34:39]
  wire  _reg_write_T_33 = _inst_type_T_21 ? 1'h0 : _reg_write_T_32; // @[Lookup.scala 34:39]
  wire  _reg_write_T_34 = _inst_type_T_75 ? 1'h0 : _reg_write_T_33; // @[Lookup.scala 34:39]
  wire  _reg_write_T_35 = _inst_type_T_37 ? 1'h0 : _reg_write_T_34; // @[Lookup.scala 34:39]
  wire  _reg_write_T_36 = _inst_type_T_35 ? 1'h0 : _reg_write_T_35; // @[Lookup.scala 34:39]
  wire  _reg_write_T_37 = _inst_type_T_11 ? 1'h0 : _reg_write_T_36; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_8 = _inst_type_T_75 ? 4'hf : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_9 = _inst_type_T_37 ? 4'h1 : _Wmask_T_8; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_10 = _inst_type_T_35 ? 4'h3 : _Wmask_T_9; // @[Lookup.scala 34:39]
  assign io_inst_now = {{25'd0}, _inst_now_T_194}; // @[IDU.scala 132:24 226:14]
  assign io_rs1 = io_inst[19:15]; // @[IDU.scala 149:16]
  assign io_rs2 = io_inst[24:20]; // @[IDU.scala 148:16]
  assign io_rd = io_inst[11:7]; // @[IDU.scala 150:15]
  assign io_imm = 32'h45 == inst_type ? _imm_T_20 : _imm_T_28; // @[Mux.scala 81:58]
  assign io_ctrl_sign_reg_write = _inst_now_T_3 ? 1'h0 : _reg_write_T_37; // @[Lookup.scala 34:39]
  assign io_ctrl_sign_csr_write = _inst_type_T_121 | (_inst_type_T_123 | _inst_type_T_125); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_src2_is_imm = 32'h45 == inst_type | (32'h43 == inst_type | (32'h44 == inst_type | (32'h42 ==
    inst_type | 32'h40 == inst_type))); // @[Mux.scala 81:58]
  assign io_ctrl_sign_src1_is_pc = _inst_type_T_7 | (_inst_type_T_3 | (_inst_type_T_21 | (_inst_type_T_23 | (
    _inst_type_T_69 | (_inst_type_T_71 | (_inst_type_T_73 | _inst_type_T_117)))))); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Writemem_en = 32'h44 == inst_type; // @[Mux.scala 81:61]
  assign io_ctrl_sign_Readmem_en = _inst_type_T_25 | (_inst_type_T_15 | (_inst_type_T_113 | (_inst_type_T_77 | (
    _inst_type_T_79 | (_inst_type_T_115 | _inst_type_T_33))))); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Wmask = _inst_type_T_11 ? 8'hff : {{4'd0}, _Wmask_T_10}; // @[Lookup.scala 34:39]
endmodule
module EXU_AXI(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  output [63:0] io_pc_next,
  input  [31:0] io_inst_now,
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [4:0]  io_rd,
  input  [63:0] io_imm,
  input         io_ctrl_sign_reg_write,
  input         io_ctrl_sign_csr_write,
  input         io_ctrl_sign_src2_is_imm,
  input         io_ctrl_sign_src1_is_pc,
  input         io_ctrl_sign_Writemem_en,
  input         io_ctrl_sign_Readmem_en,
  input  [7:0]  io_ctrl_sign_Wmask,
  output [63:0] io_res2rd,
  input         io_inst_valid,
  output        io_inst_store,
  output        io_inst_load,
  output [31:0] io_Mem_addr,
  input  [63:0] io_Mem_rdata,
  output [63:0] io_Mem_wdata,
  output [7:0]  io_Mem_wstrb,
  input         io_rdata_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] Regfile [0:31]; // @[EXU_AXI.scala 37:22]
  wire  Regfile_src1_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_src1_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_src1_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_src2_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_src2_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_src2_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_4_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_MPORT_4_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_MPORT_4_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_1_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_1_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_1_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_2_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_2_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_2_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_3_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_3_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_3_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_4_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_4_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_4_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_5_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_5_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_5_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_6_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_6_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_6_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_7_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_7_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_7_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_8_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_8_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_8_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_9_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_9_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_9_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_10_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_10_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_10_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_11_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_11_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_11_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_0_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_0_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_0_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_1_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_1_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_1_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_2_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_2_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_2_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_3_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_3_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_3_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_4_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_4_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_4_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_5_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_5_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_5_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_6_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_6_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_6_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_7_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_7_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_7_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_8_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_8_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_8_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_9_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_9_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_9_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_10_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_10_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_10_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_11_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_11_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_11_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_12_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_12_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_12_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_13_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_13_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_13_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_14_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_14_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_14_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_15_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_15_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_15_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_16_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_16_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_16_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_17_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_17_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_17_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_18_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_18_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_18_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_19_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_19_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_19_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_20_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_20_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_20_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_21_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_21_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_21_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_22_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_22_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_22_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_23_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_23_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_23_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_24_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_24_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_24_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_25_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_25_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_25_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_26_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_26_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_26_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_27_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_27_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_27_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_28_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_28_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_28_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_29_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_29_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_29_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_30_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_30_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_30_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_31_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_31_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_31_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_1_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_1_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_1_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_2_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_2_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_2_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_3_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_3_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_3_data; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_mask; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_en; // @[EXU_AXI.scala 37:22]
  reg [63:0] CSR_Reg [0:3]; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_2_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_2_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_2_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_csr_wdata_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_csr_wdata_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_csr_wdata_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_csr_wdata_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_csr_wdata_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_csr_wdata_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_2_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_2_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_2_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_5_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_5_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_5_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_7_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_7_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_7_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_j_pc_MPORT_12_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_j_pc_MPORT_12_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_j_pc_MPORT_12_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_j_pc_MPORT_13_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_j_pc_MPORT_13_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_j_pc_MPORT_13_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_0_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_1_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_2_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_1_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_3_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_3_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_3_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_3_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_6_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_6_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_6_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_6_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] reg_trace_input_reg_0; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_1; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_2; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_3; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_4; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_5; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_6; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_7; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_8; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_9; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_10; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_11; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_12; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_13; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_14; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_15; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_16; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_17; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_18; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_19; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_20; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_21; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_22; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_23; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_24; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_25; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_26; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_27; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_28; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_29; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_30; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_31; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_0; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_1; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_2; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_3; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_pc; // @[EXU_AXI.scala 163:27]
  wire [11:0] csr_addr = io_imm[11:0]; // @[EXU_AXI.scala 39:26]
  wire [1:0] _csr_index_T_5 = 12'h300 == csr_addr ? 2'h2 : {{1'd0}, 12'h341 == csr_addr}; // @[Mux.scala 81:58]
  wire  _csr_index_T_6 = 12'h342 == csr_addr; // @[Mux.scala 81:61]
  wire [63:0] _src1_value_T_1 = io_rs1 == 5'h0 ? 64'h0 : Regfile_src1_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] src1_value = io_ctrl_sign_src1_is_pc ? io_pc : _src1_value_T_1; // @[EXU_AXI.scala 49:25]
  wire [63:0] _src2_value_T_1 = io_rs2 == 5'h0 ? 64'h0 : Regfile_src2_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] src2_value = io_ctrl_sign_src2_is_imm ? io_imm : _src2_value_T_1; // @[EXU_AXI.scala 50:25]
  wire [63:0] add_res = src1_value + src2_value; // @[EXU_AXI.scala 51:30]
  wire [63:0] sub_res = src1_value - src2_value; // @[EXU_AXI.scala 52:30]
  wire [63:0] _sra_res_T = io_ctrl_sign_src1_is_pc ? io_pc : _src1_value_T_1; // @[EXU_AXI.scala 53:37]
  wire [63:0] sra_res = $signed(_sra_res_T) >>> src2_value[5:0]; // @[EXU_AXI.scala 53:60]
  wire [63:0] srl_res = src1_value >> src2_value[5:0]; // @[EXU_AXI.scala 54:30]
  wire [126:0] _GEN_1 = {{63'd0}, src1_value}; // @[EXU_AXI.scala 55:30]
  wire [126:0] sll_res = _GEN_1 << src2_value[5:0]; // @[EXU_AXI.scala 55:30]
  wire [31:0] _sraw_res_T_1 = src1_value[31:0]; // @[EXU_AXI.scala 56:43]
  wire [31:0] sraw_res = $signed(_sraw_res_T_1) >>> src2_value[4:0]; // @[EXU_AXI.scala 56:46]
  wire [31:0] srlw_res = src1_value[31:0] >> src2_value[4:0]; // @[EXU_AXI.scala 57:37]
  wire [62:0] _GEN_2 = {{31'd0}, src1_value[31:0]}; // @[EXU_AXI.scala 58:37]
  wire [62:0] sllw_res = _GEN_2 << src2_value[4:0]; // @[EXU_AXI.scala 58:37]
  wire [63:0] or_res = src1_value | src2_value; // @[EXU_AXI.scala 59:29]
  wire [63:0] xor_res = src1_value ^ src2_value; // @[EXU_AXI.scala 60:30]
  wire [63:0] and_res = src1_value & src2_value; // @[EXU_AXI.scala 61:30]
  wire [127:0] _mlu_res_T = src1_value * src2_value; // @[EXU_AXI.scala 62:31]
  wire [63:0] mlu_res = _mlu_res_T[63:0]; // @[EXU_AXI.scala 62:44]
  wire [63:0] _mluw_res_T_2 = src1_value[31:0] * src2_value[31:0]; // @[EXU_AXI.scala 63:38]
  wire [31:0] mluw_res = _mluw_res_T_2[31:0]; // @[EXU_AXI.scala 63:57]
  wire [31:0] _divw_res_T_3 = src2_value[31:0]; // @[EXU_AXI.scala 64:64]
  wire [32:0] _divw_res_T_4 = $signed(_sraw_res_T_1) / $signed(_divw_res_T_3); // @[EXU_AXI.scala 64:45]
  wire [31:0] divw_res = _divw_res_T_4[31:0]; // @[EXU_AXI.scala 64:71]
  wire [31:0] divuw_res = src1_value[31:0] / src2_value[31:0]; // @[EXU_AXI.scala 65:39]
  wire [31:0] remw_res = $signed(_sraw_res_T_1) % $signed(_divw_res_T_3); // @[EXU_AXI.scala 66:71]
  wire [31:0] remuw_res = src1_value[31:0] % src2_value[31:0]; // @[EXU_AXI.scala 67:39]
  wire [63:0] _div_res_T_1 = io_ctrl_sign_src2_is_imm ? io_imm : _src2_value_T_1; // @[EXU_AXI.scala 68:51]
  wire [64:0] div_res = $signed(_sra_res_T) / $signed(_div_res_T_1); // @[EXU_AXI.scala 68:59]
  wire [63:0] divu_res = src1_value / src2_value; // @[EXU_AXI.scala 69:31]
  wire [63:0] rem_res = $signed(_sra_res_T) % $signed(_div_res_T_1); // @[EXU_AXI.scala 70:59]
  wire [63:0] remu_res = src1_value % src2_value; // @[EXU_AXI.scala 71:31]
  wire [63:0] _io_res2rd_T_1 = io_pc + 64'h4; // @[EXU_AXI.scala 76:24]
  wire  _io_res2rd_T_4 = src1_value < src2_value; // @[EXU_AXI.scala 78:34]
  wire  _io_res2rd_T_10 = $signed(_sra_res_T) < $signed(_div_res_T_1); // @[EXU_AXI.scala 80:42]
  wire [31:0] _io_res2rd_T_18 = io_Mem_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_20 = {_io_res2rd_T_18,io_Mem_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_23 = {56'h0,io_Mem_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_26 = {32'h0,io_Mem_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [47:0] _io_res2rd_T_29 = io_Mem_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_31 = {_io_res2rd_T_29,io_Mem_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [55:0] _io_res2rd_T_34 = io_Mem_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_36 = {_io_res2rd_T_34,io_Mem_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_39 = {48'h0,io_Mem_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_42 = add_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_44 = {_io_res2rd_T_42,add_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_52 = sub_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_54 = {_io_res2rd_T_52,sub_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_57 = sllw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_59 = {_io_res2rd_T_57,sllw_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_67 = sraw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _io_res2rd_T_68 = $signed(_sraw_res_T_1) >>> src2_value[4:0]; // @[EXU_AXI.scala 105:56]
  wire [63:0] _io_res2rd_T_69 = {_io_res2rd_T_67,_io_res2rd_T_68}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_72 = srlw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_74 = {_io_res2rd_T_72,srlw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_87 = mluw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_88 = {_io_res2rd_T_87,mluw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_91 = divw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_92 = {_io_res2rd_T_91,divw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_95 = divuw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_96 = {_io_res2rd_T_95,divuw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_99 = remw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_100 = {_io_res2rd_T_99,remw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_103 = remuw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_104 = {_io_res2rd_T_103,remuw_res}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_106 = 32'h1 == io_inst_now ? add_res : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_108 = 32'h3 == io_inst_now ? add_res : _io_res2rd_T_106; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_110 = 32'h4 == io_inst_now ? io_imm : _io_res2rd_T_108; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_112 = 32'h5 == io_inst_now ? _io_res2rd_T_1 : _io_res2rd_T_110; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_114 = 32'h6 == io_inst_now ? _io_res2rd_T_1 : _io_res2rd_T_112; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_116 = 32'h20 == io_inst_now ? {{63'd0}, _io_res2rd_T_4} : _io_res2rd_T_114; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_118 = 32'h1e == io_inst_now ? {{63'd0}, _io_res2rd_T_4} : _io_res2rd_T_116; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_120 = 32'h36 == io_inst_now ? {{63'd0}, _io_res2rd_T_10} : _io_res2rd_T_118; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_122 = 32'h1f == io_inst_now ? {{63'd0}, _io_res2rd_T_10} : _io_res2rd_T_120; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_124 = 32'h21 == io_inst_now ? _io_res2rd_T_20 : _io_res2rd_T_122; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_126 = 32'h22 == io_inst_now ? io_Mem_rdata : _io_res2rd_T_124; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_128 = 32'h23 == io_inst_now ? _io_res2rd_T_23 : _io_res2rd_T_126; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_130 = 32'h3a == io_inst_now ? _io_res2rd_T_26 : _io_res2rd_T_128; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_132 = 32'h24 == io_inst_now ? _io_res2rd_T_31 : _io_res2rd_T_130; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_134 = 32'h3b == io_inst_now ? _io_res2rd_T_36 : _io_res2rd_T_132; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_136 = 32'h25 == io_inst_now ? _io_res2rd_T_39 : _io_res2rd_T_134; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_138 = 32'hc == io_inst_now ? _io_res2rd_T_44 : _io_res2rd_T_136; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_140 = 32'he == io_inst_now ? sub_res : _io_res2rd_T_138; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_142 = 32'h10 == io_inst_now ? _io_res2rd_T_44 : _io_res2rd_T_140; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_144 = 32'hf == io_inst_now ? add_res : _io_res2rd_T_142; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_146 = 32'h15 == io_inst_now ? sra_res : _io_res2rd_T_144; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_148 = 32'hb == io_inst_now ? or_res : _io_res2rd_T_146; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_150 = 32'h2f == io_inst_now ? or_res : _io_res2rd_T_148; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_152 = 32'h2e == io_inst_now ? xor_res : _io_res2rd_T_150; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_154 = 32'ha == io_inst_now ? xor_res : _io_res2rd_T_152; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_156 = 32'h8 == io_inst_now ? and_res : _io_res2rd_T_154; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_158 = 32'h9 == io_inst_now ? and_res : _io_res2rd_T_156; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_160 = 32'hd == io_inst_now ? _io_res2rd_T_54 : _io_res2rd_T_158; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_162 = 32'h16 == io_inst_now ? _io_res2rd_T_59 : _io_res2rd_T_160; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_164 = 32'h17 == io_inst_now ? sll_res : {{63'd0}, _io_res2rd_T_162}; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_166 = 32'h18 == io_inst_now ? {{63'd0}, srl_res} : _io_res2rd_T_164; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_168 = 32'h19 == io_inst_now ? {{63'd0}, _io_res2rd_T_59} : _io_res2rd_T_166; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_170 = 32'h1a == io_inst_now ? {{63'd0}, _io_res2rd_T_69} : _io_res2rd_T_168; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_172 = 32'h1b == io_inst_now ? {{63'd0}, _io_res2rd_T_74} : _io_res2rd_T_170; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_174 = 32'h1c == io_inst_now ? {{63'd0}, _io_res2rd_T_69} : _io_res2rd_T_172; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_176 = 32'h1d == io_inst_now ? {{63'd0}, _io_res2rd_T_74} : _io_res2rd_T_174; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_178 = 32'h11 == io_inst_now ? {{63'd0}, mlu_res} : _io_res2rd_T_176; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_180 = 32'h12 == io_inst_now ? {{63'd0}, _io_res2rd_T_88} : _io_res2rd_T_178; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_182 = 32'h13 == io_inst_now ? {{63'd0}, _io_res2rd_T_92} : _io_res2rd_T_180; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_184 = 32'h30 == io_inst_now ? {{63'd0}, divu_res} : _io_res2rd_T_182; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_186 = 32'h31 == io_inst_now ? {{62'd0}, div_res} : _io_res2rd_T_184; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_188 = 32'h35 == io_inst_now ? {{63'd0}, _io_res2rd_T_96} : _io_res2rd_T_186; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_190 = 32'h14 == io_inst_now ? {{63'd0}, _io_res2rd_T_100} : _io_res2rd_T_188; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_192 = 32'h32 == io_inst_now ? {{63'd0}, _io_res2rd_T_104} : _io_res2rd_T_190; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_194 = 32'h33 == io_inst_now ? {{63'd0}, remu_res} : _io_res2rd_T_192; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_196 = 32'h34 == io_inst_now ? {{63'd0}, rem_res} : _io_res2rd_T_194; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_198 = 32'h37 == io_inst_now ? sll_res : _io_res2rd_T_196; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_200 = 32'h39 == io_inst_now ? {{63'd0}, sra_res} : _io_res2rd_T_198; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_202 = 32'h38 == io_inst_now ? {{63'd0}, srl_res} : _io_res2rd_T_200; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_204 = 32'h3f == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_data} : _io_res2rd_T_202; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_206 = 32'h46 == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_1_data} : _io_res2rd_T_204; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_208 = 32'h47 == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_2_data} : _io_res2rd_T_206; // @[Mux.scala 81:58]
  wire [63:0] reg_value = io_rd == 5'h0 ? 64'h0 : Regfile_reg_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire  _T_6 = io_ctrl_sign_reg_write & io_rd != 5'h0 & (io_inst_valid & ~io_ctrl_sign_Readmem_en |
    io_ctrl_sign_Readmem_en & io_rdata_valid); // @[EXU_AXI.scala 129:63]
  wire [63:0] _csr_wdata_T = src1_value | CSR_Reg_csr_wdata_MPORT_data; // @[EXU_AXI.scala 134:32]
  wire [63:0] _csr_wdata_T_1 = ~CSR_Reg_csr_wdata_MPORT_1_data; // @[EXU_AXI.scala 135:35]
  wire [63:0] _csr_wdata_T_2 = src1_value & _csr_wdata_T_1; // @[EXU_AXI.scala 135:32]
  wire [63:0] _csr_wdata_T_4 = 32'h3f == io_inst_now ? src1_value : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _csr_wdata_T_6 = 32'h46 == io_inst_now ? _csr_wdata_T : _csr_wdata_T_4; // @[Mux.scala 81:58]
  wire [63:0] csr_wdata = 32'h47 == io_inst_now ? _csr_wdata_T_2 : _csr_wdata_T_6; // @[Mux.scala 81:58]
  wire  _T_9 = io_inst_now == 32'h3d & io_inst_valid; // @[EXU_AXI.scala 138:48]
  wire  _T_14 = io_ctrl_sign_csr_write & io_inst_valid; // @[EXU_AXI.scala 141:53]
  wire [63:0] _j_pc_T = add_res & 64'hfffffffffffffffe; // @[EXU_AXI.scala 148:28]
  wire [63:0] _j_pc_T_3 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_data; // @[EXU_AXI.scala 149:39]
  wire [63:0] _j_pc_T_6 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_1_data; // @[EXU_AXI.scala 149:67]
  wire [63:0] _j_pc_T_8 = $signed(_j_pc_T_3) != $signed(_j_pc_T_6) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 149:21]
  wire [63:0] _j_pc_T_11 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_2_data; // @[EXU_AXI.scala 150:39]
  wire [63:0] _j_pc_T_14 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_3_data; // @[EXU_AXI.scala 150:67]
  wire [63:0] _j_pc_T_16 = $signed(_j_pc_T_11) == $signed(_j_pc_T_14) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 150:21]
  wire [63:0] _j_pc_T_19 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_4_data; // @[EXU_AXI.scala 151:39]
  wire [63:0] _j_pc_T_22 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_5_data; // @[EXU_AXI.scala 151:66]
  wire [63:0] _j_pc_T_24 = $signed(_j_pc_T_19) >= $signed(_j_pc_T_22) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 151:21]
  wire [63:0] _j_pc_T_27 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_6_data; // @[EXU_AXI.scala 152:39]
  wire [63:0] _j_pc_T_30 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_7_data; // @[EXU_AXI.scala 152:65]
  wire [63:0] _j_pc_T_32 = $signed(_j_pc_T_27) < $signed(_j_pc_T_30) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 152:21]
  wire [63:0] _j_pc_T_34 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_8_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_36 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_9_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_38 = _j_pc_T_34 < _j_pc_T_36 ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 153:22]
  wire [63:0] _j_pc_T_40 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_10_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_42 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_11_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_44 = _j_pc_T_40 >= _j_pc_T_42 ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 154:22]
  wire [63:0] _j_pc_T_46 = CSR_Reg_j_pc_MPORT_13_data + 64'h4; // @[EXU_AXI.scala 156:33]
  wire [63:0] _j_pc_T_48 = 32'h5 == io_inst_now ? add_res : _io_res2rd_T_1; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_50 = 32'h6 == io_inst_now ? _j_pc_T : _j_pc_T_48; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_52 = 32'h2a == io_inst_now ? _j_pc_T_8 : _j_pc_T_50; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_54 = 32'h29 == io_inst_now ? _j_pc_T_16 : _j_pc_T_52; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_56 = 32'h2b == io_inst_now ? _j_pc_T_24 : _j_pc_T_54; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_58 = 32'h2c == io_inst_now ? _j_pc_T_32 : _j_pc_T_56; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_60 = 32'h2d == io_inst_now ? _j_pc_T_38 : _j_pc_T_58; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_62 = 32'h3c == io_inst_now ? _j_pc_T_44 : _j_pc_T_60; // @[Mux.scala 81:58]
  reg [63:0] pc_next; // @[EXU_AXI.scala 158:26]
  wire [63:0] _mem_wdata_T_1 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_3 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_1_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_6 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_2_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_9 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_3_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_12 = 32'h7 == io_inst_now ? _mem_wdata_T_1 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _mem_wdata_T_14 = 32'h26 == io_inst_now ? {{48'd0}, _mem_wdata_T_3[15:0]} : _mem_wdata_T_12; // @[Mux.scala 81:58]
  wire [63:0] _mem_wdata_T_16 = 32'h28 == io_inst_now ? {{56'd0}, _mem_wdata_T_6[7:0]} : _mem_wdata_T_14; // @[Mux.scala 81:58]
  traceregs reg_trace ( // @[EXU_AXI.scala 163:27]
    .input_reg_0(reg_trace_input_reg_0),
    .input_reg_1(reg_trace_input_reg_1),
    .input_reg_2(reg_trace_input_reg_2),
    .input_reg_3(reg_trace_input_reg_3),
    .input_reg_4(reg_trace_input_reg_4),
    .input_reg_5(reg_trace_input_reg_5),
    .input_reg_6(reg_trace_input_reg_6),
    .input_reg_7(reg_trace_input_reg_7),
    .input_reg_8(reg_trace_input_reg_8),
    .input_reg_9(reg_trace_input_reg_9),
    .input_reg_10(reg_trace_input_reg_10),
    .input_reg_11(reg_trace_input_reg_11),
    .input_reg_12(reg_trace_input_reg_12),
    .input_reg_13(reg_trace_input_reg_13),
    .input_reg_14(reg_trace_input_reg_14),
    .input_reg_15(reg_trace_input_reg_15),
    .input_reg_16(reg_trace_input_reg_16),
    .input_reg_17(reg_trace_input_reg_17),
    .input_reg_18(reg_trace_input_reg_18),
    .input_reg_19(reg_trace_input_reg_19),
    .input_reg_20(reg_trace_input_reg_20),
    .input_reg_21(reg_trace_input_reg_21),
    .input_reg_22(reg_trace_input_reg_22),
    .input_reg_23(reg_trace_input_reg_23),
    .input_reg_24(reg_trace_input_reg_24),
    .input_reg_25(reg_trace_input_reg_25),
    .input_reg_26(reg_trace_input_reg_26),
    .input_reg_27(reg_trace_input_reg_27),
    .input_reg_28(reg_trace_input_reg_28),
    .input_reg_29(reg_trace_input_reg_29),
    .input_reg_30(reg_trace_input_reg_30),
    .input_reg_31(reg_trace_input_reg_31),
    .csr_reg_0(reg_trace_csr_reg_0),
    .csr_reg_1(reg_trace_csr_reg_1),
    .csr_reg_2(reg_trace_csr_reg_2),
    .csr_reg_3(reg_trace_csr_reg_3),
    .pc(reg_trace_pc)
  );
  assign Regfile_src1_value_MPORT_en = 1'h1;
  assign Regfile_src1_value_MPORT_addr = io_rs1;
  assign Regfile_src1_value_MPORT_data = Regfile[Regfile_src1_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_src2_value_MPORT_en = 1'h1;
  assign Regfile_src2_value_MPORT_addr = io_rs2;
  assign Regfile_src2_value_MPORT_data = Regfile[Regfile_src2_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_value_MPORT_en = 1'h1;
  assign Regfile_reg_value_MPORT_addr = io_rd;
  assign Regfile_reg_value_MPORT_data = Regfile[Regfile_reg_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_MPORT_4_en = 1'h1;
  assign Regfile_MPORT_4_addr = 5'h11;
  assign Regfile_MPORT_4_data = Regfile[Regfile_MPORT_4_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_en = 1'h1;
  assign Regfile_j_pc_MPORT_addr = io_rs1;
  assign Regfile_j_pc_MPORT_data = Regfile[Regfile_j_pc_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_1_en = 1'h1;
  assign Regfile_j_pc_MPORT_1_addr = io_rs2;
  assign Regfile_j_pc_MPORT_1_data = Regfile[Regfile_j_pc_MPORT_1_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_2_en = 1'h1;
  assign Regfile_j_pc_MPORT_2_addr = io_rs1;
  assign Regfile_j_pc_MPORT_2_data = Regfile[Regfile_j_pc_MPORT_2_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_3_en = 1'h1;
  assign Regfile_j_pc_MPORT_3_addr = io_rs2;
  assign Regfile_j_pc_MPORT_3_data = Regfile[Regfile_j_pc_MPORT_3_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_4_en = 1'h1;
  assign Regfile_j_pc_MPORT_4_addr = io_rs1;
  assign Regfile_j_pc_MPORT_4_data = Regfile[Regfile_j_pc_MPORT_4_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_5_en = 1'h1;
  assign Regfile_j_pc_MPORT_5_addr = io_rs2;
  assign Regfile_j_pc_MPORT_5_data = Regfile[Regfile_j_pc_MPORT_5_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_6_en = 1'h1;
  assign Regfile_j_pc_MPORT_6_addr = io_rs1;
  assign Regfile_j_pc_MPORT_6_data = Regfile[Regfile_j_pc_MPORT_6_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_7_en = 1'h1;
  assign Regfile_j_pc_MPORT_7_addr = io_rs2;
  assign Regfile_j_pc_MPORT_7_data = Regfile[Regfile_j_pc_MPORT_7_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_8_en = 1'h1;
  assign Regfile_j_pc_MPORT_8_addr = io_rs1;
  assign Regfile_j_pc_MPORT_8_data = Regfile[Regfile_j_pc_MPORT_8_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_9_en = 1'h1;
  assign Regfile_j_pc_MPORT_9_addr = io_rs2;
  assign Regfile_j_pc_MPORT_9_data = Regfile[Regfile_j_pc_MPORT_9_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_10_en = 1'h1;
  assign Regfile_j_pc_MPORT_10_addr = io_rs1;
  assign Regfile_j_pc_MPORT_10_data = Regfile[Regfile_j_pc_MPORT_10_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_11_en = 1'h1;
  assign Regfile_j_pc_MPORT_11_addr = io_rs2;
  assign Regfile_j_pc_MPORT_11_data = Regfile[Regfile_j_pc_MPORT_11_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_0_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_0_MPORT_addr = 5'h0;
  assign Regfile_reg_trace_io_input_reg_0_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_0_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_1_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_1_MPORT_addr = 5'h1;
  assign Regfile_reg_trace_io_input_reg_1_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_1_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_2_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_2_MPORT_addr = 5'h2;
  assign Regfile_reg_trace_io_input_reg_2_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_2_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_3_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_3_MPORT_addr = 5'h3;
  assign Regfile_reg_trace_io_input_reg_3_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_3_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_4_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_4_MPORT_addr = 5'h4;
  assign Regfile_reg_trace_io_input_reg_4_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_4_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_5_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_5_MPORT_addr = 5'h5;
  assign Regfile_reg_trace_io_input_reg_5_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_5_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_6_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_6_MPORT_addr = 5'h6;
  assign Regfile_reg_trace_io_input_reg_6_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_6_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_7_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_7_MPORT_addr = 5'h7;
  assign Regfile_reg_trace_io_input_reg_7_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_7_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_8_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_8_MPORT_addr = 5'h8;
  assign Regfile_reg_trace_io_input_reg_8_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_8_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_9_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_9_MPORT_addr = 5'h9;
  assign Regfile_reg_trace_io_input_reg_9_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_9_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_10_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_10_MPORT_addr = 5'ha;
  assign Regfile_reg_trace_io_input_reg_10_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_10_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_11_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_11_MPORT_addr = 5'hb;
  assign Regfile_reg_trace_io_input_reg_11_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_11_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_12_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_12_MPORT_addr = 5'hc;
  assign Regfile_reg_trace_io_input_reg_12_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_12_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_13_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_13_MPORT_addr = 5'hd;
  assign Regfile_reg_trace_io_input_reg_13_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_13_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_14_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_14_MPORT_addr = 5'he;
  assign Regfile_reg_trace_io_input_reg_14_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_14_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_15_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_15_MPORT_addr = 5'hf;
  assign Regfile_reg_trace_io_input_reg_15_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_15_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_16_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_16_MPORT_addr = 5'h10;
  assign Regfile_reg_trace_io_input_reg_16_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_16_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_17_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_17_MPORT_addr = 5'h11;
  assign Regfile_reg_trace_io_input_reg_17_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_17_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_18_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_18_MPORT_addr = 5'h12;
  assign Regfile_reg_trace_io_input_reg_18_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_18_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_19_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_19_MPORT_addr = 5'h13;
  assign Regfile_reg_trace_io_input_reg_19_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_19_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_20_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_20_MPORT_addr = 5'h14;
  assign Regfile_reg_trace_io_input_reg_20_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_20_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_21_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_21_MPORT_addr = 5'h15;
  assign Regfile_reg_trace_io_input_reg_21_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_21_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_22_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_22_MPORT_addr = 5'h16;
  assign Regfile_reg_trace_io_input_reg_22_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_22_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_23_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_23_MPORT_addr = 5'h17;
  assign Regfile_reg_trace_io_input_reg_23_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_23_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_24_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_24_MPORT_addr = 5'h18;
  assign Regfile_reg_trace_io_input_reg_24_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_24_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_25_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_25_MPORT_addr = 5'h19;
  assign Regfile_reg_trace_io_input_reg_25_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_25_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_26_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_26_MPORT_addr = 5'h1a;
  assign Regfile_reg_trace_io_input_reg_26_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_26_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_27_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_27_MPORT_addr = 5'h1b;
  assign Regfile_reg_trace_io_input_reg_27_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_27_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_28_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_28_MPORT_addr = 5'h1c;
  assign Regfile_reg_trace_io_input_reg_28_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_28_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_29_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_29_MPORT_addr = 5'h1d;
  assign Regfile_reg_trace_io_input_reg_29_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_29_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_30_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_30_MPORT_addr = 5'h1e;
  assign Regfile_reg_trace_io_input_reg_30_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_30_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_31_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_31_MPORT_addr = 5'h1f;
  assign Regfile_reg_trace_io_input_reg_31_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_31_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_data = Regfile[Regfile_mem_wdata_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_1_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_1_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_1_data = Regfile[Regfile_mem_wdata_MPORT_1_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_2_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_2_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_2_data = Regfile[Regfile_mem_wdata_MPORT_2_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_3_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_3_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_3_data = Regfile[Regfile_mem_wdata_MPORT_3_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_MPORT_data = _T_6 ? io_res2rd : reg_value;
  assign Regfile_MPORT_addr = io_rd;
  assign Regfile_MPORT_mask = 1'h1;
  assign Regfile_MPORT_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_io_res2rd_MPORT_1_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_1_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_1_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_1_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_io_res2rd_MPORT_2_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_2_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_2_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_2_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_csr_wdata_MPORT_en = 1'h1;
  assign CSR_Reg_csr_wdata_MPORT_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_csr_wdata_MPORT_data = CSR_Reg[CSR_Reg_csr_wdata_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_csr_wdata_MPORT_1_en = 1'h1;
  assign CSR_Reg_csr_wdata_MPORT_1_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_csr_wdata_MPORT_1_data = CSR_Reg[CSR_Reg_csr_wdata_MPORT_1_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_2_en = 1'h1;
  assign CSR_Reg_MPORT_2_addr = 2'h1;
  assign CSR_Reg_MPORT_2_data = CSR_Reg[CSR_Reg_MPORT_2_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_5_en = 1'h1;
  assign CSR_Reg_MPORT_5_addr = 2'h3;
  assign CSR_Reg_MPORT_5_data = CSR_Reg[CSR_Reg_MPORT_5_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_7_en = 1'h1;
  assign CSR_Reg_MPORT_7_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_MPORT_7_data = CSR_Reg[CSR_Reg_MPORT_7_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_j_pc_MPORT_12_en = 1'h1;
  assign CSR_Reg_j_pc_MPORT_12_addr = 2'h0;
  assign CSR_Reg_j_pc_MPORT_12_data = CSR_Reg[CSR_Reg_j_pc_MPORT_12_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_j_pc_MPORT_13_en = 1'h1;
  assign CSR_Reg_j_pc_MPORT_13_addr = 2'h1;
  assign CSR_Reg_j_pc_MPORT_13_data = CSR_Reg[CSR_Reg_j_pc_MPORT_13_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr = 2'h0;
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr = 2'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr = 2'h2;
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_1_data = _T_9 ? io_pc : CSR_Reg_MPORT_2_data;
  assign CSR_Reg_MPORT_1_addr = 2'h1;
  assign CSR_Reg_MPORT_1_mask = 1'h1;
  assign CSR_Reg_MPORT_1_en = 1'h1;
  assign CSR_Reg_MPORT_3_data = _T_9 ? Regfile_MPORT_4_data : CSR_Reg_MPORT_5_data;
  assign CSR_Reg_MPORT_3_addr = 2'h3;
  assign CSR_Reg_MPORT_3_mask = 1'h1;
  assign CSR_Reg_MPORT_3_en = 1'h1;
  assign CSR_Reg_MPORT_6_data = _T_14 ? csr_wdata : CSR_Reg_MPORT_7_data;
  assign CSR_Reg_MPORT_6_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_MPORT_6_mask = 1'h1;
  assign CSR_Reg_MPORT_6_en = 1'h1;
  assign io_pc_next = pc_next; // @[EXU_AXI.scala 162:16]
  assign io_res2rd = _io_res2rd_T_208[63:0]; // @[EXU_AXI.scala 72:15]
  assign io_inst_store = io_ctrl_sign_Writemem_en; // @[EXU_AXI.scala 188:19]
  assign io_inst_load = io_ctrl_sign_Readmem_en; // @[EXU_AXI.scala 189:18]
  assign io_Mem_addr = add_res[31:0]; // @[EXU_AXI.scala 190:17]
  assign io_Mem_wdata = 32'h27 == io_inst_now ? {{32'd0}, _mem_wdata_T_9[31:0]} : _mem_wdata_T_16; // @[Mux.scala 81:58]
  assign io_Mem_wstrb = io_ctrl_sign_Wmask; // @[EXU_AXI.scala 192:18]
  assign reg_trace_input_reg_0 = Regfile_reg_trace_io_input_reg_0_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_1 = Regfile_reg_trace_io_input_reg_1_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_2 = Regfile_reg_trace_io_input_reg_2_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_3 = Regfile_reg_trace_io_input_reg_3_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_4 = Regfile_reg_trace_io_input_reg_4_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_5 = Regfile_reg_trace_io_input_reg_5_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_6 = Regfile_reg_trace_io_input_reg_6_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_7 = Regfile_reg_trace_io_input_reg_7_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_8 = Regfile_reg_trace_io_input_reg_8_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_9 = Regfile_reg_trace_io_input_reg_9_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_10 = Regfile_reg_trace_io_input_reg_10_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_11 = Regfile_reg_trace_io_input_reg_11_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_12 = Regfile_reg_trace_io_input_reg_12_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_13 = Regfile_reg_trace_io_input_reg_13_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_14 = Regfile_reg_trace_io_input_reg_14_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_15 = Regfile_reg_trace_io_input_reg_15_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_16 = Regfile_reg_trace_io_input_reg_16_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_17 = Regfile_reg_trace_io_input_reg_17_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_18 = Regfile_reg_trace_io_input_reg_18_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_19 = Regfile_reg_trace_io_input_reg_19_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_20 = Regfile_reg_trace_io_input_reg_20_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_21 = Regfile_reg_trace_io_input_reg_21_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_22 = Regfile_reg_trace_io_input_reg_22_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_23 = Regfile_reg_trace_io_input_reg_23_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_24 = Regfile_reg_trace_io_input_reg_24_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_25 = Regfile_reg_trace_io_input_reg_25_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_26 = Regfile_reg_trace_io_input_reg_26_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_27 = Regfile_reg_trace_io_input_reg_27_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_28 = Regfile_reg_trace_io_input_reg_28_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_29 = Regfile_reg_trace_io_input_reg_29_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_30 = Regfile_reg_trace_io_input_reg_30_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_31 = Regfile_reg_trace_io_input_reg_31_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_csr_reg_0 = CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_1 = CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_2 = CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_3 = 64'h0; // @[EXU_AXI.scala 167:{36,36}]
  assign reg_trace_pc = io_pc; // @[EXU_AXI.scala 166:21]
  always @(posedge clock) begin
    if (Regfile_MPORT_en & Regfile_MPORT_mask) begin
      Regfile[Regfile_MPORT_addr] <= Regfile_MPORT_data; // @[EXU_AXI.scala 37:22]
    end
    if (CSR_Reg_MPORT_1_en & CSR_Reg_MPORT_1_mask) begin
      CSR_Reg[CSR_Reg_MPORT_1_addr] <= CSR_Reg_MPORT_1_data; // @[EXU_AXI.scala 38:22]
    end
    if (CSR_Reg_MPORT_3_en & CSR_Reg_MPORT_3_mask) begin
      CSR_Reg[CSR_Reg_MPORT_3_addr] <= CSR_Reg_MPORT_3_data; // @[EXU_AXI.scala 38:22]
    end
    if (CSR_Reg_MPORT_6_en & CSR_Reg_MPORT_6_mask) begin
      CSR_Reg[CSR_Reg_MPORT_6_addr] <= CSR_Reg_MPORT_6_data; // @[EXU_AXI.scala 38:22]
    end
    if (reset) begin // @[EXU_AXI.scala 158:26]
      pc_next <= 64'h0; // @[EXU_AXI.scala 158:26]
    end else if (io_inst_valid) begin // @[EXU_AXI.scala 159:24]
      if (32'h3e == io_inst_now) begin // @[Mux.scala 81:58]
        pc_next <= _j_pc_T_46;
      end else if (32'h3d == io_inst_now) begin // @[Mux.scala 81:58]
        pc_next <= CSR_Reg_j_pc_MPORT_12_data;
      end else begin
        pc_next <= _j_pc_T_62;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    Regfile[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    CSR_Reg[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  pc_next = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top(
  input         clock,
  input         reset,
  output [31:0] io_inst,
  output [63:0] io_pc,
  output [63:0] io_pc_next,
  output [63:0] io_outval,
  output        io_step
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  axi_clock; // @[top.scala 18:21]
  wire  axi_reset; // @[top.scala 18:21]
  wire [31:0] axi_io_axi_in_araddr; // @[top.scala 18:21]
  wire  axi_io_axi_in_arvalid; // @[top.scala 18:21]
  wire  axi_io_axi_in_rready; // @[top.scala 18:21]
  wire [31:0] axi_io_axi_in_awaddr; // @[top.scala 18:21]
  wire  axi_io_axi_in_awvalid; // @[top.scala 18:21]
  wire [31:0] axi_io_axi_in_wdata; // @[top.scala 18:21]
  wire [7:0] axi_io_axi_in_wstrb; // @[top.scala 18:21]
  wire  axi_io_axi_in_wvalid; // @[top.scala 18:21]
  wire  axi_io_axi_in_bready; // @[top.scala 18:21]
  wire  axi_io_axi_out_arready; // @[top.scala 18:21]
  wire [63:0] axi_io_axi_out_rdata; // @[top.scala 18:21]
  wire  axi_io_axi_out_rvalid; // @[top.scala 18:21]
  wire  axi_io_axi_out_awready; // @[top.scala 18:21]
  wire  axi_io_axi_out_wready; // @[top.scala 18:21]
  wire  axi_io_axi_out_bvalid; // @[top.scala 18:21]
  wire  lsu_step_clock; // @[top.scala 19:26]
  wire  lsu_step_reset; // @[top.scala 19:26]
  wire  lsu_step_io_inst_store; // @[top.scala 19:26]
  wire  lsu_step_io_inst_load; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_mem_addr; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_mem_wdata; // @[top.scala 19:26]
  wire [7:0] lsu_step_io_mem_wstrb; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_mem_rdata; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_arready; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_axi_in_rdata; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_rvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_awready; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_wready; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_bvalid; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_axi_out_araddr; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_arvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_rready; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_axi_out_awaddr; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_awvalid; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_axi_out_wdata; // @[top.scala 19:26]
  wire [7:0] lsu_step_io_axi_out_wstrb; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_wvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_bready; // @[top.scala 19:26]
  wire  arbiter_clock; // @[top.scala 20:25]
  wire  arbiter_reset; // @[top.scala 20:25]
  wire [31:0] arbiter_io_ifu_axi_in_araddr; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_in_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_in_rready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_ifu_axi_out_rdata; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_out_rvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_lsu_axi_in_araddr; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_rready; // @[top.scala 20:25]
  wire [31:0] arbiter_io_lsu_axi_in_awaddr; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_awvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_lsu_axi_in_wdata; // @[top.scala 20:25]
  wire [7:0] arbiter_io_lsu_axi_in_wstrb; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_wvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_bready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_arready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_lsu_axi_out_rdata; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_rvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_awready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_wready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_bvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_arready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_axi_in_rdata; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_rvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_awready; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_wready; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_bvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_axi_out_araddr; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_rready; // @[top.scala 20:25]
  wire [31:0] arbiter_io_axi_out_awaddr; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_awvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_axi_out_wdata; // @[top.scala 20:25]
  wire [7:0] arbiter_io_axi_out_wstrb; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_wvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_bready; // @[top.scala 20:25]
  wire  ifu_step_clock; // @[top.scala 21:26]
  wire  ifu_step_reset; // @[top.scala 21:26]
  wire [63:0] ifu_step_io_pc; // @[top.scala 21:26]
  wire  ifu_step_io_pc_valid; // @[top.scala 21:26]
  wire  ifu_step_io_inst_valid; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_inst; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_inst_reg; // @[top.scala 21:26]
  wire [63:0] ifu_step_io_axi_in_rdata; // @[top.scala 21:26]
  wire  ifu_step_io_axi_in_rvalid; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_axi_out_araddr; // @[top.scala 21:26]
  wire  ifu_step_io_axi_out_arvalid; // @[top.scala 21:26]
  wire  ifu_step_io_axi_out_rready; // @[top.scala 21:26]
  wire  i_cache_clock; // @[top.scala 22:25]
  wire  i_cache_reset; // @[top.scala 22:25]
  wire [31:0] i_cache_io_from_ifu_araddr; // @[top.scala 22:25]
  wire  i_cache_io_from_ifu_arvalid; // @[top.scala 22:25]
  wire  i_cache_io_from_ifu_rready; // @[top.scala 22:25]
  wire [63:0] i_cache_io_to_ifu_rdata; // @[top.scala 22:25]
  wire  i_cache_io_to_ifu_rvalid; // @[top.scala 22:25]
  wire [31:0] i_cache_io_to_axi_araddr; // @[top.scala 22:25]
  wire  i_cache_io_to_axi_arvalid; // @[top.scala 22:25]
  wire  i_cache_io_to_axi_rready; // @[top.scala 22:25]
  wire [63:0] i_cache_io_from_axi_rdata; // @[top.scala 22:25]
  wire  i_cache_io_from_axi_rvalid; // @[top.scala 22:25]
  wire  d_cache_clock; // @[top.scala 23:25]
  wire  d_cache_reset; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_araddr; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_arvalid; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_rready; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_awaddr; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_awvalid; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_wdata; // @[top.scala 23:25]
  wire [7:0] d_cache_io_from_lsu_wstrb; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_wvalid; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_bready; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_arready; // @[top.scala 23:25]
  wire [63:0] d_cache_io_to_lsu_rdata; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_rvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_awready; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_wready; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_bvalid; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_araddr; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_arvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_rready; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_awaddr; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_awvalid; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_wdata; // @[top.scala 23:25]
  wire [7:0] d_cache_io_to_axi_wstrb; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_wvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_bready; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_arready; // @[top.scala 23:25]
  wire [63:0] d_cache_io_from_axi_rdata; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_rvalid; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_awready; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_wready; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_bvalid; // @[top.scala 23:25]
  wire [31:0] idu_step_io_inst; // @[top.scala 46:26]
  wire [31:0] idu_step_io_inst_now; // @[top.scala 46:26]
  wire [4:0] idu_step_io_rs1; // @[top.scala 46:26]
  wire [4:0] idu_step_io_rs2; // @[top.scala 46:26]
  wire [4:0] idu_step_io_rd; // @[top.scala 46:26]
  wire [63:0] idu_step_io_imm; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_reg_write; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_csr_write; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_Writemem_en; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_Readmem_en; // @[top.scala 46:26]
  wire [7:0] idu_step_io_ctrl_sign_Wmask; // @[top.scala 46:26]
  wire  exu_step_clock; // @[top.scala 51:26]
  wire  exu_step_reset; // @[top.scala 51:26]
  wire [63:0] exu_step_io_pc; // @[top.scala 51:26]
  wire [63:0] exu_step_io_pc_next; // @[top.scala 51:26]
  wire [31:0] exu_step_io_inst_now; // @[top.scala 51:26]
  wire [4:0] exu_step_io_rs1; // @[top.scala 51:26]
  wire [4:0] exu_step_io_rs2; // @[top.scala 51:26]
  wire [4:0] exu_step_io_rd; // @[top.scala 51:26]
  wire [63:0] exu_step_io_imm; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_reg_write; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_csr_write; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_Writemem_en; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_Readmem_en; // @[top.scala 51:26]
  wire [7:0] exu_step_io_ctrl_sign_Wmask; // @[top.scala 51:26]
  wire [63:0] exu_step_io_res2rd; // @[top.scala 51:26]
  wire  exu_step_io_inst_valid; // @[top.scala 51:26]
  wire  exu_step_io_inst_store; // @[top.scala 51:26]
  wire  exu_step_io_inst_load; // @[top.scala 51:26]
  wire [31:0] exu_step_io_Mem_addr; // @[top.scala 51:26]
  wire [63:0] exu_step_io_Mem_rdata; // @[top.scala 51:26]
  wire [63:0] exu_step_io_Mem_wdata; // @[top.scala 51:26]
  wire [7:0] exu_step_io_Mem_wstrb; // @[top.scala 51:26]
  wire  exu_step_io_rdata_valid; // @[top.scala 51:26]
  wire [31:0] dpi_flag; // @[top.scala 73:21]
  wire [31:0] dpi_ecall_flag; // @[top.scala 73:21]
  reg [63:0] pc_now; // @[top.scala 15:25]
  reg  execute_end; // @[top.scala 17:30]
  reg  pc_valid; // @[top.scala 87:27]
  reg  diff_step; // @[top.scala 90:28]
  AXI axi ( // @[top.scala 18:21]
    .clock(axi_clock),
    .reset(axi_reset),
    .io_axi_in_araddr(axi_io_axi_in_araddr),
    .io_axi_in_arvalid(axi_io_axi_in_arvalid),
    .io_axi_in_rready(axi_io_axi_in_rready),
    .io_axi_in_awaddr(axi_io_axi_in_awaddr),
    .io_axi_in_awvalid(axi_io_axi_in_awvalid),
    .io_axi_in_wdata(axi_io_axi_in_wdata),
    .io_axi_in_wstrb(axi_io_axi_in_wstrb),
    .io_axi_in_wvalid(axi_io_axi_in_wvalid),
    .io_axi_in_bready(axi_io_axi_in_bready),
    .io_axi_out_arready(axi_io_axi_out_arready),
    .io_axi_out_rdata(axi_io_axi_out_rdata),
    .io_axi_out_rvalid(axi_io_axi_out_rvalid),
    .io_axi_out_awready(axi_io_axi_out_awready),
    .io_axi_out_wready(axi_io_axi_out_wready),
    .io_axi_out_bvalid(axi_io_axi_out_bvalid)
  );
  LSU lsu_step ( // @[top.scala 19:26]
    .clock(lsu_step_clock),
    .reset(lsu_step_reset),
    .io_inst_store(lsu_step_io_inst_store),
    .io_inst_load(lsu_step_io_inst_load),
    .io_mem_addr(lsu_step_io_mem_addr),
    .io_mem_wdata(lsu_step_io_mem_wdata),
    .io_mem_wstrb(lsu_step_io_mem_wstrb),
    .io_mem_rdata(lsu_step_io_mem_rdata),
    .io_axi_in_arready(lsu_step_io_axi_in_arready),
    .io_axi_in_rdata(lsu_step_io_axi_in_rdata),
    .io_axi_in_rvalid(lsu_step_io_axi_in_rvalid),
    .io_axi_in_awready(lsu_step_io_axi_in_awready),
    .io_axi_in_wready(lsu_step_io_axi_in_wready),
    .io_axi_in_bvalid(lsu_step_io_axi_in_bvalid),
    .io_axi_out_araddr(lsu_step_io_axi_out_araddr),
    .io_axi_out_arvalid(lsu_step_io_axi_out_arvalid),
    .io_axi_out_rready(lsu_step_io_axi_out_rready),
    .io_axi_out_awaddr(lsu_step_io_axi_out_awaddr),
    .io_axi_out_awvalid(lsu_step_io_axi_out_awvalid),
    .io_axi_out_wdata(lsu_step_io_axi_out_wdata),
    .io_axi_out_wstrb(lsu_step_io_axi_out_wstrb),
    .io_axi_out_wvalid(lsu_step_io_axi_out_wvalid),
    .io_axi_out_bready(lsu_step_io_axi_out_bready)
  );
  AXI_ARBITER arbiter ( // @[top.scala 20:25]
    .clock(arbiter_clock),
    .reset(arbiter_reset),
    .io_ifu_axi_in_araddr(arbiter_io_ifu_axi_in_araddr),
    .io_ifu_axi_in_arvalid(arbiter_io_ifu_axi_in_arvalid),
    .io_ifu_axi_in_rready(arbiter_io_ifu_axi_in_rready),
    .io_ifu_axi_out_rdata(arbiter_io_ifu_axi_out_rdata),
    .io_ifu_axi_out_rvalid(arbiter_io_ifu_axi_out_rvalid),
    .io_lsu_axi_in_araddr(arbiter_io_lsu_axi_in_araddr),
    .io_lsu_axi_in_arvalid(arbiter_io_lsu_axi_in_arvalid),
    .io_lsu_axi_in_rready(arbiter_io_lsu_axi_in_rready),
    .io_lsu_axi_in_awaddr(arbiter_io_lsu_axi_in_awaddr),
    .io_lsu_axi_in_awvalid(arbiter_io_lsu_axi_in_awvalid),
    .io_lsu_axi_in_wdata(arbiter_io_lsu_axi_in_wdata),
    .io_lsu_axi_in_wstrb(arbiter_io_lsu_axi_in_wstrb),
    .io_lsu_axi_in_wvalid(arbiter_io_lsu_axi_in_wvalid),
    .io_lsu_axi_in_bready(arbiter_io_lsu_axi_in_bready),
    .io_lsu_axi_out_arready(arbiter_io_lsu_axi_out_arready),
    .io_lsu_axi_out_rdata(arbiter_io_lsu_axi_out_rdata),
    .io_lsu_axi_out_rvalid(arbiter_io_lsu_axi_out_rvalid),
    .io_lsu_axi_out_awready(arbiter_io_lsu_axi_out_awready),
    .io_lsu_axi_out_wready(arbiter_io_lsu_axi_out_wready),
    .io_lsu_axi_out_bvalid(arbiter_io_lsu_axi_out_bvalid),
    .io_axi_in_arready(arbiter_io_axi_in_arready),
    .io_axi_in_rdata(arbiter_io_axi_in_rdata),
    .io_axi_in_rvalid(arbiter_io_axi_in_rvalid),
    .io_axi_in_awready(arbiter_io_axi_in_awready),
    .io_axi_in_wready(arbiter_io_axi_in_wready),
    .io_axi_in_bvalid(arbiter_io_axi_in_bvalid),
    .io_axi_out_araddr(arbiter_io_axi_out_araddr),
    .io_axi_out_arvalid(arbiter_io_axi_out_arvalid),
    .io_axi_out_rready(arbiter_io_axi_out_rready),
    .io_axi_out_awaddr(arbiter_io_axi_out_awaddr),
    .io_axi_out_awvalid(arbiter_io_axi_out_awvalid),
    .io_axi_out_wdata(arbiter_io_axi_out_wdata),
    .io_axi_out_wstrb(arbiter_io_axi_out_wstrb),
    .io_axi_out_wvalid(arbiter_io_axi_out_wvalid),
    .io_axi_out_bready(arbiter_io_axi_out_bready)
  );
  IFU_AXI ifu_step ( // @[top.scala 21:26]
    .clock(ifu_step_clock),
    .reset(ifu_step_reset),
    .io_pc(ifu_step_io_pc),
    .io_pc_valid(ifu_step_io_pc_valid),
    .io_inst_valid(ifu_step_io_inst_valid),
    .io_inst(ifu_step_io_inst),
    .io_inst_reg(ifu_step_io_inst_reg),
    .io_axi_in_rdata(ifu_step_io_axi_in_rdata),
    .io_axi_in_rvalid(ifu_step_io_axi_in_rvalid),
    .io_axi_out_araddr(ifu_step_io_axi_out_araddr),
    .io_axi_out_arvalid(ifu_step_io_axi_out_arvalid),
    .io_axi_out_rready(ifu_step_io_axi_out_rready)
  );
  I_CACHE i_cache ( // @[top.scala 22:25]
    .clock(i_cache_clock),
    .reset(i_cache_reset),
    .io_from_ifu_araddr(i_cache_io_from_ifu_araddr),
    .io_from_ifu_arvalid(i_cache_io_from_ifu_arvalid),
    .io_from_ifu_rready(i_cache_io_from_ifu_rready),
    .io_to_ifu_rdata(i_cache_io_to_ifu_rdata),
    .io_to_ifu_rvalid(i_cache_io_to_ifu_rvalid),
    .io_to_axi_araddr(i_cache_io_to_axi_araddr),
    .io_to_axi_arvalid(i_cache_io_to_axi_arvalid),
    .io_to_axi_rready(i_cache_io_to_axi_rready),
    .io_from_axi_rdata(i_cache_io_from_axi_rdata),
    .io_from_axi_rvalid(i_cache_io_from_axi_rvalid)
  );
  D_CACHE d_cache ( // @[top.scala 23:25]
    .clock(d_cache_clock),
    .reset(d_cache_reset),
    .io_from_lsu_araddr(d_cache_io_from_lsu_araddr),
    .io_from_lsu_arvalid(d_cache_io_from_lsu_arvalid),
    .io_from_lsu_rready(d_cache_io_from_lsu_rready),
    .io_from_lsu_awaddr(d_cache_io_from_lsu_awaddr),
    .io_from_lsu_awvalid(d_cache_io_from_lsu_awvalid),
    .io_from_lsu_wdata(d_cache_io_from_lsu_wdata),
    .io_from_lsu_wstrb(d_cache_io_from_lsu_wstrb),
    .io_from_lsu_wvalid(d_cache_io_from_lsu_wvalid),
    .io_from_lsu_bready(d_cache_io_from_lsu_bready),
    .io_to_lsu_arready(d_cache_io_to_lsu_arready),
    .io_to_lsu_rdata(d_cache_io_to_lsu_rdata),
    .io_to_lsu_rvalid(d_cache_io_to_lsu_rvalid),
    .io_to_lsu_awready(d_cache_io_to_lsu_awready),
    .io_to_lsu_wready(d_cache_io_to_lsu_wready),
    .io_to_lsu_bvalid(d_cache_io_to_lsu_bvalid),
    .io_to_axi_araddr(d_cache_io_to_axi_araddr),
    .io_to_axi_arvalid(d_cache_io_to_axi_arvalid),
    .io_to_axi_rready(d_cache_io_to_axi_rready),
    .io_to_axi_awaddr(d_cache_io_to_axi_awaddr),
    .io_to_axi_awvalid(d_cache_io_to_axi_awvalid),
    .io_to_axi_wdata(d_cache_io_to_axi_wdata),
    .io_to_axi_wstrb(d_cache_io_to_axi_wstrb),
    .io_to_axi_wvalid(d_cache_io_to_axi_wvalid),
    .io_to_axi_bready(d_cache_io_to_axi_bready),
    .io_from_axi_arready(d_cache_io_from_axi_arready),
    .io_from_axi_rdata(d_cache_io_from_axi_rdata),
    .io_from_axi_rvalid(d_cache_io_from_axi_rvalid),
    .io_from_axi_awready(d_cache_io_from_axi_awready),
    .io_from_axi_wready(d_cache_io_from_axi_wready),
    .io_from_axi_bvalid(d_cache_io_from_axi_bvalid)
  );
  IDU idu_step ( // @[top.scala 46:26]
    .io_inst(idu_step_io_inst),
    .io_inst_now(idu_step_io_inst_now),
    .io_rs1(idu_step_io_rs1),
    .io_rs2(idu_step_io_rs2),
    .io_rd(idu_step_io_rd),
    .io_imm(idu_step_io_imm),
    .io_ctrl_sign_reg_write(idu_step_io_ctrl_sign_reg_write),
    .io_ctrl_sign_csr_write(idu_step_io_ctrl_sign_csr_write),
    .io_ctrl_sign_src2_is_imm(idu_step_io_ctrl_sign_src2_is_imm),
    .io_ctrl_sign_src1_is_pc(idu_step_io_ctrl_sign_src1_is_pc),
    .io_ctrl_sign_Writemem_en(idu_step_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(idu_step_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(idu_step_io_ctrl_sign_Wmask)
  );
  EXU_AXI exu_step ( // @[top.scala 51:26]
    .clock(exu_step_clock),
    .reset(exu_step_reset),
    .io_pc(exu_step_io_pc),
    .io_pc_next(exu_step_io_pc_next),
    .io_inst_now(exu_step_io_inst_now),
    .io_rs1(exu_step_io_rs1),
    .io_rs2(exu_step_io_rs2),
    .io_rd(exu_step_io_rd),
    .io_imm(exu_step_io_imm),
    .io_ctrl_sign_reg_write(exu_step_io_ctrl_sign_reg_write),
    .io_ctrl_sign_csr_write(exu_step_io_ctrl_sign_csr_write),
    .io_ctrl_sign_src2_is_imm(exu_step_io_ctrl_sign_src2_is_imm),
    .io_ctrl_sign_src1_is_pc(exu_step_io_ctrl_sign_src1_is_pc),
    .io_ctrl_sign_Writemem_en(exu_step_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(exu_step_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(exu_step_io_ctrl_sign_Wmask),
    .io_res2rd(exu_step_io_res2rd),
    .io_inst_valid(exu_step_io_inst_valid),
    .io_inst_store(exu_step_io_inst_store),
    .io_inst_load(exu_step_io_inst_load),
    .io_Mem_addr(exu_step_io_Mem_addr),
    .io_Mem_rdata(exu_step_io_Mem_rdata),
    .io_Mem_wdata(exu_step_io_Mem_wdata),
    .io_Mem_wstrb(exu_step_io_Mem_wstrb),
    .io_rdata_valid(exu_step_io_rdata_valid)
  );
  DPI dpi ( // @[top.scala 73:21]
    .flag(dpi_flag),
    .ecall_flag(dpi_ecall_flag)
  );
  assign io_inst = ifu_step_io_inst; // @[top.scala 25:13]
  assign io_pc = pc_now; // @[top.scala 16:11]
  assign io_pc_next = exu_step_io_pc_next; // @[top.scala 94:16]
  assign io_outval = exu_step_io_res2rd; // @[top.scala 69:15]
  assign io_step = diff_step; // @[top.scala 92:13]
  assign axi_clock = clock;
  assign axi_reset = reset;
  assign axi_io_axi_in_araddr = arbiter_io_axi_out_araddr; // @[top.scala 43:19]
  assign axi_io_axi_in_arvalid = arbiter_io_axi_out_arvalid; // @[top.scala 43:19]
  assign axi_io_axi_in_rready = arbiter_io_axi_out_rready; // @[top.scala 43:19]
  assign axi_io_axi_in_awaddr = arbiter_io_axi_out_awaddr; // @[top.scala 43:19]
  assign axi_io_axi_in_awvalid = arbiter_io_axi_out_awvalid; // @[top.scala 43:19]
  assign axi_io_axi_in_wdata = arbiter_io_axi_out_wdata; // @[top.scala 43:19]
  assign axi_io_axi_in_wstrb = arbiter_io_axi_out_wstrb; // @[top.scala 43:19]
  assign axi_io_axi_in_wvalid = arbiter_io_axi_out_wvalid; // @[top.scala 43:19]
  assign axi_io_axi_in_bready = arbiter_io_axi_out_bready; // @[top.scala 43:19]
  assign lsu_step_clock = clock;
  assign lsu_step_reset = reset;
  assign lsu_step_io_inst_store = exu_step_io_inst_store; // @[top.scala 61:28]
  assign lsu_step_io_inst_load = exu_step_io_inst_load; // @[top.scala 60:27]
  assign lsu_step_io_mem_addr = exu_step_io_Mem_addr; // @[top.scala 62:26]
  assign lsu_step_io_mem_wdata = exu_step_io_Mem_wdata; // @[top.scala 63:27]
  assign lsu_step_io_mem_wstrb = exu_step_io_Mem_wstrb; // @[top.scala 64:27]
  assign lsu_step_io_axi_in_arready = d_cache_io_to_lsu_arready; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_rdata = d_cache_io_to_lsu_rdata; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_rvalid = d_cache_io_to_lsu_rvalid; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_awready = d_cache_io_to_lsu_awready; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_wready = d_cache_io_to_lsu_wready; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_bvalid = d_cache_io_to_lsu_bvalid; // @[top.scala 36:24]
  assign arbiter_clock = clock;
  assign arbiter_reset = reset;
  assign arbiter_io_ifu_axi_in_araddr = i_cache_io_to_axi_araddr; // @[top.scala 26:27]
  assign arbiter_io_ifu_axi_in_arvalid = i_cache_io_to_axi_arvalid; // @[top.scala 26:27]
  assign arbiter_io_ifu_axi_in_rready = i_cache_io_to_axi_rready; // @[top.scala 26:27]
  assign arbiter_io_lsu_axi_in_araddr = d_cache_io_to_axi_araddr; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_arvalid = d_cache_io_to_axi_arvalid; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_rready = d_cache_io_to_axi_rready; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_awaddr = d_cache_io_to_axi_awaddr; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_awvalid = d_cache_io_to_axi_awvalid; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_wdata = d_cache_io_to_axi_wdata; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_wstrb = d_cache_io_to_axi_wstrb; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_wvalid = d_cache_io_to_axi_wvalid; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_bready = d_cache_io_to_axi_bready; // @[top.scala 34:27]
  assign arbiter_io_axi_in_arready = axi_io_axi_out_arready; // @[top.scala 42:23]
  assign arbiter_io_axi_in_rdata = axi_io_axi_out_rdata; // @[top.scala 42:23]
  assign arbiter_io_axi_in_rvalid = axi_io_axi_out_rvalid; // @[top.scala 42:23]
  assign arbiter_io_axi_in_awready = axi_io_axi_out_awready; // @[top.scala 42:23]
  assign arbiter_io_axi_in_wready = axi_io_axi_out_wready; // @[top.scala 42:23]
  assign arbiter_io_axi_in_bvalid = axi_io_axi_out_bvalid; // @[top.scala 42:23]
  assign ifu_step_clock = clock;
  assign ifu_step_reset = reset;
  assign ifu_step_io_pc = pc_now; // @[top.scala 24:20]
  assign ifu_step_io_pc_valid = pc_valid; // @[top.scala 89:26]
  assign ifu_step_io_axi_in_rdata = i_cache_io_to_ifu_rdata; // @[top.scala 28:24]
  assign ifu_step_io_axi_in_rvalid = i_cache_io_to_ifu_rvalid; // @[top.scala 28:24]
  assign i_cache_clock = clock;
  assign i_cache_reset = reset;
  assign i_cache_io_from_ifu_araddr = ifu_step_io_axi_out_araddr; // @[top.scala 29:25]
  assign i_cache_io_from_ifu_arvalid = ifu_step_io_axi_out_arvalid; // @[top.scala 29:25]
  assign i_cache_io_from_ifu_rready = ifu_step_io_axi_out_rready; // @[top.scala 29:25]
  assign i_cache_io_from_axi_rdata = arbiter_io_ifu_axi_out_rdata; // @[top.scala 27:25]
  assign i_cache_io_from_axi_rvalid = arbiter_io_ifu_axi_out_rvalid; // @[top.scala 27:25]
  assign d_cache_clock = clock;
  assign d_cache_reset = reset;
  assign d_cache_io_from_lsu_araddr = lsu_step_io_axi_out_araddr; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_arvalid = lsu_step_io_axi_out_arvalid; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_rready = lsu_step_io_axi_out_rready; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_awaddr = lsu_step_io_axi_out_awaddr; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_awvalid = lsu_step_io_axi_out_awvalid; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_wdata = lsu_step_io_axi_out_wdata; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_wstrb = lsu_step_io_axi_out_wstrb; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_wvalid = lsu_step_io_axi_out_wvalid; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_bready = lsu_step_io_axi_out_bready; // @[top.scala 37:25]
  assign d_cache_io_from_axi_arready = arbiter_io_lsu_axi_out_arready; // @[top.scala 35:25]
  assign d_cache_io_from_axi_rdata = arbiter_io_lsu_axi_out_rdata; // @[top.scala 35:25]
  assign d_cache_io_from_axi_rvalid = arbiter_io_lsu_axi_out_rvalid; // @[top.scala 35:25]
  assign d_cache_io_from_axi_awready = arbiter_io_lsu_axi_out_awready; // @[top.scala 35:25]
  assign d_cache_io_from_axi_wready = arbiter_io_lsu_axi_out_wready; // @[top.scala 35:25]
  assign d_cache_io_from_axi_bvalid = arbiter_io_lsu_axi_out_bvalid; // @[top.scala 35:25]
  assign idu_step_io_inst = ~ifu_step_io_inst_valid & ~pc_valid & ~execute_end ? ifu_step_io_inst_reg : ifu_step_io_inst
    ; // @[top.scala 96:28]
  assign exu_step_clock = clock;
  assign exu_step_reset = reset;
  assign exu_step_io_pc = pc_now; // @[top.scala 52:20]
  assign exu_step_io_inst_now = idu_step_io_inst_now; // @[top.scala 53:26]
  assign exu_step_io_rs1 = idu_step_io_rs1; // @[top.scala 55:21]
  assign exu_step_io_rs2 = idu_step_io_rs2; // @[top.scala 56:21]
  assign exu_step_io_rd = idu_step_io_rd; // @[top.scala 57:20]
  assign exu_step_io_imm = idu_step_io_imm; // @[top.scala 58:21]
  assign exu_step_io_ctrl_sign_reg_write = idu_step_io_ctrl_sign_reg_write; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_csr_write = idu_step_io_ctrl_sign_csr_write; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_src2_is_imm = idu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_src1_is_pc = idu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_Writemem_en = idu_step_io_ctrl_sign_Writemem_en; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_Readmem_en = idu_step_io_ctrl_sign_Readmem_en; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_Wmask = idu_step_io_ctrl_sign_Wmask; // @[top.scala 59:27]
  assign exu_step_io_inst_valid = ifu_step_io_inst_valid; // @[top.scala 68:28]
  assign exu_step_io_Mem_rdata = lsu_step_io_mem_rdata; // @[top.scala 65:27]
  assign exu_step_io_rdata_valid = lsu_step_io_axi_in_rvalid; // @[top.scala 66:29]
  assign dpi_flag = {{31'd0}, idu_step_io_inst_now == 32'h2}; // @[top.scala 74:17]
  assign dpi_ecall_flag = {{31'd0}, idu_step_io_inst_now == 32'h3d}; // @[top.scala 75:23]
  always @(posedge clock) begin
    if (reset) begin // @[top.scala 15:25]
      pc_now <= 64'h80000000; // @[top.scala 15:25]
    end else if (execute_end) begin // @[top.scala 93:18]
      pc_now <= exu_step_io_pc_next;
    end
    if (reset) begin // @[top.scala 17:30]
      execute_end <= 1'h0; // @[top.scala 17:30]
    end else if (exu_step_io_inst_store) begin // @[top.scala 85:23]
      execute_end <= lsu_step_io_axi_in_bvalid;
    end else if (exu_step_io_inst_load) begin // @[top.scala 85:76]
      execute_end <= lsu_step_io_axi_in_rvalid;
    end else begin
      execute_end <= ifu_step_io_inst_valid;
    end
    pc_valid <= reset | execute_end; // @[top.scala 87:{27,27} 88:14]
    if (reset) begin // @[top.scala 90:28]
      diff_step <= 1'h0; // @[top.scala 90:28]
    end else begin
      diff_step <= execute_end; // @[top.scala 91:15]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"pc : %x inst:%x execute_end : %d\n\n",pc_now,idu_step_io_inst,execute_end); // @[top.scala 86:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc_now = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  execute_end = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pc_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  diff_step = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
