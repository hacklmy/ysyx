module D_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_lsu_araddr,
  input         io_from_lsu_arvalid,
  input         io_from_lsu_rready,
  input  [31:0] io_from_lsu_awaddr,
  input         io_from_lsu_awvalid,
  input  [31:0] io_from_lsu_wdata,
  input  [7:0]  io_from_lsu_wstrb,
  input         io_from_lsu_wvalid,
  input         io_from_lsu_bready,
  output        io_to_lsu_arready,
  output [63:0] io_to_lsu_rdata,
  output        io_to_lsu_rvalid,
  output        io_to_lsu_awready,
  output        io_to_lsu_wready,
  output        io_to_lsu_bvalid,
  output [31:0] io_to_axi_araddr,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  output [31:0] io_to_axi_awaddr,
  output        io_to_axi_awvalid,
  output [31:0] io_to_axi_wdata,
  output [7:0]  io_to_axi_wstrb,
  output        io_to_axi_wvalid,
  output        io_to_axi_bready,
  input         io_from_axi_arready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rvalid,
  input         io_from_axi_awready,
  input         io_from_axi_wready,
  input         io_from_axi_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [63:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [63:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = ~reset; // @[d_cache.scala 15:11]
  reg [63:0] ram_0_0; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_1; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_2; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_3; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_4; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_5; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_6; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_7; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_8; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_9; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_10; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_11; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_12; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_13; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_14; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_15; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_16; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_17; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_18; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_19; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_20; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_21; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_22; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_23; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_24; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_25; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_26; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_27; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_28; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_29; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_30; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_31; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_32; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_33; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_34; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_35; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_36; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_37; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_38; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_39; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_40; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_41; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_42; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_43; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_44; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_45; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_46; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_47; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_48; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_49; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_50; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_51; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_52; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_53; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_54; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_55; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_56; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_57; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_58; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_59; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_60; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_61; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_62; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_63; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_64; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_65; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_66; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_67; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_68; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_69; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_70; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_71; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_72; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_73; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_74; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_75; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_76; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_77; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_78; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_79; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_80; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_81; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_82; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_83; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_84; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_85; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_86; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_87; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_88; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_89; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_90; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_91; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_92; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_93; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_94; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_95; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_96; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_97; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_98; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_99; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_100; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_101; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_102; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_103; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_104; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_105; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_106; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_107; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_108; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_109; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_110; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_111; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_112; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_113; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_114; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_115; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_116; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_117; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_118; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_119; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_120; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_121; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_122; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_123; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_124; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_125; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_126; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_127; // @[d_cache.scala 18:24]
  reg [63:0] ram_1_0; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_1; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_2; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_3; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_4; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_5; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_6; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_7; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_8; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_9; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_10; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_11; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_12; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_13; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_14; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_15; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_16; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_17; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_18; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_19; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_20; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_21; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_22; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_23; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_24; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_25; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_26; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_27; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_28; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_29; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_30; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_31; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_32; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_33; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_34; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_35; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_36; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_37; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_38; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_39; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_40; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_41; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_42; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_43; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_44; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_45; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_46; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_47; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_48; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_49; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_50; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_51; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_52; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_53; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_54; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_55; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_56; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_57; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_58; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_59; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_60; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_61; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_62; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_63; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_64; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_65; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_66; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_67; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_68; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_69; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_70; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_71; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_72; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_73; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_74; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_75; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_76; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_77; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_78; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_79; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_80; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_81; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_82; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_83; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_84; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_85; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_86; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_87; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_88; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_89; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_90; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_91; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_92; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_93; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_94; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_95; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_96; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_97; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_98; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_99; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_100; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_101; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_102; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_103; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_104; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_105; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_106; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_107; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_108; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_109; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_110; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_111; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_112; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_113; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_114; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_115; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_116; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_117; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_118; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_119; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_120; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_121; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_122; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_123; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_124; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_125; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_126; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_127; // @[d_cache.scala 19:24]
  reg [31:0] tag_0_0; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_1; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_2; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_3; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_4; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_5; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_6; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_7; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_8; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_9; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_10; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_11; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_12; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_13; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_14; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_15; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_16; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_17; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_18; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_19; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_20; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_21; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_22; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_23; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_24; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_25; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_26; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_27; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_28; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_29; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_30; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_31; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_32; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_33; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_34; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_35; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_36; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_37; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_38; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_39; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_40; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_41; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_42; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_43; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_44; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_45; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_46; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_47; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_48; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_49; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_50; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_51; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_52; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_53; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_54; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_55; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_56; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_57; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_58; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_59; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_60; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_61; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_62; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_63; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_64; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_65; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_66; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_67; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_68; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_69; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_70; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_71; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_72; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_73; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_74; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_75; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_76; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_77; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_78; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_79; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_80; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_81; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_82; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_83; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_84; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_85; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_86; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_87; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_88; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_89; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_90; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_91; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_92; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_93; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_94; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_95; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_96; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_97; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_98; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_99; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_100; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_101; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_102; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_103; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_104; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_105; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_106; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_107; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_108; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_109; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_110; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_111; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_112; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_113; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_114; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_115; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_116; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_117; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_118; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_119; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_120; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_121; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_122; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_123; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_124; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_125; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_126; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_127; // @[d_cache.scala 20:24]
  reg [31:0] tag_1_0; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_1; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_2; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_3; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_4; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_5; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_6; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_7; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_8; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_9; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_10; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_11; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_12; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_13; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_14; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_15; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_16; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_17; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_18; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_19; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_20; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_21; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_22; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_23; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_24; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_25; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_26; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_27; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_28; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_29; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_30; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_31; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_32; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_33; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_34; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_35; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_36; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_37; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_38; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_39; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_40; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_41; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_42; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_43; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_44; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_45; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_46; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_47; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_48; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_49; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_50; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_51; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_52; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_53; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_54; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_55; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_56; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_57; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_58; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_59; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_60; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_61; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_62; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_63; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_64; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_65; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_66; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_67; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_68; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_69; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_70; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_71; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_72; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_73; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_74; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_75; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_76; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_77; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_78; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_79; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_80; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_81; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_82; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_83; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_84; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_85; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_86; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_87; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_88; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_89; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_90; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_91; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_92; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_93; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_94; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_95; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_96; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_97; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_98; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_99; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_100; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_101; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_102; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_103; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_104; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_105; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_106; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_107; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_108; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_109; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_110; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_111; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_112; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_113; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_114; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_115; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_116; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_117; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_118; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_119; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_120; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_121; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_122; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_123; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_124; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_125; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_126; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_127; // @[d_cache.scala 21:24]
  reg  valid_0_0; // @[d_cache.scala 22:26]
  reg  valid_0_1; // @[d_cache.scala 22:26]
  reg  valid_0_2; // @[d_cache.scala 22:26]
  reg  valid_0_3; // @[d_cache.scala 22:26]
  reg  valid_0_4; // @[d_cache.scala 22:26]
  reg  valid_0_5; // @[d_cache.scala 22:26]
  reg  valid_0_6; // @[d_cache.scala 22:26]
  reg  valid_0_7; // @[d_cache.scala 22:26]
  reg  valid_0_8; // @[d_cache.scala 22:26]
  reg  valid_0_9; // @[d_cache.scala 22:26]
  reg  valid_0_10; // @[d_cache.scala 22:26]
  reg  valid_0_11; // @[d_cache.scala 22:26]
  reg  valid_0_12; // @[d_cache.scala 22:26]
  reg  valid_0_13; // @[d_cache.scala 22:26]
  reg  valid_0_14; // @[d_cache.scala 22:26]
  reg  valid_0_15; // @[d_cache.scala 22:26]
  reg  valid_0_16; // @[d_cache.scala 22:26]
  reg  valid_0_17; // @[d_cache.scala 22:26]
  reg  valid_0_18; // @[d_cache.scala 22:26]
  reg  valid_0_19; // @[d_cache.scala 22:26]
  reg  valid_0_20; // @[d_cache.scala 22:26]
  reg  valid_0_21; // @[d_cache.scala 22:26]
  reg  valid_0_22; // @[d_cache.scala 22:26]
  reg  valid_0_23; // @[d_cache.scala 22:26]
  reg  valid_0_24; // @[d_cache.scala 22:26]
  reg  valid_0_25; // @[d_cache.scala 22:26]
  reg  valid_0_26; // @[d_cache.scala 22:26]
  reg  valid_0_27; // @[d_cache.scala 22:26]
  reg  valid_0_28; // @[d_cache.scala 22:26]
  reg  valid_0_29; // @[d_cache.scala 22:26]
  reg  valid_0_30; // @[d_cache.scala 22:26]
  reg  valid_0_31; // @[d_cache.scala 22:26]
  reg  valid_0_32; // @[d_cache.scala 22:26]
  reg  valid_0_33; // @[d_cache.scala 22:26]
  reg  valid_0_34; // @[d_cache.scala 22:26]
  reg  valid_0_35; // @[d_cache.scala 22:26]
  reg  valid_0_36; // @[d_cache.scala 22:26]
  reg  valid_0_37; // @[d_cache.scala 22:26]
  reg  valid_0_38; // @[d_cache.scala 22:26]
  reg  valid_0_39; // @[d_cache.scala 22:26]
  reg  valid_0_40; // @[d_cache.scala 22:26]
  reg  valid_0_41; // @[d_cache.scala 22:26]
  reg  valid_0_42; // @[d_cache.scala 22:26]
  reg  valid_0_43; // @[d_cache.scala 22:26]
  reg  valid_0_44; // @[d_cache.scala 22:26]
  reg  valid_0_45; // @[d_cache.scala 22:26]
  reg  valid_0_46; // @[d_cache.scala 22:26]
  reg  valid_0_47; // @[d_cache.scala 22:26]
  reg  valid_0_48; // @[d_cache.scala 22:26]
  reg  valid_0_49; // @[d_cache.scala 22:26]
  reg  valid_0_50; // @[d_cache.scala 22:26]
  reg  valid_0_51; // @[d_cache.scala 22:26]
  reg  valid_0_52; // @[d_cache.scala 22:26]
  reg  valid_0_53; // @[d_cache.scala 22:26]
  reg  valid_0_54; // @[d_cache.scala 22:26]
  reg  valid_0_55; // @[d_cache.scala 22:26]
  reg  valid_0_56; // @[d_cache.scala 22:26]
  reg  valid_0_57; // @[d_cache.scala 22:26]
  reg  valid_0_58; // @[d_cache.scala 22:26]
  reg  valid_0_59; // @[d_cache.scala 22:26]
  reg  valid_0_60; // @[d_cache.scala 22:26]
  reg  valid_0_61; // @[d_cache.scala 22:26]
  reg  valid_0_62; // @[d_cache.scala 22:26]
  reg  valid_0_63; // @[d_cache.scala 22:26]
  reg  valid_0_64; // @[d_cache.scala 22:26]
  reg  valid_0_65; // @[d_cache.scala 22:26]
  reg  valid_0_66; // @[d_cache.scala 22:26]
  reg  valid_0_67; // @[d_cache.scala 22:26]
  reg  valid_0_68; // @[d_cache.scala 22:26]
  reg  valid_0_69; // @[d_cache.scala 22:26]
  reg  valid_0_70; // @[d_cache.scala 22:26]
  reg  valid_0_71; // @[d_cache.scala 22:26]
  reg  valid_0_72; // @[d_cache.scala 22:26]
  reg  valid_0_73; // @[d_cache.scala 22:26]
  reg  valid_0_74; // @[d_cache.scala 22:26]
  reg  valid_0_75; // @[d_cache.scala 22:26]
  reg  valid_0_76; // @[d_cache.scala 22:26]
  reg  valid_0_77; // @[d_cache.scala 22:26]
  reg  valid_0_78; // @[d_cache.scala 22:26]
  reg  valid_0_79; // @[d_cache.scala 22:26]
  reg  valid_0_80; // @[d_cache.scala 22:26]
  reg  valid_0_81; // @[d_cache.scala 22:26]
  reg  valid_0_82; // @[d_cache.scala 22:26]
  reg  valid_0_83; // @[d_cache.scala 22:26]
  reg  valid_0_84; // @[d_cache.scala 22:26]
  reg  valid_0_85; // @[d_cache.scala 22:26]
  reg  valid_0_86; // @[d_cache.scala 22:26]
  reg  valid_0_87; // @[d_cache.scala 22:26]
  reg  valid_0_88; // @[d_cache.scala 22:26]
  reg  valid_0_89; // @[d_cache.scala 22:26]
  reg  valid_0_90; // @[d_cache.scala 22:26]
  reg  valid_0_91; // @[d_cache.scala 22:26]
  reg  valid_0_92; // @[d_cache.scala 22:26]
  reg  valid_0_93; // @[d_cache.scala 22:26]
  reg  valid_0_94; // @[d_cache.scala 22:26]
  reg  valid_0_95; // @[d_cache.scala 22:26]
  reg  valid_0_96; // @[d_cache.scala 22:26]
  reg  valid_0_97; // @[d_cache.scala 22:26]
  reg  valid_0_98; // @[d_cache.scala 22:26]
  reg  valid_0_99; // @[d_cache.scala 22:26]
  reg  valid_0_100; // @[d_cache.scala 22:26]
  reg  valid_0_101; // @[d_cache.scala 22:26]
  reg  valid_0_102; // @[d_cache.scala 22:26]
  reg  valid_0_103; // @[d_cache.scala 22:26]
  reg  valid_0_104; // @[d_cache.scala 22:26]
  reg  valid_0_105; // @[d_cache.scala 22:26]
  reg  valid_0_106; // @[d_cache.scala 22:26]
  reg  valid_0_107; // @[d_cache.scala 22:26]
  reg  valid_0_108; // @[d_cache.scala 22:26]
  reg  valid_0_109; // @[d_cache.scala 22:26]
  reg  valid_0_110; // @[d_cache.scala 22:26]
  reg  valid_0_111; // @[d_cache.scala 22:26]
  reg  valid_0_112; // @[d_cache.scala 22:26]
  reg  valid_0_113; // @[d_cache.scala 22:26]
  reg  valid_0_114; // @[d_cache.scala 22:26]
  reg  valid_0_115; // @[d_cache.scala 22:26]
  reg  valid_0_116; // @[d_cache.scala 22:26]
  reg  valid_0_117; // @[d_cache.scala 22:26]
  reg  valid_0_118; // @[d_cache.scala 22:26]
  reg  valid_0_119; // @[d_cache.scala 22:26]
  reg  valid_0_120; // @[d_cache.scala 22:26]
  reg  valid_0_121; // @[d_cache.scala 22:26]
  reg  valid_0_122; // @[d_cache.scala 22:26]
  reg  valid_0_123; // @[d_cache.scala 22:26]
  reg  valid_0_124; // @[d_cache.scala 22:26]
  reg  valid_0_125; // @[d_cache.scala 22:26]
  reg  valid_0_126; // @[d_cache.scala 22:26]
  reg  valid_0_127; // @[d_cache.scala 22:26]
  reg  valid_1_0; // @[d_cache.scala 23:26]
  reg  valid_1_1; // @[d_cache.scala 23:26]
  reg  valid_1_2; // @[d_cache.scala 23:26]
  reg  valid_1_3; // @[d_cache.scala 23:26]
  reg  valid_1_4; // @[d_cache.scala 23:26]
  reg  valid_1_5; // @[d_cache.scala 23:26]
  reg  valid_1_6; // @[d_cache.scala 23:26]
  reg  valid_1_7; // @[d_cache.scala 23:26]
  reg  valid_1_8; // @[d_cache.scala 23:26]
  reg  valid_1_9; // @[d_cache.scala 23:26]
  reg  valid_1_10; // @[d_cache.scala 23:26]
  reg  valid_1_11; // @[d_cache.scala 23:26]
  reg  valid_1_12; // @[d_cache.scala 23:26]
  reg  valid_1_13; // @[d_cache.scala 23:26]
  reg  valid_1_14; // @[d_cache.scala 23:26]
  reg  valid_1_15; // @[d_cache.scala 23:26]
  reg  valid_1_16; // @[d_cache.scala 23:26]
  reg  valid_1_17; // @[d_cache.scala 23:26]
  reg  valid_1_18; // @[d_cache.scala 23:26]
  reg  valid_1_19; // @[d_cache.scala 23:26]
  reg  valid_1_20; // @[d_cache.scala 23:26]
  reg  valid_1_21; // @[d_cache.scala 23:26]
  reg  valid_1_22; // @[d_cache.scala 23:26]
  reg  valid_1_23; // @[d_cache.scala 23:26]
  reg  valid_1_24; // @[d_cache.scala 23:26]
  reg  valid_1_25; // @[d_cache.scala 23:26]
  reg  valid_1_26; // @[d_cache.scala 23:26]
  reg  valid_1_27; // @[d_cache.scala 23:26]
  reg  valid_1_28; // @[d_cache.scala 23:26]
  reg  valid_1_29; // @[d_cache.scala 23:26]
  reg  valid_1_30; // @[d_cache.scala 23:26]
  reg  valid_1_31; // @[d_cache.scala 23:26]
  reg  valid_1_32; // @[d_cache.scala 23:26]
  reg  valid_1_33; // @[d_cache.scala 23:26]
  reg  valid_1_34; // @[d_cache.scala 23:26]
  reg  valid_1_35; // @[d_cache.scala 23:26]
  reg  valid_1_36; // @[d_cache.scala 23:26]
  reg  valid_1_37; // @[d_cache.scala 23:26]
  reg  valid_1_38; // @[d_cache.scala 23:26]
  reg  valid_1_39; // @[d_cache.scala 23:26]
  reg  valid_1_40; // @[d_cache.scala 23:26]
  reg  valid_1_41; // @[d_cache.scala 23:26]
  reg  valid_1_42; // @[d_cache.scala 23:26]
  reg  valid_1_43; // @[d_cache.scala 23:26]
  reg  valid_1_44; // @[d_cache.scala 23:26]
  reg  valid_1_45; // @[d_cache.scala 23:26]
  reg  valid_1_46; // @[d_cache.scala 23:26]
  reg  valid_1_47; // @[d_cache.scala 23:26]
  reg  valid_1_48; // @[d_cache.scala 23:26]
  reg  valid_1_49; // @[d_cache.scala 23:26]
  reg  valid_1_50; // @[d_cache.scala 23:26]
  reg  valid_1_51; // @[d_cache.scala 23:26]
  reg  valid_1_52; // @[d_cache.scala 23:26]
  reg  valid_1_53; // @[d_cache.scala 23:26]
  reg  valid_1_54; // @[d_cache.scala 23:26]
  reg  valid_1_55; // @[d_cache.scala 23:26]
  reg  valid_1_56; // @[d_cache.scala 23:26]
  reg  valid_1_57; // @[d_cache.scala 23:26]
  reg  valid_1_58; // @[d_cache.scala 23:26]
  reg  valid_1_59; // @[d_cache.scala 23:26]
  reg  valid_1_60; // @[d_cache.scala 23:26]
  reg  valid_1_61; // @[d_cache.scala 23:26]
  reg  valid_1_62; // @[d_cache.scala 23:26]
  reg  valid_1_63; // @[d_cache.scala 23:26]
  reg  valid_1_64; // @[d_cache.scala 23:26]
  reg  valid_1_65; // @[d_cache.scala 23:26]
  reg  valid_1_66; // @[d_cache.scala 23:26]
  reg  valid_1_67; // @[d_cache.scala 23:26]
  reg  valid_1_68; // @[d_cache.scala 23:26]
  reg  valid_1_69; // @[d_cache.scala 23:26]
  reg  valid_1_70; // @[d_cache.scala 23:26]
  reg  valid_1_71; // @[d_cache.scala 23:26]
  reg  valid_1_72; // @[d_cache.scala 23:26]
  reg  valid_1_73; // @[d_cache.scala 23:26]
  reg  valid_1_74; // @[d_cache.scala 23:26]
  reg  valid_1_75; // @[d_cache.scala 23:26]
  reg  valid_1_76; // @[d_cache.scala 23:26]
  reg  valid_1_77; // @[d_cache.scala 23:26]
  reg  valid_1_78; // @[d_cache.scala 23:26]
  reg  valid_1_79; // @[d_cache.scala 23:26]
  reg  valid_1_80; // @[d_cache.scala 23:26]
  reg  valid_1_81; // @[d_cache.scala 23:26]
  reg  valid_1_82; // @[d_cache.scala 23:26]
  reg  valid_1_83; // @[d_cache.scala 23:26]
  reg  valid_1_84; // @[d_cache.scala 23:26]
  reg  valid_1_85; // @[d_cache.scala 23:26]
  reg  valid_1_86; // @[d_cache.scala 23:26]
  reg  valid_1_87; // @[d_cache.scala 23:26]
  reg  valid_1_88; // @[d_cache.scala 23:26]
  reg  valid_1_89; // @[d_cache.scala 23:26]
  reg  valid_1_90; // @[d_cache.scala 23:26]
  reg  valid_1_91; // @[d_cache.scala 23:26]
  reg  valid_1_92; // @[d_cache.scala 23:26]
  reg  valid_1_93; // @[d_cache.scala 23:26]
  reg  valid_1_94; // @[d_cache.scala 23:26]
  reg  valid_1_95; // @[d_cache.scala 23:26]
  reg  valid_1_96; // @[d_cache.scala 23:26]
  reg  valid_1_97; // @[d_cache.scala 23:26]
  reg  valid_1_98; // @[d_cache.scala 23:26]
  reg  valid_1_99; // @[d_cache.scala 23:26]
  reg  valid_1_100; // @[d_cache.scala 23:26]
  reg  valid_1_101; // @[d_cache.scala 23:26]
  reg  valid_1_102; // @[d_cache.scala 23:26]
  reg  valid_1_103; // @[d_cache.scala 23:26]
  reg  valid_1_104; // @[d_cache.scala 23:26]
  reg  valid_1_105; // @[d_cache.scala 23:26]
  reg  valid_1_106; // @[d_cache.scala 23:26]
  reg  valid_1_107; // @[d_cache.scala 23:26]
  reg  valid_1_108; // @[d_cache.scala 23:26]
  reg  valid_1_109; // @[d_cache.scala 23:26]
  reg  valid_1_110; // @[d_cache.scala 23:26]
  reg  valid_1_111; // @[d_cache.scala 23:26]
  reg  valid_1_112; // @[d_cache.scala 23:26]
  reg  valid_1_113; // @[d_cache.scala 23:26]
  reg  valid_1_114; // @[d_cache.scala 23:26]
  reg  valid_1_115; // @[d_cache.scala 23:26]
  reg  valid_1_116; // @[d_cache.scala 23:26]
  reg  valid_1_117; // @[d_cache.scala 23:26]
  reg  valid_1_118; // @[d_cache.scala 23:26]
  reg  valid_1_119; // @[d_cache.scala 23:26]
  reg  valid_1_120; // @[d_cache.scala 23:26]
  reg  valid_1_121; // @[d_cache.scala 23:26]
  reg  valid_1_122; // @[d_cache.scala 23:26]
  reg  valid_1_123; // @[d_cache.scala 23:26]
  reg  valid_1_124; // @[d_cache.scala 23:26]
  reg  valid_1_125; // @[d_cache.scala 23:26]
  reg  valid_1_126; // @[d_cache.scala 23:26]
  reg  valid_1_127; // @[d_cache.scala 23:26]
  reg  dirty_0_0; // @[d_cache.scala 24:26]
  reg  dirty_0_1; // @[d_cache.scala 24:26]
  reg  dirty_0_2; // @[d_cache.scala 24:26]
  reg  dirty_0_3; // @[d_cache.scala 24:26]
  reg  dirty_0_4; // @[d_cache.scala 24:26]
  reg  dirty_0_5; // @[d_cache.scala 24:26]
  reg  dirty_0_6; // @[d_cache.scala 24:26]
  reg  dirty_0_7; // @[d_cache.scala 24:26]
  reg  dirty_0_8; // @[d_cache.scala 24:26]
  reg  dirty_0_9; // @[d_cache.scala 24:26]
  reg  dirty_0_10; // @[d_cache.scala 24:26]
  reg  dirty_0_11; // @[d_cache.scala 24:26]
  reg  dirty_0_12; // @[d_cache.scala 24:26]
  reg  dirty_0_13; // @[d_cache.scala 24:26]
  reg  dirty_0_14; // @[d_cache.scala 24:26]
  reg  dirty_0_15; // @[d_cache.scala 24:26]
  reg  dirty_0_16; // @[d_cache.scala 24:26]
  reg  dirty_0_17; // @[d_cache.scala 24:26]
  reg  dirty_0_18; // @[d_cache.scala 24:26]
  reg  dirty_0_19; // @[d_cache.scala 24:26]
  reg  dirty_0_20; // @[d_cache.scala 24:26]
  reg  dirty_0_21; // @[d_cache.scala 24:26]
  reg  dirty_0_22; // @[d_cache.scala 24:26]
  reg  dirty_0_23; // @[d_cache.scala 24:26]
  reg  dirty_0_24; // @[d_cache.scala 24:26]
  reg  dirty_0_25; // @[d_cache.scala 24:26]
  reg  dirty_0_26; // @[d_cache.scala 24:26]
  reg  dirty_0_27; // @[d_cache.scala 24:26]
  reg  dirty_0_28; // @[d_cache.scala 24:26]
  reg  dirty_0_29; // @[d_cache.scala 24:26]
  reg  dirty_0_30; // @[d_cache.scala 24:26]
  reg  dirty_0_31; // @[d_cache.scala 24:26]
  reg  dirty_0_32; // @[d_cache.scala 24:26]
  reg  dirty_0_33; // @[d_cache.scala 24:26]
  reg  dirty_0_34; // @[d_cache.scala 24:26]
  reg  dirty_0_35; // @[d_cache.scala 24:26]
  reg  dirty_0_36; // @[d_cache.scala 24:26]
  reg  dirty_0_37; // @[d_cache.scala 24:26]
  reg  dirty_0_38; // @[d_cache.scala 24:26]
  reg  dirty_0_39; // @[d_cache.scala 24:26]
  reg  dirty_0_40; // @[d_cache.scala 24:26]
  reg  dirty_0_41; // @[d_cache.scala 24:26]
  reg  dirty_0_42; // @[d_cache.scala 24:26]
  reg  dirty_0_43; // @[d_cache.scala 24:26]
  reg  dirty_0_44; // @[d_cache.scala 24:26]
  reg  dirty_0_45; // @[d_cache.scala 24:26]
  reg  dirty_0_46; // @[d_cache.scala 24:26]
  reg  dirty_0_47; // @[d_cache.scala 24:26]
  reg  dirty_0_48; // @[d_cache.scala 24:26]
  reg  dirty_0_49; // @[d_cache.scala 24:26]
  reg  dirty_0_50; // @[d_cache.scala 24:26]
  reg  dirty_0_51; // @[d_cache.scala 24:26]
  reg  dirty_0_52; // @[d_cache.scala 24:26]
  reg  dirty_0_53; // @[d_cache.scala 24:26]
  reg  dirty_0_54; // @[d_cache.scala 24:26]
  reg  dirty_0_55; // @[d_cache.scala 24:26]
  reg  dirty_0_56; // @[d_cache.scala 24:26]
  reg  dirty_0_57; // @[d_cache.scala 24:26]
  reg  dirty_0_58; // @[d_cache.scala 24:26]
  reg  dirty_0_59; // @[d_cache.scala 24:26]
  reg  dirty_0_60; // @[d_cache.scala 24:26]
  reg  dirty_0_61; // @[d_cache.scala 24:26]
  reg  dirty_0_62; // @[d_cache.scala 24:26]
  reg  dirty_0_63; // @[d_cache.scala 24:26]
  reg  dirty_0_64; // @[d_cache.scala 24:26]
  reg  dirty_0_65; // @[d_cache.scala 24:26]
  reg  dirty_0_66; // @[d_cache.scala 24:26]
  reg  dirty_0_67; // @[d_cache.scala 24:26]
  reg  dirty_0_68; // @[d_cache.scala 24:26]
  reg  dirty_0_69; // @[d_cache.scala 24:26]
  reg  dirty_0_70; // @[d_cache.scala 24:26]
  reg  dirty_0_71; // @[d_cache.scala 24:26]
  reg  dirty_0_72; // @[d_cache.scala 24:26]
  reg  dirty_0_73; // @[d_cache.scala 24:26]
  reg  dirty_0_74; // @[d_cache.scala 24:26]
  reg  dirty_0_75; // @[d_cache.scala 24:26]
  reg  dirty_0_76; // @[d_cache.scala 24:26]
  reg  dirty_0_77; // @[d_cache.scala 24:26]
  reg  dirty_0_78; // @[d_cache.scala 24:26]
  reg  dirty_0_79; // @[d_cache.scala 24:26]
  reg  dirty_0_80; // @[d_cache.scala 24:26]
  reg  dirty_0_81; // @[d_cache.scala 24:26]
  reg  dirty_0_82; // @[d_cache.scala 24:26]
  reg  dirty_0_83; // @[d_cache.scala 24:26]
  reg  dirty_0_84; // @[d_cache.scala 24:26]
  reg  dirty_0_85; // @[d_cache.scala 24:26]
  reg  dirty_0_86; // @[d_cache.scala 24:26]
  reg  dirty_0_87; // @[d_cache.scala 24:26]
  reg  dirty_0_88; // @[d_cache.scala 24:26]
  reg  dirty_0_89; // @[d_cache.scala 24:26]
  reg  dirty_0_90; // @[d_cache.scala 24:26]
  reg  dirty_0_91; // @[d_cache.scala 24:26]
  reg  dirty_0_92; // @[d_cache.scala 24:26]
  reg  dirty_0_93; // @[d_cache.scala 24:26]
  reg  dirty_0_94; // @[d_cache.scala 24:26]
  reg  dirty_0_95; // @[d_cache.scala 24:26]
  reg  dirty_0_96; // @[d_cache.scala 24:26]
  reg  dirty_0_97; // @[d_cache.scala 24:26]
  reg  dirty_0_98; // @[d_cache.scala 24:26]
  reg  dirty_0_99; // @[d_cache.scala 24:26]
  reg  dirty_0_100; // @[d_cache.scala 24:26]
  reg  dirty_0_101; // @[d_cache.scala 24:26]
  reg  dirty_0_102; // @[d_cache.scala 24:26]
  reg  dirty_0_103; // @[d_cache.scala 24:26]
  reg  dirty_0_104; // @[d_cache.scala 24:26]
  reg  dirty_0_105; // @[d_cache.scala 24:26]
  reg  dirty_0_106; // @[d_cache.scala 24:26]
  reg  dirty_0_107; // @[d_cache.scala 24:26]
  reg  dirty_0_108; // @[d_cache.scala 24:26]
  reg  dirty_0_109; // @[d_cache.scala 24:26]
  reg  dirty_0_110; // @[d_cache.scala 24:26]
  reg  dirty_0_111; // @[d_cache.scala 24:26]
  reg  dirty_0_112; // @[d_cache.scala 24:26]
  reg  dirty_0_113; // @[d_cache.scala 24:26]
  reg  dirty_0_114; // @[d_cache.scala 24:26]
  reg  dirty_0_115; // @[d_cache.scala 24:26]
  reg  dirty_0_116; // @[d_cache.scala 24:26]
  reg  dirty_0_117; // @[d_cache.scala 24:26]
  reg  dirty_0_118; // @[d_cache.scala 24:26]
  reg  dirty_0_119; // @[d_cache.scala 24:26]
  reg  dirty_0_120; // @[d_cache.scala 24:26]
  reg  dirty_0_121; // @[d_cache.scala 24:26]
  reg  dirty_0_122; // @[d_cache.scala 24:26]
  reg  dirty_0_123; // @[d_cache.scala 24:26]
  reg  dirty_0_124; // @[d_cache.scala 24:26]
  reg  dirty_0_125; // @[d_cache.scala 24:26]
  reg  dirty_0_126; // @[d_cache.scala 24:26]
  reg  dirty_0_127; // @[d_cache.scala 24:26]
  reg  dirty_1_0; // @[d_cache.scala 25:26]
  reg  dirty_1_1; // @[d_cache.scala 25:26]
  reg  dirty_1_2; // @[d_cache.scala 25:26]
  reg  dirty_1_3; // @[d_cache.scala 25:26]
  reg  dirty_1_4; // @[d_cache.scala 25:26]
  reg  dirty_1_5; // @[d_cache.scala 25:26]
  reg  dirty_1_6; // @[d_cache.scala 25:26]
  reg  dirty_1_7; // @[d_cache.scala 25:26]
  reg  dirty_1_8; // @[d_cache.scala 25:26]
  reg  dirty_1_9; // @[d_cache.scala 25:26]
  reg  dirty_1_10; // @[d_cache.scala 25:26]
  reg  dirty_1_11; // @[d_cache.scala 25:26]
  reg  dirty_1_12; // @[d_cache.scala 25:26]
  reg  dirty_1_13; // @[d_cache.scala 25:26]
  reg  dirty_1_14; // @[d_cache.scala 25:26]
  reg  dirty_1_15; // @[d_cache.scala 25:26]
  reg  dirty_1_16; // @[d_cache.scala 25:26]
  reg  dirty_1_17; // @[d_cache.scala 25:26]
  reg  dirty_1_18; // @[d_cache.scala 25:26]
  reg  dirty_1_19; // @[d_cache.scala 25:26]
  reg  dirty_1_20; // @[d_cache.scala 25:26]
  reg  dirty_1_21; // @[d_cache.scala 25:26]
  reg  dirty_1_22; // @[d_cache.scala 25:26]
  reg  dirty_1_23; // @[d_cache.scala 25:26]
  reg  dirty_1_24; // @[d_cache.scala 25:26]
  reg  dirty_1_25; // @[d_cache.scala 25:26]
  reg  dirty_1_26; // @[d_cache.scala 25:26]
  reg  dirty_1_27; // @[d_cache.scala 25:26]
  reg  dirty_1_28; // @[d_cache.scala 25:26]
  reg  dirty_1_29; // @[d_cache.scala 25:26]
  reg  dirty_1_30; // @[d_cache.scala 25:26]
  reg  dirty_1_31; // @[d_cache.scala 25:26]
  reg  dirty_1_32; // @[d_cache.scala 25:26]
  reg  dirty_1_33; // @[d_cache.scala 25:26]
  reg  dirty_1_34; // @[d_cache.scala 25:26]
  reg  dirty_1_35; // @[d_cache.scala 25:26]
  reg  dirty_1_36; // @[d_cache.scala 25:26]
  reg  dirty_1_37; // @[d_cache.scala 25:26]
  reg  dirty_1_38; // @[d_cache.scala 25:26]
  reg  dirty_1_39; // @[d_cache.scala 25:26]
  reg  dirty_1_40; // @[d_cache.scala 25:26]
  reg  dirty_1_41; // @[d_cache.scala 25:26]
  reg  dirty_1_42; // @[d_cache.scala 25:26]
  reg  dirty_1_43; // @[d_cache.scala 25:26]
  reg  dirty_1_44; // @[d_cache.scala 25:26]
  reg  dirty_1_45; // @[d_cache.scala 25:26]
  reg  dirty_1_46; // @[d_cache.scala 25:26]
  reg  dirty_1_47; // @[d_cache.scala 25:26]
  reg  dirty_1_48; // @[d_cache.scala 25:26]
  reg  dirty_1_49; // @[d_cache.scala 25:26]
  reg  dirty_1_50; // @[d_cache.scala 25:26]
  reg  dirty_1_51; // @[d_cache.scala 25:26]
  reg  dirty_1_52; // @[d_cache.scala 25:26]
  reg  dirty_1_53; // @[d_cache.scala 25:26]
  reg  dirty_1_54; // @[d_cache.scala 25:26]
  reg  dirty_1_55; // @[d_cache.scala 25:26]
  reg  dirty_1_56; // @[d_cache.scala 25:26]
  reg  dirty_1_57; // @[d_cache.scala 25:26]
  reg  dirty_1_58; // @[d_cache.scala 25:26]
  reg  dirty_1_59; // @[d_cache.scala 25:26]
  reg  dirty_1_60; // @[d_cache.scala 25:26]
  reg  dirty_1_61; // @[d_cache.scala 25:26]
  reg  dirty_1_62; // @[d_cache.scala 25:26]
  reg  dirty_1_63; // @[d_cache.scala 25:26]
  reg  dirty_1_64; // @[d_cache.scala 25:26]
  reg  dirty_1_65; // @[d_cache.scala 25:26]
  reg  dirty_1_66; // @[d_cache.scala 25:26]
  reg  dirty_1_67; // @[d_cache.scala 25:26]
  reg  dirty_1_68; // @[d_cache.scala 25:26]
  reg  dirty_1_69; // @[d_cache.scala 25:26]
  reg  dirty_1_70; // @[d_cache.scala 25:26]
  reg  dirty_1_71; // @[d_cache.scala 25:26]
  reg  dirty_1_72; // @[d_cache.scala 25:26]
  reg  dirty_1_73; // @[d_cache.scala 25:26]
  reg  dirty_1_74; // @[d_cache.scala 25:26]
  reg  dirty_1_75; // @[d_cache.scala 25:26]
  reg  dirty_1_76; // @[d_cache.scala 25:26]
  reg  dirty_1_77; // @[d_cache.scala 25:26]
  reg  dirty_1_78; // @[d_cache.scala 25:26]
  reg  dirty_1_79; // @[d_cache.scala 25:26]
  reg  dirty_1_80; // @[d_cache.scala 25:26]
  reg  dirty_1_81; // @[d_cache.scala 25:26]
  reg  dirty_1_82; // @[d_cache.scala 25:26]
  reg  dirty_1_83; // @[d_cache.scala 25:26]
  reg  dirty_1_84; // @[d_cache.scala 25:26]
  reg  dirty_1_85; // @[d_cache.scala 25:26]
  reg  dirty_1_86; // @[d_cache.scala 25:26]
  reg  dirty_1_87; // @[d_cache.scala 25:26]
  reg  dirty_1_88; // @[d_cache.scala 25:26]
  reg  dirty_1_89; // @[d_cache.scala 25:26]
  reg  dirty_1_90; // @[d_cache.scala 25:26]
  reg  dirty_1_91; // @[d_cache.scala 25:26]
  reg  dirty_1_92; // @[d_cache.scala 25:26]
  reg  dirty_1_93; // @[d_cache.scala 25:26]
  reg  dirty_1_94; // @[d_cache.scala 25:26]
  reg  dirty_1_95; // @[d_cache.scala 25:26]
  reg  dirty_1_96; // @[d_cache.scala 25:26]
  reg  dirty_1_97; // @[d_cache.scala 25:26]
  reg  dirty_1_98; // @[d_cache.scala 25:26]
  reg  dirty_1_99; // @[d_cache.scala 25:26]
  reg  dirty_1_100; // @[d_cache.scala 25:26]
  reg  dirty_1_101; // @[d_cache.scala 25:26]
  reg  dirty_1_102; // @[d_cache.scala 25:26]
  reg  dirty_1_103; // @[d_cache.scala 25:26]
  reg  dirty_1_104; // @[d_cache.scala 25:26]
  reg  dirty_1_105; // @[d_cache.scala 25:26]
  reg  dirty_1_106; // @[d_cache.scala 25:26]
  reg  dirty_1_107; // @[d_cache.scala 25:26]
  reg  dirty_1_108; // @[d_cache.scala 25:26]
  reg  dirty_1_109; // @[d_cache.scala 25:26]
  reg  dirty_1_110; // @[d_cache.scala 25:26]
  reg  dirty_1_111; // @[d_cache.scala 25:26]
  reg  dirty_1_112; // @[d_cache.scala 25:26]
  reg  dirty_1_113; // @[d_cache.scala 25:26]
  reg  dirty_1_114; // @[d_cache.scala 25:26]
  reg  dirty_1_115; // @[d_cache.scala 25:26]
  reg  dirty_1_116; // @[d_cache.scala 25:26]
  reg  dirty_1_117; // @[d_cache.scala 25:26]
  reg  dirty_1_118; // @[d_cache.scala 25:26]
  reg  dirty_1_119; // @[d_cache.scala 25:26]
  reg  dirty_1_120; // @[d_cache.scala 25:26]
  reg  dirty_1_121; // @[d_cache.scala 25:26]
  reg  dirty_1_122; // @[d_cache.scala 25:26]
  reg  dirty_1_123; // @[d_cache.scala 25:26]
  reg  dirty_1_124; // @[d_cache.scala 25:26]
  reg  dirty_1_125; // @[d_cache.scala 25:26]
  reg  dirty_1_126; // @[d_cache.scala 25:26]
  reg  dirty_1_127; // @[d_cache.scala 25:26]
  reg  way0_hit; // @[d_cache.scala 26:27]
  reg  way1_hit; // @[d_cache.scala 27:27]
  reg [63:0] write_back_data; // @[d_cache.scala 29:34]
  reg [31:0] write_back_addr; // @[d_cache.scala 30:34]
  reg [1:0] unuse_way; // @[d_cache.scala 33:28]
  reg [63:0] receive_data; // @[d_cache.scala 34:31]
  reg  quene; // @[d_cache.scala 35:24]
  wire [6:0] index = io_from_lsu_araddr[6:0]; // @[d_cache.scala 38:35]
  wire [24:0] tag = io_from_lsu_araddr[31:7]; // @[d_cache.scala 39:33]
  wire [31:0] _GEN_1 = 7'h1 == index ? tag_0_1 : tag_0_0; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_2 = 7'h2 == index ? tag_0_2 : _GEN_1; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_3 = 7'h3 == index ? tag_0_3 : _GEN_2; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_4 = 7'h4 == index ? tag_0_4 : _GEN_3; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_5 = 7'h5 == index ? tag_0_5 : _GEN_4; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_6 = 7'h6 == index ? tag_0_6 : _GEN_5; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_7 = 7'h7 == index ? tag_0_7 : _GEN_6; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_8 = 7'h8 == index ? tag_0_8 : _GEN_7; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_9 = 7'h9 == index ? tag_0_9 : _GEN_8; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_10 = 7'ha == index ? tag_0_10 : _GEN_9; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_11 = 7'hb == index ? tag_0_11 : _GEN_10; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_12 = 7'hc == index ? tag_0_12 : _GEN_11; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_13 = 7'hd == index ? tag_0_13 : _GEN_12; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_14 = 7'he == index ? tag_0_14 : _GEN_13; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_15 = 7'hf == index ? tag_0_15 : _GEN_14; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_16 = 7'h10 == index ? tag_0_16 : _GEN_15; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_17 = 7'h11 == index ? tag_0_17 : _GEN_16; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_18 = 7'h12 == index ? tag_0_18 : _GEN_17; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_19 = 7'h13 == index ? tag_0_19 : _GEN_18; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_20 = 7'h14 == index ? tag_0_20 : _GEN_19; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_21 = 7'h15 == index ? tag_0_21 : _GEN_20; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_22 = 7'h16 == index ? tag_0_22 : _GEN_21; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_23 = 7'h17 == index ? tag_0_23 : _GEN_22; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_24 = 7'h18 == index ? tag_0_24 : _GEN_23; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_25 = 7'h19 == index ? tag_0_25 : _GEN_24; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_26 = 7'h1a == index ? tag_0_26 : _GEN_25; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_27 = 7'h1b == index ? tag_0_27 : _GEN_26; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_28 = 7'h1c == index ? tag_0_28 : _GEN_27; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_29 = 7'h1d == index ? tag_0_29 : _GEN_28; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_30 = 7'h1e == index ? tag_0_30 : _GEN_29; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_31 = 7'h1f == index ? tag_0_31 : _GEN_30; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_32 = 7'h20 == index ? tag_0_32 : _GEN_31; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_33 = 7'h21 == index ? tag_0_33 : _GEN_32; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_34 = 7'h22 == index ? tag_0_34 : _GEN_33; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_35 = 7'h23 == index ? tag_0_35 : _GEN_34; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_36 = 7'h24 == index ? tag_0_36 : _GEN_35; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_37 = 7'h25 == index ? tag_0_37 : _GEN_36; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_38 = 7'h26 == index ? tag_0_38 : _GEN_37; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_39 = 7'h27 == index ? tag_0_39 : _GEN_38; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_40 = 7'h28 == index ? tag_0_40 : _GEN_39; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_41 = 7'h29 == index ? tag_0_41 : _GEN_40; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_42 = 7'h2a == index ? tag_0_42 : _GEN_41; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_43 = 7'h2b == index ? tag_0_43 : _GEN_42; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_44 = 7'h2c == index ? tag_0_44 : _GEN_43; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_45 = 7'h2d == index ? tag_0_45 : _GEN_44; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_46 = 7'h2e == index ? tag_0_46 : _GEN_45; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_47 = 7'h2f == index ? tag_0_47 : _GEN_46; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_48 = 7'h30 == index ? tag_0_48 : _GEN_47; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_49 = 7'h31 == index ? tag_0_49 : _GEN_48; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_50 = 7'h32 == index ? tag_0_50 : _GEN_49; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_51 = 7'h33 == index ? tag_0_51 : _GEN_50; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_52 = 7'h34 == index ? tag_0_52 : _GEN_51; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_53 = 7'h35 == index ? tag_0_53 : _GEN_52; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_54 = 7'h36 == index ? tag_0_54 : _GEN_53; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_55 = 7'h37 == index ? tag_0_55 : _GEN_54; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_56 = 7'h38 == index ? tag_0_56 : _GEN_55; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_57 = 7'h39 == index ? tag_0_57 : _GEN_56; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_58 = 7'h3a == index ? tag_0_58 : _GEN_57; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_59 = 7'h3b == index ? tag_0_59 : _GEN_58; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_60 = 7'h3c == index ? tag_0_60 : _GEN_59; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_61 = 7'h3d == index ? tag_0_61 : _GEN_60; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_62 = 7'h3e == index ? tag_0_62 : _GEN_61; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_63 = 7'h3f == index ? tag_0_63 : _GEN_62; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_64 = 7'h40 == index ? tag_0_64 : _GEN_63; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_65 = 7'h41 == index ? tag_0_65 : _GEN_64; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_66 = 7'h42 == index ? tag_0_66 : _GEN_65; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_67 = 7'h43 == index ? tag_0_67 : _GEN_66; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_68 = 7'h44 == index ? tag_0_68 : _GEN_67; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_69 = 7'h45 == index ? tag_0_69 : _GEN_68; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_70 = 7'h46 == index ? tag_0_70 : _GEN_69; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_71 = 7'h47 == index ? tag_0_71 : _GEN_70; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_72 = 7'h48 == index ? tag_0_72 : _GEN_71; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_73 = 7'h49 == index ? tag_0_73 : _GEN_72; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_74 = 7'h4a == index ? tag_0_74 : _GEN_73; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_75 = 7'h4b == index ? tag_0_75 : _GEN_74; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_76 = 7'h4c == index ? tag_0_76 : _GEN_75; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_77 = 7'h4d == index ? tag_0_77 : _GEN_76; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_78 = 7'h4e == index ? tag_0_78 : _GEN_77; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_79 = 7'h4f == index ? tag_0_79 : _GEN_78; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_80 = 7'h50 == index ? tag_0_80 : _GEN_79; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_81 = 7'h51 == index ? tag_0_81 : _GEN_80; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_82 = 7'h52 == index ? tag_0_82 : _GEN_81; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_83 = 7'h53 == index ? tag_0_83 : _GEN_82; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_84 = 7'h54 == index ? tag_0_84 : _GEN_83; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_85 = 7'h55 == index ? tag_0_85 : _GEN_84; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_86 = 7'h56 == index ? tag_0_86 : _GEN_85; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_87 = 7'h57 == index ? tag_0_87 : _GEN_86; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_88 = 7'h58 == index ? tag_0_88 : _GEN_87; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_89 = 7'h59 == index ? tag_0_89 : _GEN_88; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_90 = 7'h5a == index ? tag_0_90 : _GEN_89; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_91 = 7'h5b == index ? tag_0_91 : _GEN_90; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_92 = 7'h5c == index ? tag_0_92 : _GEN_91; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_93 = 7'h5d == index ? tag_0_93 : _GEN_92; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_94 = 7'h5e == index ? tag_0_94 : _GEN_93; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_95 = 7'h5f == index ? tag_0_95 : _GEN_94; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_96 = 7'h60 == index ? tag_0_96 : _GEN_95; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_97 = 7'h61 == index ? tag_0_97 : _GEN_96; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_98 = 7'h62 == index ? tag_0_98 : _GEN_97; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_99 = 7'h63 == index ? tag_0_99 : _GEN_98; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_100 = 7'h64 == index ? tag_0_100 : _GEN_99; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_101 = 7'h65 == index ? tag_0_101 : _GEN_100; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_102 = 7'h66 == index ? tag_0_102 : _GEN_101; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_103 = 7'h67 == index ? tag_0_103 : _GEN_102; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_104 = 7'h68 == index ? tag_0_104 : _GEN_103; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_105 = 7'h69 == index ? tag_0_105 : _GEN_104; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_106 = 7'h6a == index ? tag_0_106 : _GEN_105; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_107 = 7'h6b == index ? tag_0_107 : _GEN_106; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_108 = 7'h6c == index ? tag_0_108 : _GEN_107; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_109 = 7'h6d == index ? tag_0_109 : _GEN_108; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_110 = 7'h6e == index ? tag_0_110 : _GEN_109; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_111 = 7'h6f == index ? tag_0_111 : _GEN_110; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_112 = 7'h70 == index ? tag_0_112 : _GEN_111; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_113 = 7'h71 == index ? tag_0_113 : _GEN_112; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_114 = 7'h72 == index ? tag_0_114 : _GEN_113; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_115 = 7'h73 == index ? tag_0_115 : _GEN_114; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_116 = 7'h74 == index ? tag_0_116 : _GEN_115; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_117 = 7'h75 == index ? tag_0_117 : _GEN_116; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_118 = 7'h76 == index ? tag_0_118 : _GEN_117; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_119 = 7'h77 == index ? tag_0_119 : _GEN_118; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_120 = 7'h78 == index ? tag_0_120 : _GEN_119; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_121 = 7'h79 == index ? tag_0_121 : _GEN_120; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_122 = 7'h7a == index ? tag_0_122 : _GEN_121; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_123 = 7'h7b == index ? tag_0_123 : _GEN_122; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_124 = 7'h7c == index ? tag_0_124 : _GEN_123; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_125 = 7'h7d == index ? tag_0_125 : _GEN_124; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_126 = 7'h7e == index ? tag_0_126 : _GEN_125; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_127 = 7'h7f == index ? tag_0_127 : _GEN_126; // @[d_cache.scala 41:{24,24}]
  wire [31:0] _GEN_15265 = {{7'd0}, tag}; // @[d_cache.scala 41:24]
  wire  _GEN_129 = 7'h1 == index ? valid_0_1 : valid_0_0; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_130 = 7'h2 == index ? valid_0_2 : _GEN_129; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_131 = 7'h3 == index ? valid_0_3 : _GEN_130; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_132 = 7'h4 == index ? valid_0_4 : _GEN_131; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_133 = 7'h5 == index ? valid_0_5 : _GEN_132; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_134 = 7'h6 == index ? valid_0_6 : _GEN_133; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_135 = 7'h7 == index ? valid_0_7 : _GEN_134; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_136 = 7'h8 == index ? valid_0_8 : _GEN_135; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_137 = 7'h9 == index ? valid_0_9 : _GEN_136; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_138 = 7'ha == index ? valid_0_10 : _GEN_137; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_139 = 7'hb == index ? valid_0_11 : _GEN_138; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_140 = 7'hc == index ? valid_0_12 : _GEN_139; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_141 = 7'hd == index ? valid_0_13 : _GEN_140; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_142 = 7'he == index ? valid_0_14 : _GEN_141; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_143 = 7'hf == index ? valid_0_15 : _GEN_142; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_144 = 7'h10 == index ? valid_0_16 : _GEN_143; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_145 = 7'h11 == index ? valid_0_17 : _GEN_144; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_146 = 7'h12 == index ? valid_0_18 : _GEN_145; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_147 = 7'h13 == index ? valid_0_19 : _GEN_146; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_148 = 7'h14 == index ? valid_0_20 : _GEN_147; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_149 = 7'h15 == index ? valid_0_21 : _GEN_148; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_150 = 7'h16 == index ? valid_0_22 : _GEN_149; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_151 = 7'h17 == index ? valid_0_23 : _GEN_150; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_152 = 7'h18 == index ? valid_0_24 : _GEN_151; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_153 = 7'h19 == index ? valid_0_25 : _GEN_152; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_154 = 7'h1a == index ? valid_0_26 : _GEN_153; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_155 = 7'h1b == index ? valid_0_27 : _GEN_154; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_156 = 7'h1c == index ? valid_0_28 : _GEN_155; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_157 = 7'h1d == index ? valid_0_29 : _GEN_156; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_158 = 7'h1e == index ? valid_0_30 : _GEN_157; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_159 = 7'h1f == index ? valid_0_31 : _GEN_158; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_160 = 7'h20 == index ? valid_0_32 : _GEN_159; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_161 = 7'h21 == index ? valid_0_33 : _GEN_160; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_162 = 7'h22 == index ? valid_0_34 : _GEN_161; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_163 = 7'h23 == index ? valid_0_35 : _GEN_162; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_164 = 7'h24 == index ? valid_0_36 : _GEN_163; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_165 = 7'h25 == index ? valid_0_37 : _GEN_164; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_166 = 7'h26 == index ? valid_0_38 : _GEN_165; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_167 = 7'h27 == index ? valid_0_39 : _GEN_166; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_168 = 7'h28 == index ? valid_0_40 : _GEN_167; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_169 = 7'h29 == index ? valid_0_41 : _GEN_168; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_170 = 7'h2a == index ? valid_0_42 : _GEN_169; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_171 = 7'h2b == index ? valid_0_43 : _GEN_170; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_172 = 7'h2c == index ? valid_0_44 : _GEN_171; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_173 = 7'h2d == index ? valid_0_45 : _GEN_172; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_174 = 7'h2e == index ? valid_0_46 : _GEN_173; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_175 = 7'h2f == index ? valid_0_47 : _GEN_174; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_176 = 7'h30 == index ? valid_0_48 : _GEN_175; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_177 = 7'h31 == index ? valid_0_49 : _GEN_176; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_178 = 7'h32 == index ? valid_0_50 : _GEN_177; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_179 = 7'h33 == index ? valid_0_51 : _GEN_178; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_180 = 7'h34 == index ? valid_0_52 : _GEN_179; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_181 = 7'h35 == index ? valid_0_53 : _GEN_180; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_182 = 7'h36 == index ? valid_0_54 : _GEN_181; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_183 = 7'h37 == index ? valid_0_55 : _GEN_182; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_184 = 7'h38 == index ? valid_0_56 : _GEN_183; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_185 = 7'h39 == index ? valid_0_57 : _GEN_184; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_186 = 7'h3a == index ? valid_0_58 : _GEN_185; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_187 = 7'h3b == index ? valid_0_59 : _GEN_186; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_188 = 7'h3c == index ? valid_0_60 : _GEN_187; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_189 = 7'h3d == index ? valid_0_61 : _GEN_188; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_190 = 7'h3e == index ? valid_0_62 : _GEN_189; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_191 = 7'h3f == index ? valid_0_63 : _GEN_190; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_192 = 7'h40 == index ? valid_0_64 : _GEN_191; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_193 = 7'h41 == index ? valid_0_65 : _GEN_192; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_194 = 7'h42 == index ? valid_0_66 : _GEN_193; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_195 = 7'h43 == index ? valid_0_67 : _GEN_194; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_196 = 7'h44 == index ? valid_0_68 : _GEN_195; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_197 = 7'h45 == index ? valid_0_69 : _GEN_196; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_198 = 7'h46 == index ? valid_0_70 : _GEN_197; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_199 = 7'h47 == index ? valid_0_71 : _GEN_198; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_200 = 7'h48 == index ? valid_0_72 : _GEN_199; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_201 = 7'h49 == index ? valid_0_73 : _GEN_200; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_202 = 7'h4a == index ? valid_0_74 : _GEN_201; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_203 = 7'h4b == index ? valid_0_75 : _GEN_202; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_204 = 7'h4c == index ? valid_0_76 : _GEN_203; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_205 = 7'h4d == index ? valid_0_77 : _GEN_204; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_206 = 7'h4e == index ? valid_0_78 : _GEN_205; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_207 = 7'h4f == index ? valid_0_79 : _GEN_206; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_208 = 7'h50 == index ? valid_0_80 : _GEN_207; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_209 = 7'h51 == index ? valid_0_81 : _GEN_208; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_210 = 7'h52 == index ? valid_0_82 : _GEN_209; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_211 = 7'h53 == index ? valid_0_83 : _GEN_210; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_212 = 7'h54 == index ? valid_0_84 : _GEN_211; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_213 = 7'h55 == index ? valid_0_85 : _GEN_212; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_214 = 7'h56 == index ? valid_0_86 : _GEN_213; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_215 = 7'h57 == index ? valid_0_87 : _GEN_214; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_216 = 7'h58 == index ? valid_0_88 : _GEN_215; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_217 = 7'h59 == index ? valid_0_89 : _GEN_216; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_218 = 7'h5a == index ? valid_0_90 : _GEN_217; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_219 = 7'h5b == index ? valid_0_91 : _GEN_218; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_220 = 7'h5c == index ? valid_0_92 : _GEN_219; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_221 = 7'h5d == index ? valid_0_93 : _GEN_220; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_222 = 7'h5e == index ? valid_0_94 : _GEN_221; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_223 = 7'h5f == index ? valid_0_95 : _GEN_222; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_224 = 7'h60 == index ? valid_0_96 : _GEN_223; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_225 = 7'h61 == index ? valid_0_97 : _GEN_224; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_226 = 7'h62 == index ? valid_0_98 : _GEN_225; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_227 = 7'h63 == index ? valid_0_99 : _GEN_226; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_228 = 7'h64 == index ? valid_0_100 : _GEN_227; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_229 = 7'h65 == index ? valid_0_101 : _GEN_228; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_230 = 7'h66 == index ? valid_0_102 : _GEN_229; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_231 = 7'h67 == index ? valid_0_103 : _GEN_230; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_232 = 7'h68 == index ? valid_0_104 : _GEN_231; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_233 = 7'h69 == index ? valid_0_105 : _GEN_232; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_234 = 7'h6a == index ? valid_0_106 : _GEN_233; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_235 = 7'h6b == index ? valid_0_107 : _GEN_234; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_236 = 7'h6c == index ? valid_0_108 : _GEN_235; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_237 = 7'h6d == index ? valid_0_109 : _GEN_236; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_238 = 7'h6e == index ? valid_0_110 : _GEN_237; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_239 = 7'h6f == index ? valid_0_111 : _GEN_238; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_240 = 7'h70 == index ? valid_0_112 : _GEN_239; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_241 = 7'h71 == index ? valid_0_113 : _GEN_240; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_242 = 7'h72 == index ? valid_0_114 : _GEN_241; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_243 = 7'h73 == index ? valid_0_115 : _GEN_242; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_244 = 7'h74 == index ? valid_0_116 : _GEN_243; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_245 = 7'h75 == index ? valid_0_117 : _GEN_244; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_246 = 7'h76 == index ? valid_0_118 : _GEN_245; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_247 = 7'h77 == index ? valid_0_119 : _GEN_246; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_248 = 7'h78 == index ? valid_0_120 : _GEN_247; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_249 = 7'h79 == index ? valid_0_121 : _GEN_248; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_250 = 7'h7a == index ? valid_0_122 : _GEN_249; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_251 = 7'h7b == index ? valid_0_123 : _GEN_250; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_252 = 7'h7c == index ? valid_0_124 : _GEN_251; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_253 = 7'h7d == index ? valid_0_125 : _GEN_252; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_254 = 7'h7e == index ? valid_0_126 : _GEN_253; // @[d_cache.scala 41:{50,50}]
  wire  _GEN_255 = 7'h7f == index ? valid_0_127 : _GEN_254; // @[d_cache.scala 41:{50,50}]
  wire  _T_4 = _GEN_127 == _GEN_15265 & _GEN_255; // @[d_cache.scala 41:33]
  wire [31:0] _GEN_258 = 7'h1 == index ? tag_1_1 : tag_1_0; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_259 = 7'h2 == index ? tag_1_2 : _GEN_258; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_260 = 7'h3 == index ? tag_1_3 : _GEN_259; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_261 = 7'h4 == index ? tag_1_4 : _GEN_260; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_262 = 7'h5 == index ? tag_1_5 : _GEN_261; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_263 = 7'h6 == index ? tag_1_6 : _GEN_262; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_264 = 7'h7 == index ? tag_1_7 : _GEN_263; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_265 = 7'h8 == index ? tag_1_8 : _GEN_264; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_266 = 7'h9 == index ? tag_1_9 : _GEN_265; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_267 = 7'ha == index ? tag_1_10 : _GEN_266; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_268 = 7'hb == index ? tag_1_11 : _GEN_267; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_269 = 7'hc == index ? tag_1_12 : _GEN_268; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_270 = 7'hd == index ? tag_1_13 : _GEN_269; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_271 = 7'he == index ? tag_1_14 : _GEN_270; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_272 = 7'hf == index ? tag_1_15 : _GEN_271; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_273 = 7'h10 == index ? tag_1_16 : _GEN_272; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_274 = 7'h11 == index ? tag_1_17 : _GEN_273; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_275 = 7'h12 == index ? tag_1_18 : _GEN_274; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_276 = 7'h13 == index ? tag_1_19 : _GEN_275; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_277 = 7'h14 == index ? tag_1_20 : _GEN_276; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_278 = 7'h15 == index ? tag_1_21 : _GEN_277; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_279 = 7'h16 == index ? tag_1_22 : _GEN_278; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_280 = 7'h17 == index ? tag_1_23 : _GEN_279; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_281 = 7'h18 == index ? tag_1_24 : _GEN_280; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_282 = 7'h19 == index ? tag_1_25 : _GEN_281; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_283 = 7'h1a == index ? tag_1_26 : _GEN_282; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_284 = 7'h1b == index ? tag_1_27 : _GEN_283; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_285 = 7'h1c == index ? tag_1_28 : _GEN_284; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_286 = 7'h1d == index ? tag_1_29 : _GEN_285; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_287 = 7'h1e == index ? tag_1_30 : _GEN_286; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_288 = 7'h1f == index ? tag_1_31 : _GEN_287; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_289 = 7'h20 == index ? tag_1_32 : _GEN_288; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_290 = 7'h21 == index ? tag_1_33 : _GEN_289; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_291 = 7'h22 == index ? tag_1_34 : _GEN_290; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_292 = 7'h23 == index ? tag_1_35 : _GEN_291; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_293 = 7'h24 == index ? tag_1_36 : _GEN_292; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_294 = 7'h25 == index ? tag_1_37 : _GEN_293; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_295 = 7'h26 == index ? tag_1_38 : _GEN_294; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_296 = 7'h27 == index ? tag_1_39 : _GEN_295; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_297 = 7'h28 == index ? tag_1_40 : _GEN_296; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_298 = 7'h29 == index ? tag_1_41 : _GEN_297; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_299 = 7'h2a == index ? tag_1_42 : _GEN_298; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_300 = 7'h2b == index ? tag_1_43 : _GEN_299; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_301 = 7'h2c == index ? tag_1_44 : _GEN_300; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_302 = 7'h2d == index ? tag_1_45 : _GEN_301; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_303 = 7'h2e == index ? tag_1_46 : _GEN_302; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_304 = 7'h2f == index ? tag_1_47 : _GEN_303; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_305 = 7'h30 == index ? tag_1_48 : _GEN_304; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_306 = 7'h31 == index ? tag_1_49 : _GEN_305; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_307 = 7'h32 == index ? tag_1_50 : _GEN_306; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_308 = 7'h33 == index ? tag_1_51 : _GEN_307; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_309 = 7'h34 == index ? tag_1_52 : _GEN_308; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_310 = 7'h35 == index ? tag_1_53 : _GEN_309; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_311 = 7'h36 == index ? tag_1_54 : _GEN_310; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_312 = 7'h37 == index ? tag_1_55 : _GEN_311; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_313 = 7'h38 == index ? tag_1_56 : _GEN_312; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_314 = 7'h39 == index ? tag_1_57 : _GEN_313; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_315 = 7'h3a == index ? tag_1_58 : _GEN_314; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_316 = 7'h3b == index ? tag_1_59 : _GEN_315; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_317 = 7'h3c == index ? tag_1_60 : _GEN_316; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_318 = 7'h3d == index ? tag_1_61 : _GEN_317; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_319 = 7'h3e == index ? tag_1_62 : _GEN_318; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_320 = 7'h3f == index ? tag_1_63 : _GEN_319; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_321 = 7'h40 == index ? tag_1_64 : _GEN_320; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_322 = 7'h41 == index ? tag_1_65 : _GEN_321; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_323 = 7'h42 == index ? tag_1_66 : _GEN_322; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_324 = 7'h43 == index ? tag_1_67 : _GEN_323; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_325 = 7'h44 == index ? tag_1_68 : _GEN_324; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_326 = 7'h45 == index ? tag_1_69 : _GEN_325; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_327 = 7'h46 == index ? tag_1_70 : _GEN_326; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_328 = 7'h47 == index ? tag_1_71 : _GEN_327; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_329 = 7'h48 == index ? tag_1_72 : _GEN_328; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_330 = 7'h49 == index ? tag_1_73 : _GEN_329; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_331 = 7'h4a == index ? tag_1_74 : _GEN_330; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_332 = 7'h4b == index ? tag_1_75 : _GEN_331; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_333 = 7'h4c == index ? tag_1_76 : _GEN_332; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_334 = 7'h4d == index ? tag_1_77 : _GEN_333; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_335 = 7'h4e == index ? tag_1_78 : _GEN_334; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_336 = 7'h4f == index ? tag_1_79 : _GEN_335; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_337 = 7'h50 == index ? tag_1_80 : _GEN_336; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_338 = 7'h51 == index ? tag_1_81 : _GEN_337; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_339 = 7'h52 == index ? tag_1_82 : _GEN_338; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_340 = 7'h53 == index ? tag_1_83 : _GEN_339; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_341 = 7'h54 == index ? tag_1_84 : _GEN_340; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_342 = 7'h55 == index ? tag_1_85 : _GEN_341; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_343 = 7'h56 == index ? tag_1_86 : _GEN_342; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_344 = 7'h57 == index ? tag_1_87 : _GEN_343; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_345 = 7'h58 == index ? tag_1_88 : _GEN_344; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_346 = 7'h59 == index ? tag_1_89 : _GEN_345; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_347 = 7'h5a == index ? tag_1_90 : _GEN_346; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_348 = 7'h5b == index ? tag_1_91 : _GEN_347; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_349 = 7'h5c == index ? tag_1_92 : _GEN_348; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_350 = 7'h5d == index ? tag_1_93 : _GEN_349; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_351 = 7'h5e == index ? tag_1_94 : _GEN_350; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_352 = 7'h5f == index ? tag_1_95 : _GEN_351; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_353 = 7'h60 == index ? tag_1_96 : _GEN_352; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_354 = 7'h61 == index ? tag_1_97 : _GEN_353; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_355 = 7'h62 == index ? tag_1_98 : _GEN_354; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_356 = 7'h63 == index ? tag_1_99 : _GEN_355; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_357 = 7'h64 == index ? tag_1_100 : _GEN_356; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_358 = 7'h65 == index ? tag_1_101 : _GEN_357; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_359 = 7'h66 == index ? tag_1_102 : _GEN_358; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_360 = 7'h67 == index ? tag_1_103 : _GEN_359; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_361 = 7'h68 == index ? tag_1_104 : _GEN_360; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_362 = 7'h69 == index ? tag_1_105 : _GEN_361; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_363 = 7'h6a == index ? tag_1_106 : _GEN_362; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_364 = 7'h6b == index ? tag_1_107 : _GEN_363; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_365 = 7'h6c == index ? tag_1_108 : _GEN_364; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_366 = 7'h6d == index ? tag_1_109 : _GEN_365; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_367 = 7'h6e == index ? tag_1_110 : _GEN_366; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_368 = 7'h6f == index ? tag_1_111 : _GEN_367; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_369 = 7'h70 == index ? tag_1_112 : _GEN_368; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_370 = 7'h71 == index ? tag_1_113 : _GEN_369; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_371 = 7'h72 == index ? tag_1_114 : _GEN_370; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_372 = 7'h73 == index ? tag_1_115 : _GEN_371; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_373 = 7'h74 == index ? tag_1_116 : _GEN_372; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_374 = 7'h75 == index ? tag_1_117 : _GEN_373; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_375 = 7'h76 == index ? tag_1_118 : _GEN_374; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_376 = 7'h77 == index ? tag_1_119 : _GEN_375; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_377 = 7'h78 == index ? tag_1_120 : _GEN_376; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_378 = 7'h79 == index ? tag_1_121 : _GEN_377; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_379 = 7'h7a == index ? tag_1_122 : _GEN_378; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_380 = 7'h7b == index ? tag_1_123 : _GEN_379; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_381 = 7'h7c == index ? tag_1_124 : _GEN_380; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_382 = 7'h7d == index ? tag_1_125 : _GEN_381; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_383 = 7'h7e == index ? tag_1_126 : _GEN_382; // @[d_cache.scala 46:{24,24}]
  wire [31:0] _GEN_384 = 7'h7f == index ? tag_1_127 : _GEN_383; // @[d_cache.scala 46:{24,24}]
  wire  _GEN_386 = 7'h1 == index ? valid_1_1 : valid_1_0; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_387 = 7'h2 == index ? valid_1_2 : _GEN_386; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_388 = 7'h3 == index ? valid_1_3 : _GEN_387; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_389 = 7'h4 == index ? valid_1_4 : _GEN_388; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_390 = 7'h5 == index ? valid_1_5 : _GEN_389; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_391 = 7'h6 == index ? valid_1_6 : _GEN_390; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_392 = 7'h7 == index ? valid_1_7 : _GEN_391; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_393 = 7'h8 == index ? valid_1_8 : _GEN_392; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_394 = 7'h9 == index ? valid_1_9 : _GEN_393; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_395 = 7'ha == index ? valid_1_10 : _GEN_394; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_396 = 7'hb == index ? valid_1_11 : _GEN_395; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_397 = 7'hc == index ? valid_1_12 : _GEN_396; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_398 = 7'hd == index ? valid_1_13 : _GEN_397; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_399 = 7'he == index ? valid_1_14 : _GEN_398; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_400 = 7'hf == index ? valid_1_15 : _GEN_399; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_401 = 7'h10 == index ? valid_1_16 : _GEN_400; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_402 = 7'h11 == index ? valid_1_17 : _GEN_401; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_403 = 7'h12 == index ? valid_1_18 : _GEN_402; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_404 = 7'h13 == index ? valid_1_19 : _GEN_403; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_405 = 7'h14 == index ? valid_1_20 : _GEN_404; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_406 = 7'h15 == index ? valid_1_21 : _GEN_405; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_407 = 7'h16 == index ? valid_1_22 : _GEN_406; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_408 = 7'h17 == index ? valid_1_23 : _GEN_407; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_409 = 7'h18 == index ? valid_1_24 : _GEN_408; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_410 = 7'h19 == index ? valid_1_25 : _GEN_409; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_411 = 7'h1a == index ? valid_1_26 : _GEN_410; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_412 = 7'h1b == index ? valid_1_27 : _GEN_411; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_413 = 7'h1c == index ? valid_1_28 : _GEN_412; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_414 = 7'h1d == index ? valid_1_29 : _GEN_413; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_415 = 7'h1e == index ? valid_1_30 : _GEN_414; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_416 = 7'h1f == index ? valid_1_31 : _GEN_415; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_417 = 7'h20 == index ? valid_1_32 : _GEN_416; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_418 = 7'h21 == index ? valid_1_33 : _GEN_417; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_419 = 7'h22 == index ? valid_1_34 : _GEN_418; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_420 = 7'h23 == index ? valid_1_35 : _GEN_419; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_421 = 7'h24 == index ? valid_1_36 : _GEN_420; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_422 = 7'h25 == index ? valid_1_37 : _GEN_421; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_423 = 7'h26 == index ? valid_1_38 : _GEN_422; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_424 = 7'h27 == index ? valid_1_39 : _GEN_423; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_425 = 7'h28 == index ? valid_1_40 : _GEN_424; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_426 = 7'h29 == index ? valid_1_41 : _GEN_425; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_427 = 7'h2a == index ? valid_1_42 : _GEN_426; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_428 = 7'h2b == index ? valid_1_43 : _GEN_427; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_429 = 7'h2c == index ? valid_1_44 : _GEN_428; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_430 = 7'h2d == index ? valid_1_45 : _GEN_429; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_431 = 7'h2e == index ? valid_1_46 : _GEN_430; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_432 = 7'h2f == index ? valid_1_47 : _GEN_431; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_433 = 7'h30 == index ? valid_1_48 : _GEN_432; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_434 = 7'h31 == index ? valid_1_49 : _GEN_433; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_435 = 7'h32 == index ? valid_1_50 : _GEN_434; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_436 = 7'h33 == index ? valid_1_51 : _GEN_435; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_437 = 7'h34 == index ? valid_1_52 : _GEN_436; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_438 = 7'h35 == index ? valid_1_53 : _GEN_437; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_439 = 7'h36 == index ? valid_1_54 : _GEN_438; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_440 = 7'h37 == index ? valid_1_55 : _GEN_439; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_441 = 7'h38 == index ? valid_1_56 : _GEN_440; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_442 = 7'h39 == index ? valid_1_57 : _GEN_441; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_443 = 7'h3a == index ? valid_1_58 : _GEN_442; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_444 = 7'h3b == index ? valid_1_59 : _GEN_443; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_445 = 7'h3c == index ? valid_1_60 : _GEN_444; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_446 = 7'h3d == index ? valid_1_61 : _GEN_445; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_447 = 7'h3e == index ? valid_1_62 : _GEN_446; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_448 = 7'h3f == index ? valid_1_63 : _GEN_447; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_449 = 7'h40 == index ? valid_1_64 : _GEN_448; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_450 = 7'h41 == index ? valid_1_65 : _GEN_449; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_451 = 7'h42 == index ? valid_1_66 : _GEN_450; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_452 = 7'h43 == index ? valid_1_67 : _GEN_451; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_453 = 7'h44 == index ? valid_1_68 : _GEN_452; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_454 = 7'h45 == index ? valid_1_69 : _GEN_453; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_455 = 7'h46 == index ? valid_1_70 : _GEN_454; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_456 = 7'h47 == index ? valid_1_71 : _GEN_455; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_457 = 7'h48 == index ? valid_1_72 : _GEN_456; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_458 = 7'h49 == index ? valid_1_73 : _GEN_457; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_459 = 7'h4a == index ? valid_1_74 : _GEN_458; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_460 = 7'h4b == index ? valid_1_75 : _GEN_459; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_461 = 7'h4c == index ? valid_1_76 : _GEN_460; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_462 = 7'h4d == index ? valid_1_77 : _GEN_461; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_463 = 7'h4e == index ? valid_1_78 : _GEN_462; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_464 = 7'h4f == index ? valid_1_79 : _GEN_463; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_465 = 7'h50 == index ? valid_1_80 : _GEN_464; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_466 = 7'h51 == index ? valid_1_81 : _GEN_465; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_467 = 7'h52 == index ? valid_1_82 : _GEN_466; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_468 = 7'h53 == index ? valid_1_83 : _GEN_467; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_469 = 7'h54 == index ? valid_1_84 : _GEN_468; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_470 = 7'h55 == index ? valid_1_85 : _GEN_469; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_471 = 7'h56 == index ? valid_1_86 : _GEN_470; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_472 = 7'h57 == index ? valid_1_87 : _GEN_471; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_473 = 7'h58 == index ? valid_1_88 : _GEN_472; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_474 = 7'h59 == index ? valid_1_89 : _GEN_473; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_475 = 7'h5a == index ? valid_1_90 : _GEN_474; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_476 = 7'h5b == index ? valid_1_91 : _GEN_475; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_477 = 7'h5c == index ? valid_1_92 : _GEN_476; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_478 = 7'h5d == index ? valid_1_93 : _GEN_477; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_479 = 7'h5e == index ? valid_1_94 : _GEN_478; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_480 = 7'h5f == index ? valid_1_95 : _GEN_479; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_481 = 7'h60 == index ? valid_1_96 : _GEN_480; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_482 = 7'h61 == index ? valid_1_97 : _GEN_481; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_483 = 7'h62 == index ? valid_1_98 : _GEN_482; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_484 = 7'h63 == index ? valid_1_99 : _GEN_483; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_485 = 7'h64 == index ? valid_1_100 : _GEN_484; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_486 = 7'h65 == index ? valid_1_101 : _GEN_485; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_487 = 7'h66 == index ? valid_1_102 : _GEN_486; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_488 = 7'h67 == index ? valid_1_103 : _GEN_487; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_489 = 7'h68 == index ? valid_1_104 : _GEN_488; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_490 = 7'h69 == index ? valid_1_105 : _GEN_489; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_491 = 7'h6a == index ? valid_1_106 : _GEN_490; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_492 = 7'h6b == index ? valid_1_107 : _GEN_491; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_493 = 7'h6c == index ? valid_1_108 : _GEN_492; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_494 = 7'h6d == index ? valid_1_109 : _GEN_493; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_495 = 7'h6e == index ? valid_1_110 : _GEN_494; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_496 = 7'h6f == index ? valid_1_111 : _GEN_495; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_497 = 7'h70 == index ? valid_1_112 : _GEN_496; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_498 = 7'h71 == index ? valid_1_113 : _GEN_497; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_499 = 7'h72 == index ? valid_1_114 : _GEN_498; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_500 = 7'h73 == index ? valid_1_115 : _GEN_499; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_501 = 7'h74 == index ? valid_1_116 : _GEN_500; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_502 = 7'h75 == index ? valid_1_117 : _GEN_501; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_503 = 7'h76 == index ? valid_1_118 : _GEN_502; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_504 = 7'h77 == index ? valid_1_119 : _GEN_503; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_505 = 7'h78 == index ? valid_1_120 : _GEN_504; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_506 = 7'h79 == index ? valid_1_121 : _GEN_505; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_507 = 7'h7a == index ? valid_1_122 : _GEN_506; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_508 = 7'h7b == index ? valid_1_123 : _GEN_507; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_509 = 7'h7c == index ? valid_1_124 : _GEN_508; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_510 = 7'h7d == index ? valid_1_125 : _GEN_509; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_511 = 7'h7e == index ? valid_1_126 : _GEN_510; // @[d_cache.scala 46:{50,50}]
  wire  _GEN_512 = 7'h7f == index ? valid_1_127 : _GEN_511; // @[d_cache.scala 46:{50,50}]
  wire  _T_7 = _GEN_384 == _GEN_15265 & _GEN_512; // @[d_cache.scala 46:33]
  reg [2:0] state; // @[d_cache.scala 60:24]
  wire  _T_16 = 3'h0 == state; // @[d_cache.scala 64:18]
  wire  _T_17 = 3'h1 == state; // @[d_cache.scala 64:18]
  wire  _GEN_519 = 7'h1 == index ? dirty_0_1 : dirty_0_0; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_520 = 7'h2 == index ? dirty_0_2 : _GEN_519; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_521 = 7'h3 == index ? dirty_0_3 : _GEN_520; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_522 = 7'h4 == index ? dirty_0_4 : _GEN_521; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_523 = 7'h5 == index ? dirty_0_5 : _GEN_522; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_524 = 7'h6 == index ? dirty_0_6 : _GEN_523; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_525 = 7'h7 == index ? dirty_0_7 : _GEN_524; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_526 = 7'h8 == index ? dirty_0_8 : _GEN_525; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_527 = 7'h9 == index ? dirty_0_9 : _GEN_526; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_528 = 7'ha == index ? dirty_0_10 : _GEN_527; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_529 = 7'hb == index ? dirty_0_11 : _GEN_528; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_530 = 7'hc == index ? dirty_0_12 : _GEN_529; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_531 = 7'hd == index ? dirty_0_13 : _GEN_530; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_532 = 7'he == index ? dirty_0_14 : _GEN_531; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_533 = 7'hf == index ? dirty_0_15 : _GEN_532; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_534 = 7'h10 == index ? dirty_0_16 : _GEN_533; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_535 = 7'h11 == index ? dirty_0_17 : _GEN_534; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_536 = 7'h12 == index ? dirty_0_18 : _GEN_535; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_537 = 7'h13 == index ? dirty_0_19 : _GEN_536; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_538 = 7'h14 == index ? dirty_0_20 : _GEN_537; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_539 = 7'h15 == index ? dirty_0_21 : _GEN_538; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_540 = 7'h16 == index ? dirty_0_22 : _GEN_539; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_541 = 7'h17 == index ? dirty_0_23 : _GEN_540; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_542 = 7'h18 == index ? dirty_0_24 : _GEN_541; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_543 = 7'h19 == index ? dirty_0_25 : _GEN_542; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_544 = 7'h1a == index ? dirty_0_26 : _GEN_543; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_545 = 7'h1b == index ? dirty_0_27 : _GEN_544; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_546 = 7'h1c == index ? dirty_0_28 : _GEN_545; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_547 = 7'h1d == index ? dirty_0_29 : _GEN_546; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_548 = 7'h1e == index ? dirty_0_30 : _GEN_547; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_549 = 7'h1f == index ? dirty_0_31 : _GEN_548; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_550 = 7'h20 == index ? dirty_0_32 : _GEN_549; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_551 = 7'h21 == index ? dirty_0_33 : _GEN_550; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_552 = 7'h22 == index ? dirty_0_34 : _GEN_551; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_553 = 7'h23 == index ? dirty_0_35 : _GEN_552; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_554 = 7'h24 == index ? dirty_0_36 : _GEN_553; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_555 = 7'h25 == index ? dirty_0_37 : _GEN_554; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_556 = 7'h26 == index ? dirty_0_38 : _GEN_555; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_557 = 7'h27 == index ? dirty_0_39 : _GEN_556; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_558 = 7'h28 == index ? dirty_0_40 : _GEN_557; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_559 = 7'h29 == index ? dirty_0_41 : _GEN_558; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_560 = 7'h2a == index ? dirty_0_42 : _GEN_559; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_561 = 7'h2b == index ? dirty_0_43 : _GEN_560; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_562 = 7'h2c == index ? dirty_0_44 : _GEN_561; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_563 = 7'h2d == index ? dirty_0_45 : _GEN_562; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_564 = 7'h2e == index ? dirty_0_46 : _GEN_563; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_565 = 7'h2f == index ? dirty_0_47 : _GEN_564; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_566 = 7'h30 == index ? dirty_0_48 : _GEN_565; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_567 = 7'h31 == index ? dirty_0_49 : _GEN_566; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_568 = 7'h32 == index ? dirty_0_50 : _GEN_567; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_569 = 7'h33 == index ? dirty_0_51 : _GEN_568; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_570 = 7'h34 == index ? dirty_0_52 : _GEN_569; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_571 = 7'h35 == index ? dirty_0_53 : _GEN_570; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_572 = 7'h36 == index ? dirty_0_54 : _GEN_571; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_573 = 7'h37 == index ? dirty_0_55 : _GEN_572; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_574 = 7'h38 == index ? dirty_0_56 : _GEN_573; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_575 = 7'h39 == index ? dirty_0_57 : _GEN_574; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_576 = 7'h3a == index ? dirty_0_58 : _GEN_575; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_577 = 7'h3b == index ? dirty_0_59 : _GEN_576; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_578 = 7'h3c == index ? dirty_0_60 : _GEN_577; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_579 = 7'h3d == index ? dirty_0_61 : _GEN_578; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_580 = 7'h3e == index ? dirty_0_62 : _GEN_579; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_581 = 7'h3f == index ? dirty_0_63 : _GEN_580; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_582 = 7'h40 == index ? dirty_0_64 : _GEN_581; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_583 = 7'h41 == index ? dirty_0_65 : _GEN_582; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_584 = 7'h42 == index ? dirty_0_66 : _GEN_583; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_585 = 7'h43 == index ? dirty_0_67 : _GEN_584; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_586 = 7'h44 == index ? dirty_0_68 : _GEN_585; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_587 = 7'h45 == index ? dirty_0_69 : _GEN_586; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_588 = 7'h46 == index ? dirty_0_70 : _GEN_587; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_589 = 7'h47 == index ? dirty_0_71 : _GEN_588; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_590 = 7'h48 == index ? dirty_0_72 : _GEN_589; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_591 = 7'h49 == index ? dirty_0_73 : _GEN_590; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_592 = 7'h4a == index ? dirty_0_74 : _GEN_591; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_593 = 7'h4b == index ? dirty_0_75 : _GEN_592; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_594 = 7'h4c == index ? dirty_0_76 : _GEN_593; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_595 = 7'h4d == index ? dirty_0_77 : _GEN_594; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_596 = 7'h4e == index ? dirty_0_78 : _GEN_595; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_597 = 7'h4f == index ? dirty_0_79 : _GEN_596; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_598 = 7'h50 == index ? dirty_0_80 : _GEN_597; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_599 = 7'h51 == index ? dirty_0_81 : _GEN_598; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_600 = 7'h52 == index ? dirty_0_82 : _GEN_599; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_601 = 7'h53 == index ? dirty_0_83 : _GEN_600; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_602 = 7'h54 == index ? dirty_0_84 : _GEN_601; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_603 = 7'h55 == index ? dirty_0_85 : _GEN_602; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_604 = 7'h56 == index ? dirty_0_86 : _GEN_603; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_605 = 7'h57 == index ? dirty_0_87 : _GEN_604; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_606 = 7'h58 == index ? dirty_0_88 : _GEN_605; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_607 = 7'h59 == index ? dirty_0_89 : _GEN_606; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_608 = 7'h5a == index ? dirty_0_90 : _GEN_607; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_609 = 7'h5b == index ? dirty_0_91 : _GEN_608; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_610 = 7'h5c == index ? dirty_0_92 : _GEN_609; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_611 = 7'h5d == index ? dirty_0_93 : _GEN_610; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_612 = 7'h5e == index ? dirty_0_94 : _GEN_611; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_613 = 7'h5f == index ? dirty_0_95 : _GEN_612; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_614 = 7'h60 == index ? dirty_0_96 : _GEN_613; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_615 = 7'h61 == index ? dirty_0_97 : _GEN_614; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_616 = 7'h62 == index ? dirty_0_98 : _GEN_615; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_617 = 7'h63 == index ? dirty_0_99 : _GEN_616; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_618 = 7'h64 == index ? dirty_0_100 : _GEN_617; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_619 = 7'h65 == index ? dirty_0_101 : _GEN_618; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_620 = 7'h66 == index ? dirty_0_102 : _GEN_619; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_621 = 7'h67 == index ? dirty_0_103 : _GEN_620; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_622 = 7'h68 == index ? dirty_0_104 : _GEN_621; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_623 = 7'h69 == index ? dirty_0_105 : _GEN_622; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_624 = 7'h6a == index ? dirty_0_106 : _GEN_623; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_625 = 7'h6b == index ? dirty_0_107 : _GEN_624; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_626 = 7'h6c == index ? dirty_0_108 : _GEN_625; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_627 = 7'h6d == index ? dirty_0_109 : _GEN_626; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_628 = 7'h6e == index ? dirty_0_110 : _GEN_627; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_629 = 7'h6f == index ? dirty_0_111 : _GEN_628; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_630 = 7'h70 == index ? dirty_0_112 : _GEN_629; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_631 = 7'h71 == index ? dirty_0_113 : _GEN_630; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_632 = 7'h72 == index ? dirty_0_114 : _GEN_631; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_633 = 7'h73 == index ? dirty_0_115 : _GEN_632; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_634 = 7'h74 == index ? dirty_0_116 : _GEN_633; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_635 = 7'h75 == index ? dirty_0_117 : _GEN_634; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_636 = 7'h76 == index ? dirty_0_118 : _GEN_635; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_637 = 7'h77 == index ? dirty_0_119 : _GEN_636; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_638 = 7'h78 == index ? dirty_0_120 : _GEN_637; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_639 = 7'h79 == index ? dirty_0_121 : _GEN_638; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_640 = 7'h7a == index ? dirty_0_122 : _GEN_639; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_641 = 7'h7b == index ? dirty_0_123 : _GEN_640; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_642 = 7'h7c == index ? dirty_0_124 : _GEN_641; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_643 = 7'h7d == index ? dirty_0_125 : _GEN_642; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_644 = 7'h7e == index ? dirty_0_126 : _GEN_643; // @[d_cache.scala 76:{27,27}]
  wire  _GEN_645 = 7'h7f == index ? dirty_0_127 : _GEN_644; // @[d_cache.scala 76:{27,27}]
  wire [2:0] _GEN_646 = io_from_lsu_rready ? 3'h0 : state; // @[d_cache.scala 60:24 75:41 77:27]
  wire  _GEN_648 = 7'h1 == index ? dirty_1_1 : dirty_1_0; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_649 = 7'h2 == index ? dirty_1_2 : _GEN_648; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_650 = 7'h3 == index ? dirty_1_3 : _GEN_649; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_651 = 7'h4 == index ? dirty_1_4 : _GEN_650; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_652 = 7'h5 == index ? dirty_1_5 : _GEN_651; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_653 = 7'h6 == index ? dirty_1_6 : _GEN_652; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_654 = 7'h7 == index ? dirty_1_7 : _GEN_653; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_655 = 7'h8 == index ? dirty_1_8 : _GEN_654; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_656 = 7'h9 == index ? dirty_1_9 : _GEN_655; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_657 = 7'ha == index ? dirty_1_10 : _GEN_656; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_658 = 7'hb == index ? dirty_1_11 : _GEN_657; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_659 = 7'hc == index ? dirty_1_12 : _GEN_658; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_660 = 7'hd == index ? dirty_1_13 : _GEN_659; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_661 = 7'he == index ? dirty_1_14 : _GEN_660; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_662 = 7'hf == index ? dirty_1_15 : _GEN_661; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_663 = 7'h10 == index ? dirty_1_16 : _GEN_662; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_664 = 7'h11 == index ? dirty_1_17 : _GEN_663; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_665 = 7'h12 == index ? dirty_1_18 : _GEN_664; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_666 = 7'h13 == index ? dirty_1_19 : _GEN_665; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_667 = 7'h14 == index ? dirty_1_20 : _GEN_666; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_668 = 7'h15 == index ? dirty_1_21 : _GEN_667; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_669 = 7'h16 == index ? dirty_1_22 : _GEN_668; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_670 = 7'h17 == index ? dirty_1_23 : _GEN_669; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_671 = 7'h18 == index ? dirty_1_24 : _GEN_670; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_672 = 7'h19 == index ? dirty_1_25 : _GEN_671; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_673 = 7'h1a == index ? dirty_1_26 : _GEN_672; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_674 = 7'h1b == index ? dirty_1_27 : _GEN_673; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_675 = 7'h1c == index ? dirty_1_28 : _GEN_674; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_676 = 7'h1d == index ? dirty_1_29 : _GEN_675; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_677 = 7'h1e == index ? dirty_1_30 : _GEN_676; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_678 = 7'h1f == index ? dirty_1_31 : _GEN_677; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_679 = 7'h20 == index ? dirty_1_32 : _GEN_678; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_680 = 7'h21 == index ? dirty_1_33 : _GEN_679; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_681 = 7'h22 == index ? dirty_1_34 : _GEN_680; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_682 = 7'h23 == index ? dirty_1_35 : _GEN_681; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_683 = 7'h24 == index ? dirty_1_36 : _GEN_682; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_684 = 7'h25 == index ? dirty_1_37 : _GEN_683; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_685 = 7'h26 == index ? dirty_1_38 : _GEN_684; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_686 = 7'h27 == index ? dirty_1_39 : _GEN_685; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_687 = 7'h28 == index ? dirty_1_40 : _GEN_686; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_688 = 7'h29 == index ? dirty_1_41 : _GEN_687; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_689 = 7'h2a == index ? dirty_1_42 : _GEN_688; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_690 = 7'h2b == index ? dirty_1_43 : _GEN_689; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_691 = 7'h2c == index ? dirty_1_44 : _GEN_690; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_692 = 7'h2d == index ? dirty_1_45 : _GEN_691; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_693 = 7'h2e == index ? dirty_1_46 : _GEN_692; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_694 = 7'h2f == index ? dirty_1_47 : _GEN_693; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_695 = 7'h30 == index ? dirty_1_48 : _GEN_694; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_696 = 7'h31 == index ? dirty_1_49 : _GEN_695; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_697 = 7'h32 == index ? dirty_1_50 : _GEN_696; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_698 = 7'h33 == index ? dirty_1_51 : _GEN_697; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_699 = 7'h34 == index ? dirty_1_52 : _GEN_698; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_700 = 7'h35 == index ? dirty_1_53 : _GEN_699; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_701 = 7'h36 == index ? dirty_1_54 : _GEN_700; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_702 = 7'h37 == index ? dirty_1_55 : _GEN_701; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_703 = 7'h38 == index ? dirty_1_56 : _GEN_702; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_704 = 7'h39 == index ? dirty_1_57 : _GEN_703; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_705 = 7'h3a == index ? dirty_1_58 : _GEN_704; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_706 = 7'h3b == index ? dirty_1_59 : _GEN_705; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_707 = 7'h3c == index ? dirty_1_60 : _GEN_706; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_708 = 7'h3d == index ? dirty_1_61 : _GEN_707; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_709 = 7'h3e == index ? dirty_1_62 : _GEN_708; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_710 = 7'h3f == index ? dirty_1_63 : _GEN_709; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_711 = 7'h40 == index ? dirty_1_64 : _GEN_710; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_712 = 7'h41 == index ? dirty_1_65 : _GEN_711; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_713 = 7'h42 == index ? dirty_1_66 : _GEN_712; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_714 = 7'h43 == index ? dirty_1_67 : _GEN_713; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_715 = 7'h44 == index ? dirty_1_68 : _GEN_714; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_716 = 7'h45 == index ? dirty_1_69 : _GEN_715; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_717 = 7'h46 == index ? dirty_1_70 : _GEN_716; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_718 = 7'h47 == index ? dirty_1_71 : _GEN_717; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_719 = 7'h48 == index ? dirty_1_72 : _GEN_718; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_720 = 7'h49 == index ? dirty_1_73 : _GEN_719; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_721 = 7'h4a == index ? dirty_1_74 : _GEN_720; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_722 = 7'h4b == index ? dirty_1_75 : _GEN_721; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_723 = 7'h4c == index ? dirty_1_76 : _GEN_722; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_724 = 7'h4d == index ? dirty_1_77 : _GEN_723; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_725 = 7'h4e == index ? dirty_1_78 : _GEN_724; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_726 = 7'h4f == index ? dirty_1_79 : _GEN_725; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_727 = 7'h50 == index ? dirty_1_80 : _GEN_726; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_728 = 7'h51 == index ? dirty_1_81 : _GEN_727; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_729 = 7'h52 == index ? dirty_1_82 : _GEN_728; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_730 = 7'h53 == index ? dirty_1_83 : _GEN_729; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_731 = 7'h54 == index ? dirty_1_84 : _GEN_730; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_732 = 7'h55 == index ? dirty_1_85 : _GEN_731; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_733 = 7'h56 == index ? dirty_1_86 : _GEN_732; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_734 = 7'h57 == index ? dirty_1_87 : _GEN_733; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_735 = 7'h58 == index ? dirty_1_88 : _GEN_734; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_736 = 7'h59 == index ? dirty_1_89 : _GEN_735; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_737 = 7'h5a == index ? dirty_1_90 : _GEN_736; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_738 = 7'h5b == index ? dirty_1_91 : _GEN_737; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_739 = 7'h5c == index ? dirty_1_92 : _GEN_738; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_740 = 7'h5d == index ? dirty_1_93 : _GEN_739; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_741 = 7'h5e == index ? dirty_1_94 : _GEN_740; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_742 = 7'h5f == index ? dirty_1_95 : _GEN_741; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_743 = 7'h60 == index ? dirty_1_96 : _GEN_742; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_744 = 7'h61 == index ? dirty_1_97 : _GEN_743; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_745 = 7'h62 == index ? dirty_1_98 : _GEN_744; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_746 = 7'h63 == index ? dirty_1_99 : _GEN_745; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_747 = 7'h64 == index ? dirty_1_100 : _GEN_746; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_748 = 7'h65 == index ? dirty_1_101 : _GEN_747; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_749 = 7'h66 == index ? dirty_1_102 : _GEN_748; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_750 = 7'h67 == index ? dirty_1_103 : _GEN_749; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_751 = 7'h68 == index ? dirty_1_104 : _GEN_750; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_752 = 7'h69 == index ? dirty_1_105 : _GEN_751; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_753 = 7'h6a == index ? dirty_1_106 : _GEN_752; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_754 = 7'h6b == index ? dirty_1_107 : _GEN_753; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_755 = 7'h6c == index ? dirty_1_108 : _GEN_754; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_756 = 7'h6d == index ? dirty_1_109 : _GEN_755; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_757 = 7'h6e == index ? dirty_1_110 : _GEN_756; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_758 = 7'h6f == index ? dirty_1_111 : _GEN_757; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_759 = 7'h70 == index ? dirty_1_112 : _GEN_758; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_760 = 7'h71 == index ? dirty_1_113 : _GEN_759; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_761 = 7'h72 == index ? dirty_1_114 : _GEN_760; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_762 = 7'h73 == index ? dirty_1_115 : _GEN_761; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_763 = 7'h74 == index ? dirty_1_116 : _GEN_762; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_764 = 7'h75 == index ? dirty_1_117 : _GEN_763; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_765 = 7'h76 == index ? dirty_1_118 : _GEN_764; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_766 = 7'h77 == index ? dirty_1_119 : _GEN_765; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_767 = 7'h78 == index ? dirty_1_120 : _GEN_766; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_768 = 7'h79 == index ? dirty_1_121 : _GEN_767; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_769 = 7'h7a == index ? dirty_1_122 : _GEN_768; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_770 = 7'h7b == index ? dirty_1_123 : _GEN_769; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_771 = 7'h7c == index ? dirty_1_124 : _GEN_770; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_772 = 7'h7d == index ? dirty_1_125 : _GEN_771; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_773 = 7'h7e == index ? dirty_1_126 : _GEN_772; // @[d_cache.scala 82:{27,27}]
  wire  _GEN_774 = 7'h7f == index ? dirty_1_127 : _GEN_773; // @[d_cache.scala 82:{27,27}]
  wire [2:0] _GEN_775 = way1_hit ? _GEN_646 : 3'h3; // @[d_cache.scala 80:33 86:23]
  wire [63:0] _ram_0_index = {{32'd0}, io_from_lsu_wdata}; // @[d_cache.scala 92:{30,30}]
  wire [63:0] _GEN_777 = 7'h0 == index ? _ram_0_index : ram_0_0; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_778 = 7'h1 == index ? _ram_0_index : ram_0_1; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_779 = 7'h2 == index ? _ram_0_index : ram_0_2; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_780 = 7'h3 == index ? _ram_0_index : ram_0_3; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_781 = 7'h4 == index ? _ram_0_index : ram_0_4; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_782 = 7'h5 == index ? _ram_0_index : ram_0_5; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_783 = 7'h6 == index ? _ram_0_index : ram_0_6; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_784 = 7'h7 == index ? _ram_0_index : ram_0_7; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_785 = 7'h8 == index ? _ram_0_index : ram_0_8; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_786 = 7'h9 == index ? _ram_0_index : ram_0_9; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_787 = 7'ha == index ? _ram_0_index : ram_0_10; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_788 = 7'hb == index ? _ram_0_index : ram_0_11; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_789 = 7'hc == index ? _ram_0_index : ram_0_12; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_790 = 7'hd == index ? _ram_0_index : ram_0_13; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_791 = 7'he == index ? _ram_0_index : ram_0_14; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_792 = 7'hf == index ? _ram_0_index : ram_0_15; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_793 = 7'h10 == index ? _ram_0_index : ram_0_16; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_794 = 7'h11 == index ? _ram_0_index : ram_0_17; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_795 = 7'h12 == index ? _ram_0_index : ram_0_18; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_796 = 7'h13 == index ? _ram_0_index : ram_0_19; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_797 = 7'h14 == index ? _ram_0_index : ram_0_20; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_798 = 7'h15 == index ? _ram_0_index : ram_0_21; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_799 = 7'h16 == index ? _ram_0_index : ram_0_22; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_800 = 7'h17 == index ? _ram_0_index : ram_0_23; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_801 = 7'h18 == index ? _ram_0_index : ram_0_24; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_802 = 7'h19 == index ? _ram_0_index : ram_0_25; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_803 = 7'h1a == index ? _ram_0_index : ram_0_26; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_804 = 7'h1b == index ? _ram_0_index : ram_0_27; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_805 = 7'h1c == index ? _ram_0_index : ram_0_28; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_806 = 7'h1d == index ? _ram_0_index : ram_0_29; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_807 = 7'h1e == index ? _ram_0_index : ram_0_30; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_808 = 7'h1f == index ? _ram_0_index : ram_0_31; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_809 = 7'h20 == index ? _ram_0_index : ram_0_32; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_810 = 7'h21 == index ? _ram_0_index : ram_0_33; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_811 = 7'h22 == index ? _ram_0_index : ram_0_34; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_812 = 7'h23 == index ? _ram_0_index : ram_0_35; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_813 = 7'h24 == index ? _ram_0_index : ram_0_36; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_814 = 7'h25 == index ? _ram_0_index : ram_0_37; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_815 = 7'h26 == index ? _ram_0_index : ram_0_38; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_816 = 7'h27 == index ? _ram_0_index : ram_0_39; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_817 = 7'h28 == index ? _ram_0_index : ram_0_40; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_818 = 7'h29 == index ? _ram_0_index : ram_0_41; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_819 = 7'h2a == index ? _ram_0_index : ram_0_42; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_820 = 7'h2b == index ? _ram_0_index : ram_0_43; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_821 = 7'h2c == index ? _ram_0_index : ram_0_44; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_822 = 7'h2d == index ? _ram_0_index : ram_0_45; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_823 = 7'h2e == index ? _ram_0_index : ram_0_46; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_824 = 7'h2f == index ? _ram_0_index : ram_0_47; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_825 = 7'h30 == index ? _ram_0_index : ram_0_48; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_826 = 7'h31 == index ? _ram_0_index : ram_0_49; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_827 = 7'h32 == index ? _ram_0_index : ram_0_50; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_828 = 7'h33 == index ? _ram_0_index : ram_0_51; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_829 = 7'h34 == index ? _ram_0_index : ram_0_52; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_830 = 7'h35 == index ? _ram_0_index : ram_0_53; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_831 = 7'h36 == index ? _ram_0_index : ram_0_54; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_832 = 7'h37 == index ? _ram_0_index : ram_0_55; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_833 = 7'h38 == index ? _ram_0_index : ram_0_56; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_834 = 7'h39 == index ? _ram_0_index : ram_0_57; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_835 = 7'h3a == index ? _ram_0_index : ram_0_58; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_836 = 7'h3b == index ? _ram_0_index : ram_0_59; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_837 = 7'h3c == index ? _ram_0_index : ram_0_60; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_838 = 7'h3d == index ? _ram_0_index : ram_0_61; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_839 = 7'h3e == index ? _ram_0_index : ram_0_62; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_840 = 7'h3f == index ? _ram_0_index : ram_0_63; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_841 = 7'h40 == index ? _ram_0_index : ram_0_64; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_842 = 7'h41 == index ? _ram_0_index : ram_0_65; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_843 = 7'h42 == index ? _ram_0_index : ram_0_66; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_844 = 7'h43 == index ? _ram_0_index : ram_0_67; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_845 = 7'h44 == index ? _ram_0_index : ram_0_68; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_846 = 7'h45 == index ? _ram_0_index : ram_0_69; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_847 = 7'h46 == index ? _ram_0_index : ram_0_70; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_848 = 7'h47 == index ? _ram_0_index : ram_0_71; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_849 = 7'h48 == index ? _ram_0_index : ram_0_72; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_850 = 7'h49 == index ? _ram_0_index : ram_0_73; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_851 = 7'h4a == index ? _ram_0_index : ram_0_74; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_852 = 7'h4b == index ? _ram_0_index : ram_0_75; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_853 = 7'h4c == index ? _ram_0_index : ram_0_76; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_854 = 7'h4d == index ? _ram_0_index : ram_0_77; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_855 = 7'h4e == index ? _ram_0_index : ram_0_78; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_856 = 7'h4f == index ? _ram_0_index : ram_0_79; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_857 = 7'h50 == index ? _ram_0_index : ram_0_80; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_858 = 7'h51 == index ? _ram_0_index : ram_0_81; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_859 = 7'h52 == index ? _ram_0_index : ram_0_82; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_860 = 7'h53 == index ? _ram_0_index : ram_0_83; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_861 = 7'h54 == index ? _ram_0_index : ram_0_84; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_862 = 7'h55 == index ? _ram_0_index : ram_0_85; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_863 = 7'h56 == index ? _ram_0_index : ram_0_86; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_864 = 7'h57 == index ? _ram_0_index : ram_0_87; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_865 = 7'h58 == index ? _ram_0_index : ram_0_88; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_866 = 7'h59 == index ? _ram_0_index : ram_0_89; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_867 = 7'h5a == index ? _ram_0_index : ram_0_90; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_868 = 7'h5b == index ? _ram_0_index : ram_0_91; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_869 = 7'h5c == index ? _ram_0_index : ram_0_92; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_870 = 7'h5d == index ? _ram_0_index : ram_0_93; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_871 = 7'h5e == index ? _ram_0_index : ram_0_94; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_872 = 7'h5f == index ? _ram_0_index : ram_0_95; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_873 = 7'h60 == index ? _ram_0_index : ram_0_96; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_874 = 7'h61 == index ? _ram_0_index : ram_0_97; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_875 = 7'h62 == index ? _ram_0_index : ram_0_98; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_876 = 7'h63 == index ? _ram_0_index : ram_0_99; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_877 = 7'h64 == index ? _ram_0_index : ram_0_100; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_878 = 7'h65 == index ? _ram_0_index : ram_0_101; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_879 = 7'h66 == index ? _ram_0_index : ram_0_102; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_880 = 7'h67 == index ? _ram_0_index : ram_0_103; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_881 = 7'h68 == index ? _ram_0_index : ram_0_104; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_882 = 7'h69 == index ? _ram_0_index : ram_0_105; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_883 = 7'h6a == index ? _ram_0_index : ram_0_106; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_884 = 7'h6b == index ? _ram_0_index : ram_0_107; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_885 = 7'h6c == index ? _ram_0_index : ram_0_108; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_886 = 7'h6d == index ? _ram_0_index : ram_0_109; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_887 = 7'h6e == index ? _ram_0_index : ram_0_110; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_888 = 7'h6f == index ? _ram_0_index : ram_0_111; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_889 = 7'h70 == index ? _ram_0_index : ram_0_112; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_890 = 7'h71 == index ? _ram_0_index : ram_0_113; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_891 = 7'h72 == index ? _ram_0_index : ram_0_114; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_892 = 7'h73 == index ? _ram_0_index : ram_0_115; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_893 = 7'h74 == index ? _ram_0_index : ram_0_116; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_894 = 7'h75 == index ? _ram_0_index : ram_0_117; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_895 = 7'h76 == index ? _ram_0_index : ram_0_118; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_896 = 7'h77 == index ? _ram_0_index : ram_0_119; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_897 = 7'h78 == index ? _ram_0_index : ram_0_120; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_898 = 7'h79 == index ? _ram_0_index : ram_0_121; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_899 = 7'h7a == index ? _ram_0_index : ram_0_122; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_900 = 7'h7b == index ? _ram_0_index : ram_0_123; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_901 = 7'h7c == index ? _ram_0_index : ram_0_124; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_902 = 7'h7d == index ? _ram_0_index : ram_0_125; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_903 = 7'h7e == index ? _ram_0_index : ram_0_126; // @[d_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_904 = 7'h7f == index ? _ram_0_index : ram_0_127; // @[d_cache.scala 18:24 92:{30,30}]
  wire  _GEN_15267 = 7'h0 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_905 = 7'h0 == index | dirty_0_0; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15268 = 7'h1 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_906 = 7'h1 == index | dirty_0_1; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15269 = 7'h2 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_907 = 7'h2 == index | dirty_0_2; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15270 = 7'h3 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_908 = 7'h3 == index | dirty_0_3; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15271 = 7'h4 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_909 = 7'h4 == index | dirty_0_4; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15272 = 7'h5 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_910 = 7'h5 == index | dirty_0_5; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15273 = 7'h6 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_911 = 7'h6 == index | dirty_0_6; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15274 = 7'h7 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_912 = 7'h7 == index | dirty_0_7; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15275 = 7'h8 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_913 = 7'h8 == index | dirty_0_8; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15276 = 7'h9 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_914 = 7'h9 == index | dirty_0_9; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15277 = 7'ha == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_915 = 7'ha == index | dirty_0_10; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15278 = 7'hb == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_916 = 7'hb == index | dirty_0_11; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15279 = 7'hc == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_917 = 7'hc == index | dirty_0_12; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15280 = 7'hd == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_918 = 7'hd == index | dirty_0_13; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15281 = 7'he == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_919 = 7'he == index | dirty_0_14; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15282 = 7'hf == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_920 = 7'hf == index | dirty_0_15; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15283 = 7'h10 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_921 = 7'h10 == index | dirty_0_16; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15284 = 7'h11 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_922 = 7'h11 == index | dirty_0_17; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15285 = 7'h12 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_923 = 7'h12 == index | dirty_0_18; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15286 = 7'h13 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_924 = 7'h13 == index | dirty_0_19; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15287 = 7'h14 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_925 = 7'h14 == index | dirty_0_20; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15288 = 7'h15 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_926 = 7'h15 == index | dirty_0_21; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15289 = 7'h16 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_927 = 7'h16 == index | dirty_0_22; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15290 = 7'h17 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_928 = 7'h17 == index | dirty_0_23; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15291 = 7'h18 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_929 = 7'h18 == index | dirty_0_24; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15292 = 7'h19 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_930 = 7'h19 == index | dirty_0_25; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15293 = 7'h1a == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_931 = 7'h1a == index | dirty_0_26; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15294 = 7'h1b == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_932 = 7'h1b == index | dirty_0_27; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15295 = 7'h1c == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_933 = 7'h1c == index | dirty_0_28; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15296 = 7'h1d == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_934 = 7'h1d == index | dirty_0_29; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15297 = 7'h1e == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_935 = 7'h1e == index | dirty_0_30; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15298 = 7'h1f == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_936 = 7'h1f == index | dirty_0_31; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15299 = 7'h20 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_937 = 7'h20 == index | dirty_0_32; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15300 = 7'h21 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_938 = 7'h21 == index | dirty_0_33; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15301 = 7'h22 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_939 = 7'h22 == index | dirty_0_34; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15302 = 7'h23 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_940 = 7'h23 == index | dirty_0_35; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15303 = 7'h24 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_941 = 7'h24 == index | dirty_0_36; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15304 = 7'h25 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_942 = 7'h25 == index | dirty_0_37; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15305 = 7'h26 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_943 = 7'h26 == index | dirty_0_38; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15306 = 7'h27 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_944 = 7'h27 == index | dirty_0_39; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15307 = 7'h28 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_945 = 7'h28 == index | dirty_0_40; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15308 = 7'h29 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_946 = 7'h29 == index | dirty_0_41; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15309 = 7'h2a == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_947 = 7'h2a == index | dirty_0_42; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15310 = 7'h2b == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_948 = 7'h2b == index | dirty_0_43; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15311 = 7'h2c == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_949 = 7'h2c == index | dirty_0_44; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15312 = 7'h2d == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_950 = 7'h2d == index | dirty_0_45; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15313 = 7'h2e == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_951 = 7'h2e == index | dirty_0_46; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15314 = 7'h2f == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_952 = 7'h2f == index | dirty_0_47; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15315 = 7'h30 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_953 = 7'h30 == index | dirty_0_48; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15316 = 7'h31 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_954 = 7'h31 == index | dirty_0_49; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15317 = 7'h32 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_955 = 7'h32 == index | dirty_0_50; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15318 = 7'h33 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_956 = 7'h33 == index | dirty_0_51; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15319 = 7'h34 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_957 = 7'h34 == index | dirty_0_52; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15320 = 7'h35 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_958 = 7'h35 == index | dirty_0_53; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15321 = 7'h36 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_959 = 7'h36 == index | dirty_0_54; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15322 = 7'h37 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_960 = 7'h37 == index | dirty_0_55; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15323 = 7'h38 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_961 = 7'h38 == index | dirty_0_56; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15324 = 7'h39 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_962 = 7'h39 == index | dirty_0_57; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15325 = 7'h3a == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_963 = 7'h3a == index | dirty_0_58; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15326 = 7'h3b == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_964 = 7'h3b == index | dirty_0_59; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15327 = 7'h3c == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_965 = 7'h3c == index | dirty_0_60; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15328 = 7'h3d == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_966 = 7'h3d == index | dirty_0_61; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15329 = 7'h3e == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_967 = 7'h3e == index | dirty_0_62; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15330 = 7'h3f == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_968 = 7'h3f == index | dirty_0_63; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15331 = 7'h40 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_969 = 7'h40 == index | dirty_0_64; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15332 = 7'h41 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_970 = 7'h41 == index | dirty_0_65; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15333 = 7'h42 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_971 = 7'h42 == index | dirty_0_66; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15334 = 7'h43 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_972 = 7'h43 == index | dirty_0_67; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15335 = 7'h44 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_973 = 7'h44 == index | dirty_0_68; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15336 = 7'h45 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_974 = 7'h45 == index | dirty_0_69; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15337 = 7'h46 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_975 = 7'h46 == index | dirty_0_70; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15338 = 7'h47 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_976 = 7'h47 == index | dirty_0_71; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15339 = 7'h48 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_977 = 7'h48 == index | dirty_0_72; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15340 = 7'h49 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_978 = 7'h49 == index | dirty_0_73; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15341 = 7'h4a == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_979 = 7'h4a == index | dirty_0_74; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15342 = 7'h4b == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_980 = 7'h4b == index | dirty_0_75; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15343 = 7'h4c == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_981 = 7'h4c == index | dirty_0_76; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15344 = 7'h4d == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_982 = 7'h4d == index | dirty_0_77; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15345 = 7'h4e == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_983 = 7'h4e == index | dirty_0_78; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15346 = 7'h4f == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_984 = 7'h4f == index | dirty_0_79; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15347 = 7'h50 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_985 = 7'h50 == index | dirty_0_80; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15348 = 7'h51 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_986 = 7'h51 == index | dirty_0_81; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15349 = 7'h52 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_987 = 7'h52 == index | dirty_0_82; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15350 = 7'h53 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_988 = 7'h53 == index | dirty_0_83; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15351 = 7'h54 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_989 = 7'h54 == index | dirty_0_84; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15352 = 7'h55 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_990 = 7'h55 == index | dirty_0_85; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15353 = 7'h56 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_991 = 7'h56 == index | dirty_0_86; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15354 = 7'h57 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_992 = 7'h57 == index | dirty_0_87; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15355 = 7'h58 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_993 = 7'h58 == index | dirty_0_88; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15356 = 7'h59 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_994 = 7'h59 == index | dirty_0_89; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15357 = 7'h5a == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_995 = 7'h5a == index | dirty_0_90; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15358 = 7'h5b == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_996 = 7'h5b == index | dirty_0_91; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15359 = 7'h5c == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_997 = 7'h5c == index | dirty_0_92; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15360 = 7'h5d == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_998 = 7'h5d == index | dirty_0_93; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15361 = 7'h5e == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_999 = 7'h5e == index | dirty_0_94; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15362 = 7'h5f == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1000 = 7'h5f == index | dirty_0_95; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15363 = 7'h60 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1001 = 7'h60 == index | dirty_0_96; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15364 = 7'h61 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1002 = 7'h61 == index | dirty_0_97; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15365 = 7'h62 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1003 = 7'h62 == index | dirty_0_98; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15366 = 7'h63 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1004 = 7'h63 == index | dirty_0_99; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15367 = 7'h64 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1005 = 7'h64 == index | dirty_0_100; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15368 = 7'h65 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1006 = 7'h65 == index | dirty_0_101; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15369 = 7'h66 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1007 = 7'h66 == index | dirty_0_102; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15370 = 7'h67 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1008 = 7'h67 == index | dirty_0_103; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15371 = 7'h68 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1009 = 7'h68 == index | dirty_0_104; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15372 = 7'h69 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1010 = 7'h69 == index | dirty_0_105; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15373 = 7'h6a == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1011 = 7'h6a == index | dirty_0_106; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15374 = 7'h6b == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1012 = 7'h6b == index | dirty_0_107; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15375 = 7'h6c == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1013 = 7'h6c == index | dirty_0_108; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15376 = 7'h6d == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1014 = 7'h6d == index | dirty_0_109; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15377 = 7'h6e == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1015 = 7'h6e == index | dirty_0_110; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15378 = 7'h6f == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1016 = 7'h6f == index | dirty_0_111; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15379 = 7'h70 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1017 = 7'h70 == index | dirty_0_112; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15380 = 7'h71 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1018 = 7'h71 == index | dirty_0_113; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15381 = 7'h72 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1019 = 7'h72 == index | dirty_0_114; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15382 = 7'h73 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1020 = 7'h73 == index | dirty_0_115; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15383 = 7'h74 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1021 = 7'h74 == index | dirty_0_116; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15384 = 7'h75 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1022 = 7'h75 == index | dirty_0_117; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15385 = 7'h76 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1023 = 7'h76 == index | dirty_0_118; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15386 = 7'h77 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1024 = 7'h77 == index | dirty_0_119; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15387 = 7'h78 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1025 = 7'h78 == index | dirty_0_120; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15388 = 7'h79 == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1026 = 7'h79 == index | dirty_0_121; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15389 = 7'h7a == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1027 = 7'h7a == index | dirty_0_122; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15390 = 7'h7b == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1028 = 7'h7b == index | dirty_0_123; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15391 = 7'h7c == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1029 = 7'h7c == index | dirty_0_124; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15392 = 7'h7d == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1030 = 7'h7d == index | dirty_0_125; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15393 = 7'h7e == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1031 = 7'h7e == index | dirty_0_126; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_15394 = 7'h7f == index; // @[d_cache.scala 24:26 94:{32,32}]
  wire  _GEN_1032 = 7'h7f == index | dirty_0_127; // @[d_cache.scala 24:26 94:{32,32}]
  wire [63:0] _GEN_1033 = 7'h0 == index ? _ram_0_index : ram_1_0; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1034 = 7'h1 == index ? _ram_0_index : ram_1_1; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1035 = 7'h2 == index ? _ram_0_index : ram_1_2; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1036 = 7'h3 == index ? _ram_0_index : ram_1_3; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1037 = 7'h4 == index ? _ram_0_index : ram_1_4; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1038 = 7'h5 == index ? _ram_0_index : ram_1_5; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1039 = 7'h6 == index ? _ram_0_index : ram_1_6; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1040 = 7'h7 == index ? _ram_0_index : ram_1_7; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1041 = 7'h8 == index ? _ram_0_index : ram_1_8; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1042 = 7'h9 == index ? _ram_0_index : ram_1_9; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1043 = 7'ha == index ? _ram_0_index : ram_1_10; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1044 = 7'hb == index ? _ram_0_index : ram_1_11; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1045 = 7'hc == index ? _ram_0_index : ram_1_12; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1046 = 7'hd == index ? _ram_0_index : ram_1_13; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1047 = 7'he == index ? _ram_0_index : ram_1_14; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1048 = 7'hf == index ? _ram_0_index : ram_1_15; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1049 = 7'h10 == index ? _ram_0_index : ram_1_16; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1050 = 7'h11 == index ? _ram_0_index : ram_1_17; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1051 = 7'h12 == index ? _ram_0_index : ram_1_18; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1052 = 7'h13 == index ? _ram_0_index : ram_1_19; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1053 = 7'h14 == index ? _ram_0_index : ram_1_20; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1054 = 7'h15 == index ? _ram_0_index : ram_1_21; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1055 = 7'h16 == index ? _ram_0_index : ram_1_22; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1056 = 7'h17 == index ? _ram_0_index : ram_1_23; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1057 = 7'h18 == index ? _ram_0_index : ram_1_24; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1058 = 7'h19 == index ? _ram_0_index : ram_1_25; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1059 = 7'h1a == index ? _ram_0_index : ram_1_26; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1060 = 7'h1b == index ? _ram_0_index : ram_1_27; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1061 = 7'h1c == index ? _ram_0_index : ram_1_28; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1062 = 7'h1d == index ? _ram_0_index : ram_1_29; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1063 = 7'h1e == index ? _ram_0_index : ram_1_30; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1064 = 7'h1f == index ? _ram_0_index : ram_1_31; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1065 = 7'h20 == index ? _ram_0_index : ram_1_32; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1066 = 7'h21 == index ? _ram_0_index : ram_1_33; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1067 = 7'h22 == index ? _ram_0_index : ram_1_34; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1068 = 7'h23 == index ? _ram_0_index : ram_1_35; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1069 = 7'h24 == index ? _ram_0_index : ram_1_36; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1070 = 7'h25 == index ? _ram_0_index : ram_1_37; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1071 = 7'h26 == index ? _ram_0_index : ram_1_38; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1072 = 7'h27 == index ? _ram_0_index : ram_1_39; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1073 = 7'h28 == index ? _ram_0_index : ram_1_40; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1074 = 7'h29 == index ? _ram_0_index : ram_1_41; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1075 = 7'h2a == index ? _ram_0_index : ram_1_42; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1076 = 7'h2b == index ? _ram_0_index : ram_1_43; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1077 = 7'h2c == index ? _ram_0_index : ram_1_44; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1078 = 7'h2d == index ? _ram_0_index : ram_1_45; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1079 = 7'h2e == index ? _ram_0_index : ram_1_46; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1080 = 7'h2f == index ? _ram_0_index : ram_1_47; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1081 = 7'h30 == index ? _ram_0_index : ram_1_48; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1082 = 7'h31 == index ? _ram_0_index : ram_1_49; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1083 = 7'h32 == index ? _ram_0_index : ram_1_50; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1084 = 7'h33 == index ? _ram_0_index : ram_1_51; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1085 = 7'h34 == index ? _ram_0_index : ram_1_52; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1086 = 7'h35 == index ? _ram_0_index : ram_1_53; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1087 = 7'h36 == index ? _ram_0_index : ram_1_54; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1088 = 7'h37 == index ? _ram_0_index : ram_1_55; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1089 = 7'h38 == index ? _ram_0_index : ram_1_56; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1090 = 7'h39 == index ? _ram_0_index : ram_1_57; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1091 = 7'h3a == index ? _ram_0_index : ram_1_58; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1092 = 7'h3b == index ? _ram_0_index : ram_1_59; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1093 = 7'h3c == index ? _ram_0_index : ram_1_60; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1094 = 7'h3d == index ? _ram_0_index : ram_1_61; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1095 = 7'h3e == index ? _ram_0_index : ram_1_62; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1096 = 7'h3f == index ? _ram_0_index : ram_1_63; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1097 = 7'h40 == index ? _ram_0_index : ram_1_64; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1098 = 7'h41 == index ? _ram_0_index : ram_1_65; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1099 = 7'h42 == index ? _ram_0_index : ram_1_66; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1100 = 7'h43 == index ? _ram_0_index : ram_1_67; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1101 = 7'h44 == index ? _ram_0_index : ram_1_68; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1102 = 7'h45 == index ? _ram_0_index : ram_1_69; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1103 = 7'h46 == index ? _ram_0_index : ram_1_70; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1104 = 7'h47 == index ? _ram_0_index : ram_1_71; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1105 = 7'h48 == index ? _ram_0_index : ram_1_72; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1106 = 7'h49 == index ? _ram_0_index : ram_1_73; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1107 = 7'h4a == index ? _ram_0_index : ram_1_74; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1108 = 7'h4b == index ? _ram_0_index : ram_1_75; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1109 = 7'h4c == index ? _ram_0_index : ram_1_76; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1110 = 7'h4d == index ? _ram_0_index : ram_1_77; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1111 = 7'h4e == index ? _ram_0_index : ram_1_78; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1112 = 7'h4f == index ? _ram_0_index : ram_1_79; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1113 = 7'h50 == index ? _ram_0_index : ram_1_80; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1114 = 7'h51 == index ? _ram_0_index : ram_1_81; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1115 = 7'h52 == index ? _ram_0_index : ram_1_82; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1116 = 7'h53 == index ? _ram_0_index : ram_1_83; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1117 = 7'h54 == index ? _ram_0_index : ram_1_84; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1118 = 7'h55 == index ? _ram_0_index : ram_1_85; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1119 = 7'h56 == index ? _ram_0_index : ram_1_86; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1120 = 7'h57 == index ? _ram_0_index : ram_1_87; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1121 = 7'h58 == index ? _ram_0_index : ram_1_88; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1122 = 7'h59 == index ? _ram_0_index : ram_1_89; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1123 = 7'h5a == index ? _ram_0_index : ram_1_90; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1124 = 7'h5b == index ? _ram_0_index : ram_1_91; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1125 = 7'h5c == index ? _ram_0_index : ram_1_92; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1126 = 7'h5d == index ? _ram_0_index : ram_1_93; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1127 = 7'h5e == index ? _ram_0_index : ram_1_94; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1128 = 7'h5f == index ? _ram_0_index : ram_1_95; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1129 = 7'h60 == index ? _ram_0_index : ram_1_96; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1130 = 7'h61 == index ? _ram_0_index : ram_1_97; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1131 = 7'h62 == index ? _ram_0_index : ram_1_98; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1132 = 7'h63 == index ? _ram_0_index : ram_1_99; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1133 = 7'h64 == index ? _ram_0_index : ram_1_100; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1134 = 7'h65 == index ? _ram_0_index : ram_1_101; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1135 = 7'h66 == index ? _ram_0_index : ram_1_102; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1136 = 7'h67 == index ? _ram_0_index : ram_1_103; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1137 = 7'h68 == index ? _ram_0_index : ram_1_104; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1138 = 7'h69 == index ? _ram_0_index : ram_1_105; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1139 = 7'h6a == index ? _ram_0_index : ram_1_106; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1140 = 7'h6b == index ? _ram_0_index : ram_1_107; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1141 = 7'h6c == index ? _ram_0_index : ram_1_108; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1142 = 7'h6d == index ? _ram_0_index : ram_1_109; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1143 = 7'h6e == index ? _ram_0_index : ram_1_110; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1144 = 7'h6f == index ? _ram_0_index : ram_1_111; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1145 = 7'h70 == index ? _ram_0_index : ram_1_112; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1146 = 7'h71 == index ? _ram_0_index : ram_1_113; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1147 = 7'h72 == index ? _ram_0_index : ram_1_114; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1148 = 7'h73 == index ? _ram_0_index : ram_1_115; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1149 = 7'h74 == index ? _ram_0_index : ram_1_116; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1150 = 7'h75 == index ? _ram_0_index : ram_1_117; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1151 = 7'h76 == index ? _ram_0_index : ram_1_118; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1152 = 7'h77 == index ? _ram_0_index : ram_1_119; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1153 = 7'h78 == index ? _ram_0_index : ram_1_120; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1154 = 7'h79 == index ? _ram_0_index : ram_1_121; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1155 = 7'h7a == index ? _ram_0_index : ram_1_122; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1156 = 7'h7b == index ? _ram_0_index : ram_1_123; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1157 = 7'h7c == index ? _ram_0_index : ram_1_124; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1158 = 7'h7d == index ? _ram_0_index : ram_1_125; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1159 = 7'h7e == index ? _ram_0_index : ram_1_126; // @[d_cache.scala 19:24 98:{30,30}]
  wire [63:0] _GEN_1160 = 7'h7f == index ? _ram_0_index : ram_1_127; // @[d_cache.scala 19:24 98:{30,30}]
  wire  _GEN_1161 = _GEN_15267 | dirty_1_0; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1162 = _GEN_15268 | dirty_1_1; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1163 = _GEN_15269 | dirty_1_2; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1164 = _GEN_15270 | dirty_1_3; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1165 = _GEN_15271 | dirty_1_4; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1166 = _GEN_15272 | dirty_1_5; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1167 = _GEN_15273 | dirty_1_6; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1168 = _GEN_15274 | dirty_1_7; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1169 = _GEN_15275 | dirty_1_8; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1170 = _GEN_15276 | dirty_1_9; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1171 = _GEN_15277 | dirty_1_10; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1172 = _GEN_15278 | dirty_1_11; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1173 = _GEN_15279 | dirty_1_12; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1174 = _GEN_15280 | dirty_1_13; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1175 = _GEN_15281 | dirty_1_14; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1176 = _GEN_15282 | dirty_1_15; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1177 = _GEN_15283 | dirty_1_16; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1178 = _GEN_15284 | dirty_1_17; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1179 = _GEN_15285 | dirty_1_18; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1180 = _GEN_15286 | dirty_1_19; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1181 = _GEN_15287 | dirty_1_20; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1182 = _GEN_15288 | dirty_1_21; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1183 = _GEN_15289 | dirty_1_22; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1184 = _GEN_15290 | dirty_1_23; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1185 = _GEN_15291 | dirty_1_24; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1186 = _GEN_15292 | dirty_1_25; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1187 = _GEN_15293 | dirty_1_26; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1188 = _GEN_15294 | dirty_1_27; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1189 = _GEN_15295 | dirty_1_28; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1190 = _GEN_15296 | dirty_1_29; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1191 = _GEN_15297 | dirty_1_30; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1192 = _GEN_15298 | dirty_1_31; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1193 = _GEN_15299 | dirty_1_32; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1194 = _GEN_15300 | dirty_1_33; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1195 = _GEN_15301 | dirty_1_34; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1196 = _GEN_15302 | dirty_1_35; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1197 = _GEN_15303 | dirty_1_36; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1198 = _GEN_15304 | dirty_1_37; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1199 = _GEN_15305 | dirty_1_38; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1200 = _GEN_15306 | dirty_1_39; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1201 = _GEN_15307 | dirty_1_40; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1202 = _GEN_15308 | dirty_1_41; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1203 = _GEN_15309 | dirty_1_42; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1204 = _GEN_15310 | dirty_1_43; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1205 = _GEN_15311 | dirty_1_44; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1206 = _GEN_15312 | dirty_1_45; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1207 = _GEN_15313 | dirty_1_46; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1208 = _GEN_15314 | dirty_1_47; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1209 = _GEN_15315 | dirty_1_48; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1210 = _GEN_15316 | dirty_1_49; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1211 = _GEN_15317 | dirty_1_50; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1212 = _GEN_15318 | dirty_1_51; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1213 = _GEN_15319 | dirty_1_52; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1214 = _GEN_15320 | dirty_1_53; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1215 = _GEN_15321 | dirty_1_54; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1216 = _GEN_15322 | dirty_1_55; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1217 = _GEN_15323 | dirty_1_56; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1218 = _GEN_15324 | dirty_1_57; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1219 = _GEN_15325 | dirty_1_58; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1220 = _GEN_15326 | dirty_1_59; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1221 = _GEN_15327 | dirty_1_60; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1222 = _GEN_15328 | dirty_1_61; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1223 = _GEN_15329 | dirty_1_62; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1224 = _GEN_15330 | dirty_1_63; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1225 = _GEN_15331 | dirty_1_64; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1226 = _GEN_15332 | dirty_1_65; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1227 = _GEN_15333 | dirty_1_66; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1228 = _GEN_15334 | dirty_1_67; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1229 = _GEN_15335 | dirty_1_68; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1230 = _GEN_15336 | dirty_1_69; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1231 = _GEN_15337 | dirty_1_70; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1232 = _GEN_15338 | dirty_1_71; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1233 = _GEN_15339 | dirty_1_72; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1234 = _GEN_15340 | dirty_1_73; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1235 = _GEN_15341 | dirty_1_74; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1236 = _GEN_15342 | dirty_1_75; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1237 = _GEN_15343 | dirty_1_76; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1238 = _GEN_15344 | dirty_1_77; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1239 = _GEN_15345 | dirty_1_78; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1240 = _GEN_15346 | dirty_1_79; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1241 = _GEN_15347 | dirty_1_80; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1242 = _GEN_15348 | dirty_1_81; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1243 = _GEN_15349 | dirty_1_82; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1244 = _GEN_15350 | dirty_1_83; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1245 = _GEN_15351 | dirty_1_84; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1246 = _GEN_15352 | dirty_1_85; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1247 = _GEN_15353 | dirty_1_86; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1248 = _GEN_15354 | dirty_1_87; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1249 = _GEN_15355 | dirty_1_88; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1250 = _GEN_15356 | dirty_1_89; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1251 = _GEN_15357 | dirty_1_90; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1252 = _GEN_15358 | dirty_1_91; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1253 = _GEN_15359 | dirty_1_92; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1254 = _GEN_15360 | dirty_1_93; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1255 = _GEN_15361 | dirty_1_94; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1256 = _GEN_15362 | dirty_1_95; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1257 = _GEN_15363 | dirty_1_96; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1258 = _GEN_15364 | dirty_1_97; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1259 = _GEN_15365 | dirty_1_98; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1260 = _GEN_15366 | dirty_1_99; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1261 = _GEN_15367 | dirty_1_100; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1262 = _GEN_15368 | dirty_1_101; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1263 = _GEN_15369 | dirty_1_102; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1264 = _GEN_15370 | dirty_1_103; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1265 = _GEN_15371 | dirty_1_104; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1266 = _GEN_15372 | dirty_1_105; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1267 = _GEN_15373 | dirty_1_106; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1268 = _GEN_15374 | dirty_1_107; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1269 = _GEN_15375 | dirty_1_108; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1270 = _GEN_15376 | dirty_1_109; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1271 = _GEN_15377 | dirty_1_110; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1272 = _GEN_15378 | dirty_1_111; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1273 = _GEN_15379 | dirty_1_112; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1274 = _GEN_15380 | dirty_1_113; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1275 = _GEN_15381 | dirty_1_114; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1276 = _GEN_15382 | dirty_1_115; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1277 = _GEN_15383 | dirty_1_116; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1278 = _GEN_15384 | dirty_1_117; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1279 = _GEN_15385 | dirty_1_118; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1280 = _GEN_15386 | dirty_1_119; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1281 = _GEN_15387 | dirty_1_120; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1282 = _GEN_15388 | dirty_1_121; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1283 = _GEN_15389 | dirty_1_122; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1284 = _GEN_15390 | dirty_1_123; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1285 = _GEN_15391 | dirty_1_124; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1286 = _GEN_15392 | dirty_1_125; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1287 = _GEN_15393 | dirty_1_126; // @[d_cache.scala 100:{32,32} 25:26]
  wire  _GEN_1288 = _GEN_15394 | dirty_1_127; // @[d_cache.scala 100:{32,32} 25:26]
  wire [2:0] _GEN_1289 = way1_hit ? 3'h0 : 3'h4; // @[d_cache.scala 102:23 96:33 97:23]
  wire [63:0] _GEN_1290 = way1_hit ? _GEN_1033 : ram_1_0; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1291 = way1_hit ? _GEN_1034 : ram_1_1; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1292 = way1_hit ? _GEN_1035 : ram_1_2; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1293 = way1_hit ? _GEN_1036 : ram_1_3; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1294 = way1_hit ? _GEN_1037 : ram_1_4; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1295 = way1_hit ? _GEN_1038 : ram_1_5; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1296 = way1_hit ? _GEN_1039 : ram_1_6; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1297 = way1_hit ? _GEN_1040 : ram_1_7; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1298 = way1_hit ? _GEN_1041 : ram_1_8; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1299 = way1_hit ? _GEN_1042 : ram_1_9; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1300 = way1_hit ? _GEN_1043 : ram_1_10; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1301 = way1_hit ? _GEN_1044 : ram_1_11; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1302 = way1_hit ? _GEN_1045 : ram_1_12; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1303 = way1_hit ? _GEN_1046 : ram_1_13; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1304 = way1_hit ? _GEN_1047 : ram_1_14; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1305 = way1_hit ? _GEN_1048 : ram_1_15; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1306 = way1_hit ? _GEN_1049 : ram_1_16; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1307 = way1_hit ? _GEN_1050 : ram_1_17; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1308 = way1_hit ? _GEN_1051 : ram_1_18; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1309 = way1_hit ? _GEN_1052 : ram_1_19; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1310 = way1_hit ? _GEN_1053 : ram_1_20; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1311 = way1_hit ? _GEN_1054 : ram_1_21; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1312 = way1_hit ? _GEN_1055 : ram_1_22; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1313 = way1_hit ? _GEN_1056 : ram_1_23; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1314 = way1_hit ? _GEN_1057 : ram_1_24; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1315 = way1_hit ? _GEN_1058 : ram_1_25; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1316 = way1_hit ? _GEN_1059 : ram_1_26; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1317 = way1_hit ? _GEN_1060 : ram_1_27; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1318 = way1_hit ? _GEN_1061 : ram_1_28; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1319 = way1_hit ? _GEN_1062 : ram_1_29; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1320 = way1_hit ? _GEN_1063 : ram_1_30; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1321 = way1_hit ? _GEN_1064 : ram_1_31; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1322 = way1_hit ? _GEN_1065 : ram_1_32; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1323 = way1_hit ? _GEN_1066 : ram_1_33; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1324 = way1_hit ? _GEN_1067 : ram_1_34; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1325 = way1_hit ? _GEN_1068 : ram_1_35; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1326 = way1_hit ? _GEN_1069 : ram_1_36; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1327 = way1_hit ? _GEN_1070 : ram_1_37; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1328 = way1_hit ? _GEN_1071 : ram_1_38; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1329 = way1_hit ? _GEN_1072 : ram_1_39; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1330 = way1_hit ? _GEN_1073 : ram_1_40; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1331 = way1_hit ? _GEN_1074 : ram_1_41; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1332 = way1_hit ? _GEN_1075 : ram_1_42; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1333 = way1_hit ? _GEN_1076 : ram_1_43; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1334 = way1_hit ? _GEN_1077 : ram_1_44; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1335 = way1_hit ? _GEN_1078 : ram_1_45; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1336 = way1_hit ? _GEN_1079 : ram_1_46; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1337 = way1_hit ? _GEN_1080 : ram_1_47; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1338 = way1_hit ? _GEN_1081 : ram_1_48; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1339 = way1_hit ? _GEN_1082 : ram_1_49; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1340 = way1_hit ? _GEN_1083 : ram_1_50; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1341 = way1_hit ? _GEN_1084 : ram_1_51; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1342 = way1_hit ? _GEN_1085 : ram_1_52; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1343 = way1_hit ? _GEN_1086 : ram_1_53; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1344 = way1_hit ? _GEN_1087 : ram_1_54; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1345 = way1_hit ? _GEN_1088 : ram_1_55; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1346 = way1_hit ? _GEN_1089 : ram_1_56; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1347 = way1_hit ? _GEN_1090 : ram_1_57; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1348 = way1_hit ? _GEN_1091 : ram_1_58; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1349 = way1_hit ? _GEN_1092 : ram_1_59; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1350 = way1_hit ? _GEN_1093 : ram_1_60; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1351 = way1_hit ? _GEN_1094 : ram_1_61; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1352 = way1_hit ? _GEN_1095 : ram_1_62; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1353 = way1_hit ? _GEN_1096 : ram_1_63; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1354 = way1_hit ? _GEN_1097 : ram_1_64; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1355 = way1_hit ? _GEN_1098 : ram_1_65; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1356 = way1_hit ? _GEN_1099 : ram_1_66; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1357 = way1_hit ? _GEN_1100 : ram_1_67; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1358 = way1_hit ? _GEN_1101 : ram_1_68; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1359 = way1_hit ? _GEN_1102 : ram_1_69; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1360 = way1_hit ? _GEN_1103 : ram_1_70; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1361 = way1_hit ? _GEN_1104 : ram_1_71; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1362 = way1_hit ? _GEN_1105 : ram_1_72; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1363 = way1_hit ? _GEN_1106 : ram_1_73; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1364 = way1_hit ? _GEN_1107 : ram_1_74; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1365 = way1_hit ? _GEN_1108 : ram_1_75; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1366 = way1_hit ? _GEN_1109 : ram_1_76; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1367 = way1_hit ? _GEN_1110 : ram_1_77; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1368 = way1_hit ? _GEN_1111 : ram_1_78; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1369 = way1_hit ? _GEN_1112 : ram_1_79; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1370 = way1_hit ? _GEN_1113 : ram_1_80; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1371 = way1_hit ? _GEN_1114 : ram_1_81; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1372 = way1_hit ? _GEN_1115 : ram_1_82; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1373 = way1_hit ? _GEN_1116 : ram_1_83; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1374 = way1_hit ? _GEN_1117 : ram_1_84; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1375 = way1_hit ? _GEN_1118 : ram_1_85; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1376 = way1_hit ? _GEN_1119 : ram_1_86; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1377 = way1_hit ? _GEN_1120 : ram_1_87; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1378 = way1_hit ? _GEN_1121 : ram_1_88; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1379 = way1_hit ? _GEN_1122 : ram_1_89; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1380 = way1_hit ? _GEN_1123 : ram_1_90; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1381 = way1_hit ? _GEN_1124 : ram_1_91; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1382 = way1_hit ? _GEN_1125 : ram_1_92; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1383 = way1_hit ? _GEN_1126 : ram_1_93; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1384 = way1_hit ? _GEN_1127 : ram_1_94; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1385 = way1_hit ? _GEN_1128 : ram_1_95; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1386 = way1_hit ? _GEN_1129 : ram_1_96; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1387 = way1_hit ? _GEN_1130 : ram_1_97; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1388 = way1_hit ? _GEN_1131 : ram_1_98; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1389 = way1_hit ? _GEN_1132 : ram_1_99; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1390 = way1_hit ? _GEN_1133 : ram_1_100; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1391 = way1_hit ? _GEN_1134 : ram_1_101; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1392 = way1_hit ? _GEN_1135 : ram_1_102; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1393 = way1_hit ? _GEN_1136 : ram_1_103; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1394 = way1_hit ? _GEN_1137 : ram_1_104; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1395 = way1_hit ? _GEN_1138 : ram_1_105; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1396 = way1_hit ? _GEN_1139 : ram_1_106; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1397 = way1_hit ? _GEN_1140 : ram_1_107; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1398 = way1_hit ? _GEN_1141 : ram_1_108; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1399 = way1_hit ? _GEN_1142 : ram_1_109; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1400 = way1_hit ? _GEN_1143 : ram_1_110; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1401 = way1_hit ? _GEN_1144 : ram_1_111; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1402 = way1_hit ? _GEN_1145 : ram_1_112; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1403 = way1_hit ? _GEN_1146 : ram_1_113; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1404 = way1_hit ? _GEN_1147 : ram_1_114; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1405 = way1_hit ? _GEN_1148 : ram_1_115; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1406 = way1_hit ? _GEN_1149 : ram_1_116; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1407 = way1_hit ? _GEN_1150 : ram_1_117; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1408 = way1_hit ? _GEN_1151 : ram_1_118; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1409 = way1_hit ? _GEN_1152 : ram_1_119; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1410 = way1_hit ? _GEN_1153 : ram_1_120; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1411 = way1_hit ? _GEN_1154 : ram_1_121; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1412 = way1_hit ? _GEN_1155 : ram_1_122; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1413 = way1_hit ? _GEN_1156 : ram_1_123; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1414 = way1_hit ? _GEN_1157 : ram_1_124; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1415 = way1_hit ? _GEN_1158 : ram_1_125; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1416 = way1_hit ? _GEN_1159 : ram_1_126; // @[d_cache.scala 19:24 96:33]
  wire [63:0] _GEN_1417 = way1_hit ? _GEN_1160 : ram_1_127; // @[d_cache.scala 19:24 96:33]
  wire  _GEN_1418 = way1_hit ? _GEN_1161 : dirty_1_0; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1419 = way1_hit ? _GEN_1162 : dirty_1_1; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1420 = way1_hit ? _GEN_1163 : dirty_1_2; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1421 = way1_hit ? _GEN_1164 : dirty_1_3; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1422 = way1_hit ? _GEN_1165 : dirty_1_4; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1423 = way1_hit ? _GEN_1166 : dirty_1_5; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1424 = way1_hit ? _GEN_1167 : dirty_1_6; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1425 = way1_hit ? _GEN_1168 : dirty_1_7; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1426 = way1_hit ? _GEN_1169 : dirty_1_8; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1427 = way1_hit ? _GEN_1170 : dirty_1_9; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1428 = way1_hit ? _GEN_1171 : dirty_1_10; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1429 = way1_hit ? _GEN_1172 : dirty_1_11; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1430 = way1_hit ? _GEN_1173 : dirty_1_12; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1431 = way1_hit ? _GEN_1174 : dirty_1_13; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1432 = way1_hit ? _GEN_1175 : dirty_1_14; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1433 = way1_hit ? _GEN_1176 : dirty_1_15; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1434 = way1_hit ? _GEN_1177 : dirty_1_16; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1435 = way1_hit ? _GEN_1178 : dirty_1_17; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1436 = way1_hit ? _GEN_1179 : dirty_1_18; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1437 = way1_hit ? _GEN_1180 : dirty_1_19; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1438 = way1_hit ? _GEN_1181 : dirty_1_20; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1439 = way1_hit ? _GEN_1182 : dirty_1_21; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1440 = way1_hit ? _GEN_1183 : dirty_1_22; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1441 = way1_hit ? _GEN_1184 : dirty_1_23; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1442 = way1_hit ? _GEN_1185 : dirty_1_24; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1443 = way1_hit ? _GEN_1186 : dirty_1_25; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1444 = way1_hit ? _GEN_1187 : dirty_1_26; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1445 = way1_hit ? _GEN_1188 : dirty_1_27; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1446 = way1_hit ? _GEN_1189 : dirty_1_28; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1447 = way1_hit ? _GEN_1190 : dirty_1_29; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1448 = way1_hit ? _GEN_1191 : dirty_1_30; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1449 = way1_hit ? _GEN_1192 : dirty_1_31; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1450 = way1_hit ? _GEN_1193 : dirty_1_32; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1451 = way1_hit ? _GEN_1194 : dirty_1_33; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1452 = way1_hit ? _GEN_1195 : dirty_1_34; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1453 = way1_hit ? _GEN_1196 : dirty_1_35; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1454 = way1_hit ? _GEN_1197 : dirty_1_36; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1455 = way1_hit ? _GEN_1198 : dirty_1_37; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1456 = way1_hit ? _GEN_1199 : dirty_1_38; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1457 = way1_hit ? _GEN_1200 : dirty_1_39; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1458 = way1_hit ? _GEN_1201 : dirty_1_40; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1459 = way1_hit ? _GEN_1202 : dirty_1_41; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1460 = way1_hit ? _GEN_1203 : dirty_1_42; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1461 = way1_hit ? _GEN_1204 : dirty_1_43; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1462 = way1_hit ? _GEN_1205 : dirty_1_44; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1463 = way1_hit ? _GEN_1206 : dirty_1_45; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1464 = way1_hit ? _GEN_1207 : dirty_1_46; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1465 = way1_hit ? _GEN_1208 : dirty_1_47; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1466 = way1_hit ? _GEN_1209 : dirty_1_48; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1467 = way1_hit ? _GEN_1210 : dirty_1_49; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1468 = way1_hit ? _GEN_1211 : dirty_1_50; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1469 = way1_hit ? _GEN_1212 : dirty_1_51; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1470 = way1_hit ? _GEN_1213 : dirty_1_52; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1471 = way1_hit ? _GEN_1214 : dirty_1_53; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1472 = way1_hit ? _GEN_1215 : dirty_1_54; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1473 = way1_hit ? _GEN_1216 : dirty_1_55; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1474 = way1_hit ? _GEN_1217 : dirty_1_56; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1475 = way1_hit ? _GEN_1218 : dirty_1_57; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1476 = way1_hit ? _GEN_1219 : dirty_1_58; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1477 = way1_hit ? _GEN_1220 : dirty_1_59; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1478 = way1_hit ? _GEN_1221 : dirty_1_60; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1479 = way1_hit ? _GEN_1222 : dirty_1_61; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1480 = way1_hit ? _GEN_1223 : dirty_1_62; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1481 = way1_hit ? _GEN_1224 : dirty_1_63; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1482 = way1_hit ? _GEN_1225 : dirty_1_64; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1483 = way1_hit ? _GEN_1226 : dirty_1_65; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1484 = way1_hit ? _GEN_1227 : dirty_1_66; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1485 = way1_hit ? _GEN_1228 : dirty_1_67; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1486 = way1_hit ? _GEN_1229 : dirty_1_68; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1487 = way1_hit ? _GEN_1230 : dirty_1_69; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1488 = way1_hit ? _GEN_1231 : dirty_1_70; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1489 = way1_hit ? _GEN_1232 : dirty_1_71; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1490 = way1_hit ? _GEN_1233 : dirty_1_72; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1491 = way1_hit ? _GEN_1234 : dirty_1_73; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1492 = way1_hit ? _GEN_1235 : dirty_1_74; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1493 = way1_hit ? _GEN_1236 : dirty_1_75; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1494 = way1_hit ? _GEN_1237 : dirty_1_76; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1495 = way1_hit ? _GEN_1238 : dirty_1_77; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1496 = way1_hit ? _GEN_1239 : dirty_1_78; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1497 = way1_hit ? _GEN_1240 : dirty_1_79; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1498 = way1_hit ? _GEN_1241 : dirty_1_80; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1499 = way1_hit ? _GEN_1242 : dirty_1_81; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1500 = way1_hit ? _GEN_1243 : dirty_1_82; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1501 = way1_hit ? _GEN_1244 : dirty_1_83; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1502 = way1_hit ? _GEN_1245 : dirty_1_84; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1503 = way1_hit ? _GEN_1246 : dirty_1_85; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1504 = way1_hit ? _GEN_1247 : dirty_1_86; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1505 = way1_hit ? _GEN_1248 : dirty_1_87; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1506 = way1_hit ? _GEN_1249 : dirty_1_88; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1507 = way1_hit ? _GEN_1250 : dirty_1_89; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1508 = way1_hit ? _GEN_1251 : dirty_1_90; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1509 = way1_hit ? _GEN_1252 : dirty_1_91; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1510 = way1_hit ? _GEN_1253 : dirty_1_92; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1511 = way1_hit ? _GEN_1254 : dirty_1_93; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1512 = way1_hit ? _GEN_1255 : dirty_1_94; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1513 = way1_hit ? _GEN_1256 : dirty_1_95; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1514 = way1_hit ? _GEN_1257 : dirty_1_96; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1515 = way1_hit ? _GEN_1258 : dirty_1_97; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1516 = way1_hit ? _GEN_1259 : dirty_1_98; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1517 = way1_hit ? _GEN_1260 : dirty_1_99; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1518 = way1_hit ? _GEN_1261 : dirty_1_100; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1519 = way1_hit ? _GEN_1262 : dirty_1_101; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1520 = way1_hit ? _GEN_1263 : dirty_1_102; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1521 = way1_hit ? _GEN_1264 : dirty_1_103; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1522 = way1_hit ? _GEN_1265 : dirty_1_104; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1523 = way1_hit ? _GEN_1266 : dirty_1_105; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1524 = way1_hit ? _GEN_1267 : dirty_1_106; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1525 = way1_hit ? _GEN_1268 : dirty_1_107; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1526 = way1_hit ? _GEN_1269 : dirty_1_108; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1527 = way1_hit ? _GEN_1270 : dirty_1_109; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1528 = way1_hit ? _GEN_1271 : dirty_1_110; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1529 = way1_hit ? _GEN_1272 : dirty_1_111; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1530 = way1_hit ? _GEN_1273 : dirty_1_112; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1531 = way1_hit ? _GEN_1274 : dirty_1_113; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1532 = way1_hit ? _GEN_1275 : dirty_1_114; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1533 = way1_hit ? _GEN_1276 : dirty_1_115; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1534 = way1_hit ? _GEN_1277 : dirty_1_116; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1535 = way1_hit ? _GEN_1278 : dirty_1_117; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1536 = way1_hit ? _GEN_1279 : dirty_1_118; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1537 = way1_hit ? _GEN_1280 : dirty_1_119; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1538 = way1_hit ? _GEN_1281 : dirty_1_120; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1539 = way1_hit ? _GEN_1282 : dirty_1_121; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1540 = way1_hit ? _GEN_1283 : dirty_1_122; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1541 = way1_hit ? _GEN_1284 : dirty_1_123; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1542 = way1_hit ? _GEN_1285 : dirty_1_124; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1543 = way1_hit ? _GEN_1286 : dirty_1_125; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1544 = way1_hit ? _GEN_1287 : dirty_1_126; // @[d_cache.scala 25:26 96:33]
  wire  _GEN_1545 = way1_hit ? _GEN_1288 : dirty_1_127; // @[d_cache.scala 25:26 96:33]
  wire [2:0] _GEN_1546 = way0_hit ? 3'h0 : _GEN_1289; // @[d_cache.scala 90:27 91:23]
  wire [63:0] _GEN_1547 = way0_hit ? _GEN_777 : ram_0_0; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1548 = way0_hit ? _GEN_778 : ram_0_1; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1549 = way0_hit ? _GEN_779 : ram_0_2; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1550 = way0_hit ? _GEN_780 : ram_0_3; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1551 = way0_hit ? _GEN_781 : ram_0_4; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1552 = way0_hit ? _GEN_782 : ram_0_5; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1553 = way0_hit ? _GEN_783 : ram_0_6; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1554 = way0_hit ? _GEN_784 : ram_0_7; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1555 = way0_hit ? _GEN_785 : ram_0_8; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1556 = way0_hit ? _GEN_786 : ram_0_9; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1557 = way0_hit ? _GEN_787 : ram_0_10; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1558 = way0_hit ? _GEN_788 : ram_0_11; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1559 = way0_hit ? _GEN_789 : ram_0_12; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1560 = way0_hit ? _GEN_790 : ram_0_13; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1561 = way0_hit ? _GEN_791 : ram_0_14; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1562 = way0_hit ? _GEN_792 : ram_0_15; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1563 = way0_hit ? _GEN_793 : ram_0_16; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1564 = way0_hit ? _GEN_794 : ram_0_17; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1565 = way0_hit ? _GEN_795 : ram_0_18; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1566 = way0_hit ? _GEN_796 : ram_0_19; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1567 = way0_hit ? _GEN_797 : ram_0_20; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1568 = way0_hit ? _GEN_798 : ram_0_21; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1569 = way0_hit ? _GEN_799 : ram_0_22; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1570 = way0_hit ? _GEN_800 : ram_0_23; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1571 = way0_hit ? _GEN_801 : ram_0_24; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1572 = way0_hit ? _GEN_802 : ram_0_25; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1573 = way0_hit ? _GEN_803 : ram_0_26; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1574 = way0_hit ? _GEN_804 : ram_0_27; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1575 = way0_hit ? _GEN_805 : ram_0_28; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1576 = way0_hit ? _GEN_806 : ram_0_29; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1577 = way0_hit ? _GEN_807 : ram_0_30; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1578 = way0_hit ? _GEN_808 : ram_0_31; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1579 = way0_hit ? _GEN_809 : ram_0_32; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1580 = way0_hit ? _GEN_810 : ram_0_33; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1581 = way0_hit ? _GEN_811 : ram_0_34; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1582 = way0_hit ? _GEN_812 : ram_0_35; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1583 = way0_hit ? _GEN_813 : ram_0_36; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1584 = way0_hit ? _GEN_814 : ram_0_37; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1585 = way0_hit ? _GEN_815 : ram_0_38; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1586 = way0_hit ? _GEN_816 : ram_0_39; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1587 = way0_hit ? _GEN_817 : ram_0_40; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1588 = way0_hit ? _GEN_818 : ram_0_41; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1589 = way0_hit ? _GEN_819 : ram_0_42; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1590 = way0_hit ? _GEN_820 : ram_0_43; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1591 = way0_hit ? _GEN_821 : ram_0_44; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1592 = way0_hit ? _GEN_822 : ram_0_45; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1593 = way0_hit ? _GEN_823 : ram_0_46; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1594 = way0_hit ? _GEN_824 : ram_0_47; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1595 = way0_hit ? _GEN_825 : ram_0_48; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1596 = way0_hit ? _GEN_826 : ram_0_49; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1597 = way0_hit ? _GEN_827 : ram_0_50; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1598 = way0_hit ? _GEN_828 : ram_0_51; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1599 = way0_hit ? _GEN_829 : ram_0_52; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1600 = way0_hit ? _GEN_830 : ram_0_53; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1601 = way0_hit ? _GEN_831 : ram_0_54; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1602 = way0_hit ? _GEN_832 : ram_0_55; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1603 = way0_hit ? _GEN_833 : ram_0_56; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1604 = way0_hit ? _GEN_834 : ram_0_57; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1605 = way0_hit ? _GEN_835 : ram_0_58; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1606 = way0_hit ? _GEN_836 : ram_0_59; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1607 = way0_hit ? _GEN_837 : ram_0_60; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1608 = way0_hit ? _GEN_838 : ram_0_61; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1609 = way0_hit ? _GEN_839 : ram_0_62; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1610 = way0_hit ? _GEN_840 : ram_0_63; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1611 = way0_hit ? _GEN_841 : ram_0_64; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1612 = way0_hit ? _GEN_842 : ram_0_65; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1613 = way0_hit ? _GEN_843 : ram_0_66; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1614 = way0_hit ? _GEN_844 : ram_0_67; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1615 = way0_hit ? _GEN_845 : ram_0_68; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1616 = way0_hit ? _GEN_846 : ram_0_69; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1617 = way0_hit ? _GEN_847 : ram_0_70; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1618 = way0_hit ? _GEN_848 : ram_0_71; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1619 = way0_hit ? _GEN_849 : ram_0_72; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1620 = way0_hit ? _GEN_850 : ram_0_73; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1621 = way0_hit ? _GEN_851 : ram_0_74; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1622 = way0_hit ? _GEN_852 : ram_0_75; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1623 = way0_hit ? _GEN_853 : ram_0_76; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1624 = way0_hit ? _GEN_854 : ram_0_77; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1625 = way0_hit ? _GEN_855 : ram_0_78; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1626 = way0_hit ? _GEN_856 : ram_0_79; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1627 = way0_hit ? _GEN_857 : ram_0_80; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1628 = way0_hit ? _GEN_858 : ram_0_81; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1629 = way0_hit ? _GEN_859 : ram_0_82; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1630 = way0_hit ? _GEN_860 : ram_0_83; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1631 = way0_hit ? _GEN_861 : ram_0_84; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1632 = way0_hit ? _GEN_862 : ram_0_85; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1633 = way0_hit ? _GEN_863 : ram_0_86; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1634 = way0_hit ? _GEN_864 : ram_0_87; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1635 = way0_hit ? _GEN_865 : ram_0_88; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1636 = way0_hit ? _GEN_866 : ram_0_89; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1637 = way0_hit ? _GEN_867 : ram_0_90; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1638 = way0_hit ? _GEN_868 : ram_0_91; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1639 = way0_hit ? _GEN_869 : ram_0_92; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1640 = way0_hit ? _GEN_870 : ram_0_93; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1641 = way0_hit ? _GEN_871 : ram_0_94; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1642 = way0_hit ? _GEN_872 : ram_0_95; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1643 = way0_hit ? _GEN_873 : ram_0_96; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1644 = way0_hit ? _GEN_874 : ram_0_97; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1645 = way0_hit ? _GEN_875 : ram_0_98; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1646 = way0_hit ? _GEN_876 : ram_0_99; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1647 = way0_hit ? _GEN_877 : ram_0_100; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1648 = way0_hit ? _GEN_878 : ram_0_101; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1649 = way0_hit ? _GEN_879 : ram_0_102; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1650 = way0_hit ? _GEN_880 : ram_0_103; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1651 = way0_hit ? _GEN_881 : ram_0_104; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1652 = way0_hit ? _GEN_882 : ram_0_105; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1653 = way0_hit ? _GEN_883 : ram_0_106; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1654 = way0_hit ? _GEN_884 : ram_0_107; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1655 = way0_hit ? _GEN_885 : ram_0_108; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1656 = way0_hit ? _GEN_886 : ram_0_109; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1657 = way0_hit ? _GEN_887 : ram_0_110; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1658 = way0_hit ? _GEN_888 : ram_0_111; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1659 = way0_hit ? _GEN_889 : ram_0_112; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1660 = way0_hit ? _GEN_890 : ram_0_113; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1661 = way0_hit ? _GEN_891 : ram_0_114; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1662 = way0_hit ? _GEN_892 : ram_0_115; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1663 = way0_hit ? _GEN_893 : ram_0_116; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1664 = way0_hit ? _GEN_894 : ram_0_117; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1665 = way0_hit ? _GEN_895 : ram_0_118; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1666 = way0_hit ? _GEN_896 : ram_0_119; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1667 = way0_hit ? _GEN_897 : ram_0_120; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1668 = way0_hit ? _GEN_898 : ram_0_121; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1669 = way0_hit ? _GEN_899 : ram_0_122; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1670 = way0_hit ? _GEN_900 : ram_0_123; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1671 = way0_hit ? _GEN_901 : ram_0_124; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1672 = way0_hit ? _GEN_902 : ram_0_125; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1673 = way0_hit ? _GEN_903 : ram_0_126; // @[d_cache.scala 18:24 90:27]
  wire [63:0] _GEN_1674 = way0_hit ? _GEN_904 : ram_0_127; // @[d_cache.scala 18:24 90:27]
  wire  _GEN_1675 = way0_hit ? _GEN_905 : dirty_0_0; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1676 = way0_hit ? _GEN_906 : dirty_0_1; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1677 = way0_hit ? _GEN_907 : dirty_0_2; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1678 = way0_hit ? _GEN_908 : dirty_0_3; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1679 = way0_hit ? _GEN_909 : dirty_0_4; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1680 = way0_hit ? _GEN_910 : dirty_0_5; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1681 = way0_hit ? _GEN_911 : dirty_0_6; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1682 = way0_hit ? _GEN_912 : dirty_0_7; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1683 = way0_hit ? _GEN_913 : dirty_0_8; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1684 = way0_hit ? _GEN_914 : dirty_0_9; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1685 = way0_hit ? _GEN_915 : dirty_0_10; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1686 = way0_hit ? _GEN_916 : dirty_0_11; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1687 = way0_hit ? _GEN_917 : dirty_0_12; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1688 = way0_hit ? _GEN_918 : dirty_0_13; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1689 = way0_hit ? _GEN_919 : dirty_0_14; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1690 = way0_hit ? _GEN_920 : dirty_0_15; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1691 = way0_hit ? _GEN_921 : dirty_0_16; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1692 = way0_hit ? _GEN_922 : dirty_0_17; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1693 = way0_hit ? _GEN_923 : dirty_0_18; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1694 = way0_hit ? _GEN_924 : dirty_0_19; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1695 = way0_hit ? _GEN_925 : dirty_0_20; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1696 = way0_hit ? _GEN_926 : dirty_0_21; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1697 = way0_hit ? _GEN_927 : dirty_0_22; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1698 = way0_hit ? _GEN_928 : dirty_0_23; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1699 = way0_hit ? _GEN_929 : dirty_0_24; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1700 = way0_hit ? _GEN_930 : dirty_0_25; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1701 = way0_hit ? _GEN_931 : dirty_0_26; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1702 = way0_hit ? _GEN_932 : dirty_0_27; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1703 = way0_hit ? _GEN_933 : dirty_0_28; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1704 = way0_hit ? _GEN_934 : dirty_0_29; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1705 = way0_hit ? _GEN_935 : dirty_0_30; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1706 = way0_hit ? _GEN_936 : dirty_0_31; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1707 = way0_hit ? _GEN_937 : dirty_0_32; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1708 = way0_hit ? _GEN_938 : dirty_0_33; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1709 = way0_hit ? _GEN_939 : dirty_0_34; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1710 = way0_hit ? _GEN_940 : dirty_0_35; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1711 = way0_hit ? _GEN_941 : dirty_0_36; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1712 = way0_hit ? _GEN_942 : dirty_0_37; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1713 = way0_hit ? _GEN_943 : dirty_0_38; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1714 = way0_hit ? _GEN_944 : dirty_0_39; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1715 = way0_hit ? _GEN_945 : dirty_0_40; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1716 = way0_hit ? _GEN_946 : dirty_0_41; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1717 = way0_hit ? _GEN_947 : dirty_0_42; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1718 = way0_hit ? _GEN_948 : dirty_0_43; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1719 = way0_hit ? _GEN_949 : dirty_0_44; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1720 = way0_hit ? _GEN_950 : dirty_0_45; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1721 = way0_hit ? _GEN_951 : dirty_0_46; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1722 = way0_hit ? _GEN_952 : dirty_0_47; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1723 = way0_hit ? _GEN_953 : dirty_0_48; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1724 = way0_hit ? _GEN_954 : dirty_0_49; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1725 = way0_hit ? _GEN_955 : dirty_0_50; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1726 = way0_hit ? _GEN_956 : dirty_0_51; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1727 = way0_hit ? _GEN_957 : dirty_0_52; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1728 = way0_hit ? _GEN_958 : dirty_0_53; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1729 = way0_hit ? _GEN_959 : dirty_0_54; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1730 = way0_hit ? _GEN_960 : dirty_0_55; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1731 = way0_hit ? _GEN_961 : dirty_0_56; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1732 = way0_hit ? _GEN_962 : dirty_0_57; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1733 = way0_hit ? _GEN_963 : dirty_0_58; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1734 = way0_hit ? _GEN_964 : dirty_0_59; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1735 = way0_hit ? _GEN_965 : dirty_0_60; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1736 = way0_hit ? _GEN_966 : dirty_0_61; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1737 = way0_hit ? _GEN_967 : dirty_0_62; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1738 = way0_hit ? _GEN_968 : dirty_0_63; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1739 = way0_hit ? _GEN_969 : dirty_0_64; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1740 = way0_hit ? _GEN_970 : dirty_0_65; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1741 = way0_hit ? _GEN_971 : dirty_0_66; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1742 = way0_hit ? _GEN_972 : dirty_0_67; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1743 = way0_hit ? _GEN_973 : dirty_0_68; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1744 = way0_hit ? _GEN_974 : dirty_0_69; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1745 = way0_hit ? _GEN_975 : dirty_0_70; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1746 = way0_hit ? _GEN_976 : dirty_0_71; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1747 = way0_hit ? _GEN_977 : dirty_0_72; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1748 = way0_hit ? _GEN_978 : dirty_0_73; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1749 = way0_hit ? _GEN_979 : dirty_0_74; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1750 = way0_hit ? _GEN_980 : dirty_0_75; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1751 = way0_hit ? _GEN_981 : dirty_0_76; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1752 = way0_hit ? _GEN_982 : dirty_0_77; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1753 = way0_hit ? _GEN_983 : dirty_0_78; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1754 = way0_hit ? _GEN_984 : dirty_0_79; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1755 = way0_hit ? _GEN_985 : dirty_0_80; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1756 = way0_hit ? _GEN_986 : dirty_0_81; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1757 = way0_hit ? _GEN_987 : dirty_0_82; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1758 = way0_hit ? _GEN_988 : dirty_0_83; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1759 = way0_hit ? _GEN_989 : dirty_0_84; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1760 = way0_hit ? _GEN_990 : dirty_0_85; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1761 = way0_hit ? _GEN_991 : dirty_0_86; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1762 = way0_hit ? _GEN_992 : dirty_0_87; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1763 = way0_hit ? _GEN_993 : dirty_0_88; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1764 = way0_hit ? _GEN_994 : dirty_0_89; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1765 = way0_hit ? _GEN_995 : dirty_0_90; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1766 = way0_hit ? _GEN_996 : dirty_0_91; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1767 = way0_hit ? _GEN_997 : dirty_0_92; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1768 = way0_hit ? _GEN_998 : dirty_0_93; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1769 = way0_hit ? _GEN_999 : dirty_0_94; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1770 = way0_hit ? _GEN_1000 : dirty_0_95; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1771 = way0_hit ? _GEN_1001 : dirty_0_96; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1772 = way0_hit ? _GEN_1002 : dirty_0_97; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1773 = way0_hit ? _GEN_1003 : dirty_0_98; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1774 = way0_hit ? _GEN_1004 : dirty_0_99; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1775 = way0_hit ? _GEN_1005 : dirty_0_100; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1776 = way0_hit ? _GEN_1006 : dirty_0_101; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1777 = way0_hit ? _GEN_1007 : dirty_0_102; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1778 = way0_hit ? _GEN_1008 : dirty_0_103; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1779 = way0_hit ? _GEN_1009 : dirty_0_104; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1780 = way0_hit ? _GEN_1010 : dirty_0_105; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1781 = way0_hit ? _GEN_1011 : dirty_0_106; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1782 = way0_hit ? _GEN_1012 : dirty_0_107; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1783 = way0_hit ? _GEN_1013 : dirty_0_108; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1784 = way0_hit ? _GEN_1014 : dirty_0_109; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1785 = way0_hit ? _GEN_1015 : dirty_0_110; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1786 = way0_hit ? _GEN_1016 : dirty_0_111; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1787 = way0_hit ? _GEN_1017 : dirty_0_112; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1788 = way0_hit ? _GEN_1018 : dirty_0_113; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1789 = way0_hit ? _GEN_1019 : dirty_0_114; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1790 = way0_hit ? _GEN_1020 : dirty_0_115; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1791 = way0_hit ? _GEN_1021 : dirty_0_116; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1792 = way0_hit ? _GEN_1022 : dirty_0_117; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1793 = way0_hit ? _GEN_1023 : dirty_0_118; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1794 = way0_hit ? _GEN_1024 : dirty_0_119; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1795 = way0_hit ? _GEN_1025 : dirty_0_120; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1796 = way0_hit ? _GEN_1026 : dirty_0_121; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1797 = way0_hit ? _GEN_1027 : dirty_0_122; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1798 = way0_hit ? _GEN_1028 : dirty_0_123; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1799 = way0_hit ? _GEN_1029 : dirty_0_124; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1800 = way0_hit ? _GEN_1030 : dirty_0_125; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1801 = way0_hit ? _GEN_1031 : dirty_0_126; // @[d_cache.scala 24:26 90:27]
  wire  _GEN_1802 = way0_hit ? _GEN_1032 : dirty_0_127; // @[d_cache.scala 24:26 90:27]
  wire [63:0] _GEN_1803 = way0_hit ? ram_1_0 : _GEN_1290; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1804 = way0_hit ? ram_1_1 : _GEN_1291; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1805 = way0_hit ? ram_1_2 : _GEN_1292; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1806 = way0_hit ? ram_1_3 : _GEN_1293; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1807 = way0_hit ? ram_1_4 : _GEN_1294; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1808 = way0_hit ? ram_1_5 : _GEN_1295; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1809 = way0_hit ? ram_1_6 : _GEN_1296; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1810 = way0_hit ? ram_1_7 : _GEN_1297; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1811 = way0_hit ? ram_1_8 : _GEN_1298; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1812 = way0_hit ? ram_1_9 : _GEN_1299; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1813 = way0_hit ? ram_1_10 : _GEN_1300; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1814 = way0_hit ? ram_1_11 : _GEN_1301; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1815 = way0_hit ? ram_1_12 : _GEN_1302; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1816 = way0_hit ? ram_1_13 : _GEN_1303; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1817 = way0_hit ? ram_1_14 : _GEN_1304; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1818 = way0_hit ? ram_1_15 : _GEN_1305; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1819 = way0_hit ? ram_1_16 : _GEN_1306; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1820 = way0_hit ? ram_1_17 : _GEN_1307; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1821 = way0_hit ? ram_1_18 : _GEN_1308; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1822 = way0_hit ? ram_1_19 : _GEN_1309; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1823 = way0_hit ? ram_1_20 : _GEN_1310; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1824 = way0_hit ? ram_1_21 : _GEN_1311; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1825 = way0_hit ? ram_1_22 : _GEN_1312; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1826 = way0_hit ? ram_1_23 : _GEN_1313; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1827 = way0_hit ? ram_1_24 : _GEN_1314; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1828 = way0_hit ? ram_1_25 : _GEN_1315; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1829 = way0_hit ? ram_1_26 : _GEN_1316; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1830 = way0_hit ? ram_1_27 : _GEN_1317; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1831 = way0_hit ? ram_1_28 : _GEN_1318; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1832 = way0_hit ? ram_1_29 : _GEN_1319; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1833 = way0_hit ? ram_1_30 : _GEN_1320; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1834 = way0_hit ? ram_1_31 : _GEN_1321; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1835 = way0_hit ? ram_1_32 : _GEN_1322; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1836 = way0_hit ? ram_1_33 : _GEN_1323; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1837 = way0_hit ? ram_1_34 : _GEN_1324; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1838 = way0_hit ? ram_1_35 : _GEN_1325; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1839 = way0_hit ? ram_1_36 : _GEN_1326; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1840 = way0_hit ? ram_1_37 : _GEN_1327; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1841 = way0_hit ? ram_1_38 : _GEN_1328; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1842 = way0_hit ? ram_1_39 : _GEN_1329; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1843 = way0_hit ? ram_1_40 : _GEN_1330; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1844 = way0_hit ? ram_1_41 : _GEN_1331; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1845 = way0_hit ? ram_1_42 : _GEN_1332; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1846 = way0_hit ? ram_1_43 : _GEN_1333; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1847 = way0_hit ? ram_1_44 : _GEN_1334; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1848 = way0_hit ? ram_1_45 : _GEN_1335; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1849 = way0_hit ? ram_1_46 : _GEN_1336; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1850 = way0_hit ? ram_1_47 : _GEN_1337; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1851 = way0_hit ? ram_1_48 : _GEN_1338; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1852 = way0_hit ? ram_1_49 : _GEN_1339; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1853 = way0_hit ? ram_1_50 : _GEN_1340; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1854 = way0_hit ? ram_1_51 : _GEN_1341; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1855 = way0_hit ? ram_1_52 : _GEN_1342; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1856 = way0_hit ? ram_1_53 : _GEN_1343; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1857 = way0_hit ? ram_1_54 : _GEN_1344; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1858 = way0_hit ? ram_1_55 : _GEN_1345; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1859 = way0_hit ? ram_1_56 : _GEN_1346; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1860 = way0_hit ? ram_1_57 : _GEN_1347; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1861 = way0_hit ? ram_1_58 : _GEN_1348; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1862 = way0_hit ? ram_1_59 : _GEN_1349; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1863 = way0_hit ? ram_1_60 : _GEN_1350; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1864 = way0_hit ? ram_1_61 : _GEN_1351; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1865 = way0_hit ? ram_1_62 : _GEN_1352; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1866 = way0_hit ? ram_1_63 : _GEN_1353; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1867 = way0_hit ? ram_1_64 : _GEN_1354; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1868 = way0_hit ? ram_1_65 : _GEN_1355; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1869 = way0_hit ? ram_1_66 : _GEN_1356; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1870 = way0_hit ? ram_1_67 : _GEN_1357; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1871 = way0_hit ? ram_1_68 : _GEN_1358; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1872 = way0_hit ? ram_1_69 : _GEN_1359; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1873 = way0_hit ? ram_1_70 : _GEN_1360; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1874 = way0_hit ? ram_1_71 : _GEN_1361; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1875 = way0_hit ? ram_1_72 : _GEN_1362; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1876 = way0_hit ? ram_1_73 : _GEN_1363; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1877 = way0_hit ? ram_1_74 : _GEN_1364; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1878 = way0_hit ? ram_1_75 : _GEN_1365; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1879 = way0_hit ? ram_1_76 : _GEN_1366; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1880 = way0_hit ? ram_1_77 : _GEN_1367; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1881 = way0_hit ? ram_1_78 : _GEN_1368; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1882 = way0_hit ? ram_1_79 : _GEN_1369; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1883 = way0_hit ? ram_1_80 : _GEN_1370; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1884 = way0_hit ? ram_1_81 : _GEN_1371; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1885 = way0_hit ? ram_1_82 : _GEN_1372; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1886 = way0_hit ? ram_1_83 : _GEN_1373; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1887 = way0_hit ? ram_1_84 : _GEN_1374; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1888 = way0_hit ? ram_1_85 : _GEN_1375; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1889 = way0_hit ? ram_1_86 : _GEN_1376; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1890 = way0_hit ? ram_1_87 : _GEN_1377; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1891 = way0_hit ? ram_1_88 : _GEN_1378; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1892 = way0_hit ? ram_1_89 : _GEN_1379; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1893 = way0_hit ? ram_1_90 : _GEN_1380; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1894 = way0_hit ? ram_1_91 : _GEN_1381; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1895 = way0_hit ? ram_1_92 : _GEN_1382; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1896 = way0_hit ? ram_1_93 : _GEN_1383; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1897 = way0_hit ? ram_1_94 : _GEN_1384; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1898 = way0_hit ? ram_1_95 : _GEN_1385; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1899 = way0_hit ? ram_1_96 : _GEN_1386; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1900 = way0_hit ? ram_1_97 : _GEN_1387; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1901 = way0_hit ? ram_1_98 : _GEN_1388; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1902 = way0_hit ? ram_1_99 : _GEN_1389; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1903 = way0_hit ? ram_1_100 : _GEN_1390; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1904 = way0_hit ? ram_1_101 : _GEN_1391; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1905 = way0_hit ? ram_1_102 : _GEN_1392; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1906 = way0_hit ? ram_1_103 : _GEN_1393; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1907 = way0_hit ? ram_1_104 : _GEN_1394; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1908 = way0_hit ? ram_1_105 : _GEN_1395; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1909 = way0_hit ? ram_1_106 : _GEN_1396; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1910 = way0_hit ? ram_1_107 : _GEN_1397; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1911 = way0_hit ? ram_1_108 : _GEN_1398; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1912 = way0_hit ? ram_1_109 : _GEN_1399; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1913 = way0_hit ? ram_1_110 : _GEN_1400; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1914 = way0_hit ? ram_1_111 : _GEN_1401; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1915 = way0_hit ? ram_1_112 : _GEN_1402; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1916 = way0_hit ? ram_1_113 : _GEN_1403; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1917 = way0_hit ? ram_1_114 : _GEN_1404; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1918 = way0_hit ? ram_1_115 : _GEN_1405; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1919 = way0_hit ? ram_1_116 : _GEN_1406; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1920 = way0_hit ? ram_1_117 : _GEN_1407; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1921 = way0_hit ? ram_1_118 : _GEN_1408; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1922 = way0_hit ? ram_1_119 : _GEN_1409; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1923 = way0_hit ? ram_1_120 : _GEN_1410; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1924 = way0_hit ? ram_1_121 : _GEN_1411; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1925 = way0_hit ? ram_1_122 : _GEN_1412; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1926 = way0_hit ? ram_1_123 : _GEN_1413; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1927 = way0_hit ? ram_1_124 : _GEN_1414; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1928 = way0_hit ? ram_1_125 : _GEN_1415; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1929 = way0_hit ? ram_1_126 : _GEN_1416; // @[d_cache.scala 19:24 90:27]
  wire [63:0] _GEN_1930 = way0_hit ? ram_1_127 : _GEN_1417; // @[d_cache.scala 19:24 90:27]
  wire  _GEN_1931 = way0_hit ? dirty_1_0 : _GEN_1418; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1932 = way0_hit ? dirty_1_1 : _GEN_1419; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1933 = way0_hit ? dirty_1_2 : _GEN_1420; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1934 = way0_hit ? dirty_1_3 : _GEN_1421; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1935 = way0_hit ? dirty_1_4 : _GEN_1422; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1936 = way0_hit ? dirty_1_5 : _GEN_1423; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1937 = way0_hit ? dirty_1_6 : _GEN_1424; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1938 = way0_hit ? dirty_1_7 : _GEN_1425; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1939 = way0_hit ? dirty_1_8 : _GEN_1426; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1940 = way0_hit ? dirty_1_9 : _GEN_1427; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1941 = way0_hit ? dirty_1_10 : _GEN_1428; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1942 = way0_hit ? dirty_1_11 : _GEN_1429; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1943 = way0_hit ? dirty_1_12 : _GEN_1430; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1944 = way0_hit ? dirty_1_13 : _GEN_1431; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1945 = way0_hit ? dirty_1_14 : _GEN_1432; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1946 = way0_hit ? dirty_1_15 : _GEN_1433; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1947 = way0_hit ? dirty_1_16 : _GEN_1434; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1948 = way0_hit ? dirty_1_17 : _GEN_1435; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1949 = way0_hit ? dirty_1_18 : _GEN_1436; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1950 = way0_hit ? dirty_1_19 : _GEN_1437; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1951 = way0_hit ? dirty_1_20 : _GEN_1438; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1952 = way0_hit ? dirty_1_21 : _GEN_1439; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1953 = way0_hit ? dirty_1_22 : _GEN_1440; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1954 = way0_hit ? dirty_1_23 : _GEN_1441; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1955 = way0_hit ? dirty_1_24 : _GEN_1442; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1956 = way0_hit ? dirty_1_25 : _GEN_1443; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1957 = way0_hit ? dirty_1_26 : _GEN_1444; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1958 = way0_hit ? dirty_1_27 : _GEN_1445; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1959 = way0_hit ? dirty_1_28 : _GEN_1446; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1960 = way0_hit ? dirty_1_29 : _GEN_1447; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1961 = way0_hit ? dirty_1_30 : _GEN_1448; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1962 = way0_hit ? dirty_1_31 : _GEN_1449; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1963 = way0_hit ? dirty_1_32 : _GEN_1450; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1964 = way0_hit ? dirty_1_33 : _GEN_1451; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1965 = way0_hit ? dirty_1_34 : _GEN_1452; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1966 = way0_hit ? dirty_1_35 : _GEN_1453; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1967 = way0_hit ? dirty_1_36 : _GEN_1454; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1968 = way0_hit ? dirty_1_37 : _GEN_1455; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1969 = way0_hit ? dirty_1_38 : _GEN_1456; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1970 = way0_hit ? dirty_1_39 : _GEN_1457; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1971 = way0_hit ? dirty_1_40 : _GEN_1458; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1972 = way0_hit ? dirty_1_41 : _GEN_1459; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1973 = way0_hit ? dirty_1_42 : _GEN_1460; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1974 = way0_hit ? dirty_1_43 : _GEN_1461; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1975 = way0_hit ? dirty_1_44 : _GEN_1462; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1976 = way0_hit ? dirty_1_45 : _GEN_1463; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1977 = way0_hit ? dirty_1_46 : _GEN_1464; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1978 = way0_hit ? dirty_1_47 : _GEN_1465; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1979 = way0_hit ? dirty_1_48 : _GEN_1466; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1980 = way0_hit ? dirty_1_49 : _GEN_1467; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1981 = way0_hit ? dirty_1_50 : _GEN_1468; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1982 = way0_hit ? dirty_1_51 : _GEN_1469; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1983 = way0_hit ? dirty_1_52 : _GEN_1470; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1984 = way0_hit ? dirty_1_53 : _GEN_1471; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1985 = way0_hit ? dirty_1_54 : _GEN_1472; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1986 = way0_hit ? dirty_1_55 : _GEN_1473; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1987 = way0_hit ? dirty_1_56 : _GEN_1474; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1988 = way0_hit ? dirty_1_57 : _GEN_1475; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1989 = way0_hit ? dirty_1_58 : _GEN_1476; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1990 = way0_hit ? dirty_1_59 : _GEN_1477; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1991 = way0_hit ? dirty_1_60 : _GEN_1478; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1992 = way0_hit ? dirty_1_61 : _GEN_1479; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1993 = way0_hit ? dirty_1_62 : _GEN_1480; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1994 = way0_hit ? dirty_1_63 : _GEN_1481; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1995 = way0_hit ? dirty_1_64 : _GEN_1482; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1996 = way0_hit ? dirty_1_65 : _GEN_1483; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1997 = way0_hit ? dirty_1_66 : _GEN_1484; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1998 = way0_hit ? dirty_1_67 : _GEN_1485; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_1999 = way0_hit ? dirty_1_68 : _GEN_1486; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2000 = way0_hit ? dirty_1_69 : _GEN_1487; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2001 = way0_hit ? dirty_1_70 : _GEN_1488; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2002 = way0_hit ? dirty_1_71 : _GEN_1489; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2003 = way0_hit ? dirty_1_72 : _GEN_1490; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2004 = way0_hit ? dirty_1_73 : _GEN_1491; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2005 = way0_hit ? dirty_1_74 : _GEN_1492; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2006 = way0_hit ? dirty_1_75 : _GEN_1493; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2007 = way0_hit ? dirty_1_76 : _GEN_1494; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2008 = way0_hit ? dirty_1_77 : _GEN_1495; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2009 = way0_hit ? dirty_1_78 : _GEN_1496; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2010 = way0_hit ? dirty_1_79 : _GEN_1497; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2011 = way0_hit ? dirty_1_80 : _GEN_1498; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2012 = way0_hit ? dirty_1_81 : _GEN_1499; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2013 = way0_hit ? dirty_1_82 : _GEN_1500; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2014 = way0_hit ? dirty_1_83 : _GEN_1501; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2015 = way0_hit ? dirty_1_84 : _GEN_1502; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2016 = way0_hit ? dirty_1_85 : _GEN_1503; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2017 = way0_hit ? dirty_1_86 : _GEN_1504; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2018 = way0_hit ? dirty_1_87 : _GEN_1505; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2019 = way0_hit ? dirty_1_88 : _GEN_1506; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2020 = way0_hit ? dirty_1_89 : _GEN_1507; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2021 = way0_hit ? dirty_1_90 : _GEN_1508; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2022 = way0_hit ? dirty_1_91 : _GEN_1509; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2023 = way0_hit ? dirty_1_92 : _GEN_1510; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2024 = way0_hit ? dirty_1_93 : _GEN_1511; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2025 = way0_hit ? dirty_1_94 : _GEN_1512; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2026 = way0_hit ? dirty_1_95 : _GEN_1513; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2027 = way0_hit ? dirty_1_96 : _GEN_1514; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2028 = way0_hit ? dirty_1_97 : _GEN_1515; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2029 = way0_hit ? dirty_1_98 : _GEN_1516; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2030 = way0_hit ? dirty_1_99 : _GEN_1517; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2031 = way0_hit ? dirty_1_100 : _GEN_1518; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2032 = way0_hit ? dirty_1_101 : _GEN_1519; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2033 = way0_hit ? dirty_1_102 : _GEN_1520; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2034 = way0_hit ? dirty_1_103 : _GEN_1521; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2035 = way0_hit ? dirty_1_104 : _GEN_1522; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2036 = way0_hit ? dirty_1_105 : _GEN_1523; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2037 = way0_hit ? dirty_1_106 : _GEN_1524; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2038 = way0_hit ? dirty_1_107 : _GEN_1525; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2039 = way0_hit ? dirty_1_108 : _GEN_1526; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2040 = way0_hit ? dirty_1_109 : _GEN_1527; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2041 = way0_hit ? dirty_1_110 : _GEN_1528; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2042 = way0_hit ? dirty_1_111 : _GEN_1529; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2043 = way0_hit ? dirty_1_112 : _GEN_1530; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2044 = way0_hit ? dirty_1_113 : _GEN_1531; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2045 = way0_hit ? dirty_1_114 : _GEN_1532; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2046 = way0_hit ? dirty_1_115 : _GEN_1533; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2047 = way0_hit ? dirty_1_116 : _GEN_1534; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2048 = way0_hit ? dirty_1_117 : _GEN_1535; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2049 = way0_hit ? dirty_1_118 : _GEN_1536; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2050 = way0_hit ? dirty_1_119 : _GEN_1537; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2051 = way0_hit ? dirty_1_120 : _GEN_1538; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2052 = way0_hit ? dirty_1_121 : _GEN_1539; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2053 = way0_hit ? dirty_1_122 : _GEN_1540; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2054 = way0_hit ? dirty_1_123 : _GEN_1541; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2055 = way0_hit ? dirty_1_124 : _GEN_1542; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2056 = way0_hit ? dirty_1_125 : _GEN_1543; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2057 = way0_hit ? dirty_1_126 : _GEN_1544; // @[d_cache.scala 25:26 90:27]
  wire  _GEN_2058 = way0_hit ? dirty_1_127 : _GEN_1545; // @[d_cache.scala 25:26 90:27]
  wire [2:0] _GEN_2059 = io_from_axi_rvalid ? 3'h5 : state; // @[d_cache.scala 106:37 107:23 60:24]
  wire [63:0] _GEN_2060 = io_from_axi_rvalid ? io_from_axi_rdata : receive_data; // @[d_cache.scala 109:37 110:30 34:31]
  wire [2:0] _GEN_2061 = io_from_axi_bvalid ? 3'h0 : state; // @[d_cache.scala 114:37 115:23 60:24]
  wire [63:0] _GEN_2062 = 7'h0 == index ? receive_data : ram_0_0; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2063 = 7'h1 == index ? receive_data : ram_0_1; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2064 = 7'h2 == index ? receive_data : ram_0_2; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2065 = 7'h3 == index ? receive_data : ram_0_3; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2066 = 7'h4 == index ? receive_data : ram_0_4; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2067 = 7'h5 == index ? receive_data : ram_0_5; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2068 = 7'h6 == index ? receive_data : ram_0_6; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2069 = 7'h7 == index ? receive_data : ram_0_7; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2070 = 7'h8 == index ? receive_data : ram_0_8; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2071 = 7'h9 == index ? receive_data : ram_0_9; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2072 = 7'ha == index ? receive_data : ram_0_10; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2073 = 7'hb == index ? receive_data : ram_0_11; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2074 = 7'hc == index ? receive_data : ram_0_12; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2075 = 7'hd == index ? receive_data : ram_0_13; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2076 = 7'he == index ? receive_data : ram_0_14; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2077 = 7'hf == index ? receive_data : ram_0_15; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2078 = 7'h10 == index ? receive_data : ram_0_16; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2079 = 7'h11 == index ? receive_data : ram_0_17; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2080 = 7'h12 == index ? receive_data : ram_0_18; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2081 = 7'h13 == index ? receive_data : ram_0_19; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2082 = 7'h14 == index ? receive_data : ram_0_20; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2083 = 7'h15 == index ? receive_data : ram_0_21; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2084 = 7'h16 == index ? receive_data : ram_0_22; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2085 = 7'h17 == index ? receive_data : ram_0_23; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2086 = 7'h18 == index ? receive_data : ram_0_24; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2087 = 7'h19 == index ? receive_data : ram_0_25; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2088 = 7'h1a == index ? receive_data : ram_0_26; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2089 = 7'h1b == index ? receive_data : ram_0_27; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2090 = 7'h1c == index ? receive_data : ram_0_28; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2091 = 7'h1d == index ? receive_data : ram_0_29; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2092 = 7'h1e == index ? receive_data : ram_0_30; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2093 = 7'h1f == index ? receive_data : ram_0_31; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2094 = 7'h20 == index ? receive_data : ram_0_32; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2095 = 7'h21 == index ? receive_data : ram_0_33; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2096 = 7'h22 == index ? receive_data : ram_0_34; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2097 = 7'h23 == index ? receive_data : ram_0_35; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2098 = 7'h24 == index ? receive_data : ram_0_36; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2099 = 7'h25 == index ? receive_data : ram_0_37; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2100 = 7'h26 == index ? receive_data : ram_0_38; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2101 = 7'h27 == index ? receive_data : ram_0_39; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2102 = 7'h28 == index ? receive_data : ram_0_40; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2103 = 7'h29 == index ? receive_data : ram_0_41; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2104 = 7'h2a == index ? receive_data : ram_0_42; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2105 = 7'h2b == index ? receive_data : ram_0_43; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2106 = 7'h2c == index ? receive_data : ram_0_44; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2107 = 7'h2d == index ? receive_data : ram_0_45; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2108 = 7'h2e == index ? receive_data : ram_0_46; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2109 = 7'h2f == index ? receive_data : ram_0_47; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2110 = 7'h30 == index ? receive_data : ram_0_48; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2111 = 7'h31 == index ? receive_data : ram_0_49; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2112 = 7'h32 == index ? receive_data : ram_0_50; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2113 = 7'h33 == index ? receive_data : ram_0_51; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2114 = 7'h34 == index ? receive_data : ram_0_52; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2115 = 7'h35 == index ? receive_data : ram_0_53; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2116 = 7'h36 == index ? receive_data : ram_0_54; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2117 = 7'h37 == index ? receive_data : ram_0_55; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2118 = 7'h38 == index ? receive_data : ram_0_56; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2119 = 7'h39 == index ? receive_data : ram_0_57; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2120 = 7'h3a == index ? receive_data : ram_0_58; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2121 = 7'h3b == index ? receive_data : ram_0_59; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2122 = 7'h3c == index ? receive_data : ram_0_60; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2123 = 7'h3d == index ? receive_data : ram_0_61; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2124 = 7'h3e == index ? receive_data : ram_0_62; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2125 = 7'h3f == index ? receive_data : ram_0_63; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2126 = 7'h40 == index ? receive_data : ram_0_64; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2127 = 7'h41 == index ? receive_data : ram_0_65; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2128 = 7'h42 == index ? receive_data : ram_0_66; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2129 = 7'h43 == index ? receive_data : ram_0_67; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2130 = 7'h44 == index ? receive_data : ram_0_68; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2131 = 7'h45 == index ? receive_data : ram_0_69; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2132 = 7'h46 == index ? receive_data : ram_0_70; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2133 = 7'h47 == index ? receive_data : ram_0_71; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2134 = 7'h48 == index ? receive_data : ram_0_72; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2135 = 7'h49 == index ? receive_data : ram_0_73; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2136 = 7'h4a == index ? receive_data : ram_0_74; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2137 = 7'h4b == index ? receive_data : ram_0_75; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2138 = 7'h4c == index ? receive_data : ram_0_76; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2139 = 7'h4d == index ? receive_data : ram_0_77; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2140 = 7'h4e == index ? receive_data : ram_0_78; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2141 = 7'h4f == index ? receive_data : ram_0_79; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2142 = 7'h50 == index ? receive_data : ram_0_80; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2143 = 7'h51 == index ? receive_data : ram_0_81; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2144 = 7'h52 == index ? receive_data : ram_0_82; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2145 = 7'h53 == index ? receive_data : ram_0_83; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2146 = 7'h54 == index ? receive_data : ram_0_84; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2147 = 7'h55 == index ? receive_data : ram_0_85; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2148 = 7'h56 == index ? receive_data : ram_0_86; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2149 = 7'h57 == index ? receive_data : ram_0_87; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2150 = 7'h58 == index ? receive_data : ram_0_88; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2151 = 7'h59 == index ? receive_data : ram_0_89; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2152 = 7'h5a == index ? receive_data : ram_0_90; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2153 = 7'h5b == index ? receive_data : ram_0_91; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2154 = 7'h5c == index ? receive_data : ram_0_92; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2155 = 7'h5d == index ? receive_data : ram_0_93; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2156 = 7'h5e == index ? receive_data : ram_0_94; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2157 = 7'h5f == index ? receive_data : ram_0_95; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2158 = 7'h60 == index ? receive_data : ram_0_96; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2159 = 7'h61 == index ? receive_data : ram_0_97; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2160 = 7'h62 == index ? receive_data : ram_0_98; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2161 = 7'h63 == index ? receive_data : ram_0_99; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2162 = 7'h64 == index ? receive_data : ram_0_100; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2163 = 7'h65 == index ? receive_data : ram_0_101; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2164 = 7'h66 == index ? receive_data : ram_0_102; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2165 = 7'h67 == index ? receive_data : ram_0_103; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2166 = 7'h68 == index ? receive_data : ram_0_104; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2167 = 7'h69 == index ? receive_data : ram_0_105; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2168 = 7'h6a == index ? receive_data : ram_0_106; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2169 = 7'h6b == index ? receive_data : ram_0_107; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2170 = 7'h6c == index ? receive_data : ram_0_108; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2171 = 7'h6d == index ? receive_data : ram_0_109; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2172 = 7'h6e == index ? receive_data : ram_0_110; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2173 = 7'h6f == index ? receive_data : ram_0_111; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2174 = 7'h70 == index ? receive_data : ram_0_112; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2175 = 7'h71 == index ? receive_data : ram_0_113; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2176 = 7'h72 == index ? receive_data : ram_0_114; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2177 = 7'h73 == index ? receive_data : ram_0_115; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2178 = 7'h74 == index ? receive_data : ram_0_116; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2179 = 7'h75 == index ? receive_data : ram_0_117; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2180 = 7'h76 == index ? receive_data : ram_0_118; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2181 = 7'h77 == index ? receive_data : ram_0_119; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2182 = 7'h78 == index ? receive_data : ram_0_120; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2183 = 7'h79 == index ? receive_data : ram_0_121; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2184 = 7'h7a == index ? receive_data : ram_0_122; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2185 = 7'h7b == index ? receive_data : ram_0_123; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2186 = 7'h7c == index ? receive_data : ram_0_124; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2187 = 7'h7d == index ? receive_data : ram_0_125; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2188 = 7'h7e == index ? receive_data : ram_0_126; // @[d_cache.scala 121:{30,30} 18:24]
  wire [63:0] _GEN_2189 = 7'h7f == index ? receive_data : ram_0_127; // @[d_cache.scala 121:{30,30} 18:24]
  wire [31:0] _GEN_2190 = 7'h0 == index ? _GEN_15265 : tag_0_0; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2191 = 7'h1 == index ? _GEN_15265 : tag_0_1; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2192 = 7'h2 == index ? _GEN_15265 : tag_0_2; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2193 = 7'h3 == index ? _GEN_15265 : tag_0_3; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2194 = 7'h4 == index ? _GEN_15265 : tag_0_4; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2195 = 7'h5 == index ? _GEN_15265 : tag_0_5; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2196 = 7'h6 == index ? _GEN_15265 : tag_0_6; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2197 = 7'h7 == index ? _GEN_15265 : tag_0_7; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2198 = 7'h8 == index ? _GEN_15265 : tag_0_8; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2199 = 7'h9 == index ? _GEN_15265 : tag_0_9; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2200 = 7'ha == index ? _GEN_15265 : tag_0_10; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2201 = 7'hb == index ? _GEN_15265 : tag_0_11; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2202 = 7'hc == index ? _GEN_15265 : tag_0_12; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2203 = 7'hd == index ? _GEN_15265 : tag_0_13; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2204 = 7'he == index ? _GEN_15265 : tag_0_14; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2205 = 7'hf == index ? _GEN_15265 : tag_0_15; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2206 = 7'h10 == index ? _GEN_15265 : tag_0_16; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2207 = 7'h11 == index ? _GEN_15265 : tag_0_17; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2208 = 7'h12 == index ? _GEN_15265 : tag_0_18; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2209 = 7'h13 == index ? _GEN_15265 : tag_0_19; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2210 = 7'h14 == index ? _GEN_15265 : tag_0_20; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2211 = 7'h15 == index ? _GEN_15265 : tag_0_21; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2212 = 7'h16 == index ? _GEN_15265 : tag_0_22; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2213 = 7'h17 == index ? _GEN_15265 : tag_0_23; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2214 = 7'h18 == index ? _GEN_15265 : tag_0_24; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2215 = 7'h19 == index ? _GEN_15265 : tag_0_25; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2216 = 7'h1a == index ? _GEN_15265 : tag_0_26; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2217 = 7'h1b == index ? _GEN_15265 : tag_0_27; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2218 = 7'h1c == index ? _GEN_15265 : tag_0_28; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2219 = 7'h1d == index ? _GEN_15265 : tag_0_29; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2220 = 7'h1e == index ? _GEN_15265 : tag_0_30; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2221 = 7'h1f == index ? _GEN_15265 : tag_0_31; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2222 = 7'h20 == index ? _GEN_15265 : tag_0_32; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2223 = 7'h21 == index ? _GEN_15265 : tag_0_33; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2224 = 7'h22 == index ? _GEN_15265 : tag_0_34; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2225 = 7'h23 == index ? _GEN_15265 : tag_0_35; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2226 = 7'h24 == index ? _GEN_15265 : tag_0_36; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2227 = 7'h25 == index ? _GEN_15265 : tag_0_37; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2228 = 7'h26 == index ? _GEN_15265 : tag_0_38; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2229 = 7'h27 == index ? _GEN_15265 : tag_0_39; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2230 = 7'h28 == index ? _GEN_15265 : tag_0_40; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2231 = 7'h29 == index ? _GEN_15265 : tag_0_41; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2232 = 7'h2a == index ? _GEN_15265 : tag_0_42; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2233 = 7'h2b == index ? _GEN_15265 : tag_0_43; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2234 = 7'h2c == index ? _GEN_15265 : tag_0_44; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2235 = 7'h2d == index ? _GEN_15265 : tag_0_45; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2236 = 7'h2e == index ? _GEN_15265 : tag_0_46; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2237 = 7'h2f == index ? _GEN_15265 : tag_0_47; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2238 = 7'h30 == index ? _GEN_15265 : tag_0_48; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2239 = 7'h31 == index ? _GEN_15265 : tag_0_49; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2240 = 7'h32 == index ? _GEN_15265 : tag_0_50; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2241 = 7'h33 == index ? _GEN_15265 : tag_0_51; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2242 = 7'h34 == index ? _GEN_15265 : tag_0_52; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2243 = 7'h35 == index ? _GEN_15265 : tag_0_53; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2244 = 7'h36 == index ? _GEN_15265 : tag_0_54; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2245 = 7'h37 == index ? _GEN_15265 : tag_0_55; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2246 = 7'h38 == index ? _GEN_15265 : tag_0_56; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2247 = 7'h39 == index ? _GEN_15265 : tag_0_57; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2248 = 7'h3a == index ? _GEN_15265 : tag_0_58; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2249 = 7'h3b == index ? _GEN_15265 : tag_0_59; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2250 = 7'h3c == index ? _GEN_15265 : tag_0_60; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2251 = 7'h3d == index ? _GEN_15265 : tag_0_61; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2252 = 7'h3e == index ? _GEN_15265 : tag_0_62; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2253 = 7'h3f == index ? _GEN_15265 : tag_0_63; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2254 = 7'h40 == index ? _GEN_15265 : tag_0_64; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2255 = 7'h41 == index ? _GEN_15265 : tag_0_65; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2256 = 7'h42 == index ? _GEN_15265 : tag_0_66; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2257 = 7'h43 == index ? _GEN_15265 : tag_0_67; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2258 = 7'h44 == index ? _GEN_15265 : tag_0_68; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2259 = 7'h45 == index ? _GEN_15265 : tag_0_69; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2260 = 7'h46 == index ? _GEN_15265 : tag_0_70; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2261 = 7'h47 == index ? _GEN_15265 : tag_0_71; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2262 = 7'h48 == index ? _GEN_15265 : tag_0_72; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2263 = 7'h49 == index ? _GEN_15265 : tag_0_73; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2264 = 7'h4a == index ? _GEN_15265 : tag_0_74; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2265 = 7'h4b == index ? _GEN_15265 : tag_0_75; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2266 = 7'h4c == index ? _GEN_15265 : tag_0_76; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2267 = 7'h4d == index ? _GEN_15265 : tag_0_77; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2268 = 7'h4e == index ? _GEN_15265 : tag_0_78; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2269 = 7'h4f == index ? _GEN_15265 : tag_0_79; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2270 = 7'h50 == index ? _GEN_15265 : tag_0_80; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2271 = 7'h51 == index ? _GEN_15265 : tag_0_81; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2272 = 7'h52 == index ? _GEN_15265 : tag_0_82; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2273 = 7'h53 == index ? _GEN_15265 : tag_0_83; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2274 = 7'h54 == index ? _GEN_15265 : tag_0_84; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2275 = 7'h55 == index ? _GEN_15265 : tag_0_85; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2276 = 7'h56 == index ? _GEN_15265 : tag_0_86; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2277 = 7'h57 == index ? _GEN_15265 : tag_0_87; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2278 = 7'h58 == index ? _GEN_15265 : tag_0_88; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2279 = 7'h59 == index ? _GEN_15265 : tag_0_89; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2280 = 7'h5a == index ? _GEN_15265 : tag_0_90; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2281 = 7'h5b == index ? _GEN_15265 : tag_0_91; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2282 = 7'h5c == index ? _GEN_15265 : tag_0_92; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2283 = 7'h5d == index ? _GEN_15265 : tag_0_93; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2284 = 7'h5e == index ? _GEN_15265 : tag_0_94; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2285 = 7'h5f == index ? _GEN_15265 : tag_0_95; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2286 = 7'h60 == index ? _GEN_15265 : tag_0_96; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2287 = 7'h61 == index ? _GEN_15265 : tag_0_97; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2288 = 7'h62 == index ? _GEN_15265 : tag_0_98; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2289 = 7'h63 == index ? _GEN_15265 : tag_0_99; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2290 = 7'h64 == index ? _GEN_15265 : tag_0_100; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2291 = 7'h65 == index ? _GEN_15265 : tag_0_101; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2292 = 7'h66 == index ? _GEN_15265 : tag_0_102; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2293 = 7'h67 == index ? _GEN_15265 : tag_0_103; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2294 = 7'h68 == index ? _GEN_15265 : tag_0_104; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2295 = 7'h69 == index ? _GEN_15265 : tag_0_105; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2296 = 7'h6a == index ? _GEN_15265 : tag_0_106; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2297 = 7'h6b == index ? _GEN_15265 : tag_0_107; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2298 = 7'h6c == index ? _GEN_15265 : tag_0_108; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2299 = 7'h6d == index ? _GEN_15265 : tag_0_109; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2300 = 7'h6e == index ? _GEN_15265 : tag_0_110; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2301 = 7'h6f == index ? _GEN_15265 : tag_0_111; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2302 = 7'h70 == index ? _GEN_15265 : tag_0_112; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2303 = 7'h71 == index ? _GEN_15265 : tag_0_113; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2304 = 7'h72 == index ? _GEN_15265 : tag_0_114; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2305 = 7'h73 == index ? _GEN_15265 : tag_0_115; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2306 = 7'h74 == index ? _GEN_15265 : tag_0_116; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2307 = 7'h75 == index ? _GEN_15265 : tag_0_117; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2308 = 7'h76 == index ? _GEN_15265 : tag_0_118; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2309 = 7'h77 == index ? _GEN_15265 : tag_0_119; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2310 = 7'h78 == index ? _GEN_15265 : tag_0_120; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2311 = 7'h79 == index ? _GEN_15265 : tag_0_121; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2312 = 7'h7a == index ? _GEN_15265 : tag_0_122; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2313 = 7'h7b == index ? _GEN_15265 : tag_0_123; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2314 = 7'h7c == index ? _GEN_15265 : tag_0_124; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2315 = 7'h7d == index ? _GEN_15265 : tag_0_125; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2316 = 7'h7e == index ? _GEN_15265 : tag_0_126; // @[d_cache.scala 122:{30,30} 20:24]
  wire [31:0] _GEN_2317 = 7'h7f == index ? _GEN_15265 : tag_0_127; // @[d_cache.scala 122:{30,30} 20:24]
  wire  _GEN_2318 = _GEN_15267 | valid_0_0; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2319 = _GEN_15268 | valid_0_1; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2320 = _GEN_15269 | valid_0_2; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2321 = _GEN_15270 | valid_0_3; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2322 = _GEN_15271 | valid_0_4; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2323 = _GEN_15272 | valid_0_5; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2324 = _GEN_15273 | valid_0_6; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2325 = _GEN_15274 | valid_0_7; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2326 = _GEN_15275 | valid_0_8; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2327 = _GEN_15276 | valid_0_9; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2328 = _GEN_15277 | valid_0_10; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2329 = _GEN_15278 | valid_0_11; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2330 = _GEN_15279 | valid_0_12; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2331 = _GEN_15280 | valid_0_13; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2332 = _GEN_15281 | valid_0_14; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2333 = _GEN_15282 | valid_0_15; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2334 = _GEN_15283 | valid_0_16; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2335 = _GEN_15284 | valid_0_17; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2336 = _GEN_15285 | valid_0_18; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2337 = _GEN_15286 | valid_0_19; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2338 = _GEN_15287 | valid_0_20; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2339 = _GEN_15288 | valid_0_21; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2340 = _GEN_15289 | valid_0_22; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2341 = _GEN_15290 | valid_0_23; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2342 = _GEN_15291 | valid_0_24; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2343 = _GEN_15292 | valid_0_25; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2344 = _GEN_15293 | valid_0_26; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2345 = _GEN_15294 | valid_0_27; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2346 = _GEN_15295 | valid_0_28; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2347 = _GEN_15296 | valid_0_29; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2348 = _GEN_15297 | valid_0_30; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2349 = _GEN_15298 | valid_0_31; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2350 = _GEN_15299 | valid_0_32; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2351 = _GEN_15300 | valid_0_33; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2352 = _GEN_15301 | valid_0_34; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2353 = _GEN_15302 | valid_0_35; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2354 = _GEN_15303 | valid_0_36; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2355 = _GEN_15304 | valid_0_37; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2356 = _GEN_15305 | valid_0_38; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2357 = _GEN_15306 | valid_0_39; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2358 = _GEN_15307 | valid_0_40; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2359 = _GEN_15308 | valid_0_41; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2360 = _GEN_15309 | valid_0_42; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2361 = _GEN_15310 | valid_0_43; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2362 = _GEN_15311 | valid_0_44; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2363 = _GEN_15312 | valid_0_45; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2364 = _GEN_15313 | valid_0_46; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2365 = _GEN_15314 | valid_0_47; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2366 = _GEN_15315 | valid_0_48; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2367 = _GEN_15316 | valid_0_49; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2368 = _GEN_15317 | valid_0_50; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2369 = _GEN_15318 | valid_0_51; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2370 = _GEN_15319 | valid_0_52; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2371 = _GEN_15320 | valid_0_53; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2372 = _GEN_15321 | valid_0_54; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2373 = _GEN_15322 | valid_0_55; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2374 = _GEN_15323 | valid_0_56; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2375 = _GEN_15324 | valid_0_57; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2376 = _GEN_15325 | valid_0_58; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2377 = _GEN_15326 | valid_0_59; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2378 = _GEN_15327 | valid_0_60; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2379 = _GEN_15328 | valid_0_61; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2380 = _GEN_15329 | valid_0_62; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2381 = _GEN_15330 | valid_0_63; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2382 = _GEN_15331 | valid_0_64; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2383 = _GEN_15332 | valid_0_65; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2384 = _GEN_15333 | valid_0_66; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2385 = _GEN_15334 | valid_0_67; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2386 = _GEN_15335 | valid_0_68; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2387 = _GEN_15336 | valid_0_69; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2388 = _GEN_15337 | valid_0_70; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2389 = _GEN_15338 | valid_0_71; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2390 = _GEN_15339 | valid_0_72; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2391 = _GEN_15340 | valid_0_73; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2392 = _GEN_15341 | valid_0_74; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2393 = _GEN_15342 | valid_0_75; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2394 = _GEN_15343 | valid_0_76; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2395 = _GEN_15344 | valid_0_77; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2396 = _GEN_15345 | valid_0_78; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2397 = _GEN_15346 | valid_0_79; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2398 = _GEN_15347 | valid_0_80; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2399 = _GEN_15348 | valid_0_81; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2400 = _GEN_15349 | valid_0_82; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2401 = _GEN_15350 | valid_0_83; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2402 = _GEN_15351 | valid_0_84; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2403 = _GEN_15352 | valid_0_85; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2404 = _GEN_15353 | valid_0_86; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2405 = _GEN_15354 | valid_0_87; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2406 = _GEN_15355 | valid_0_88; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2407 = _GEN_15356 | valid_0_89; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2408 = _GEN_15357 | valid_0_90; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2409 = _GEN_15358 | valid_0_91; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2410 = _GEN_15359 | valid_0_92; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2411 = _GEN_15360 | valid_0_93; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2412 = _GEN_15361 | valid_0_94; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2413 = _GEN_15362 | valid_0_95; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2414 = _GEN_15363 | valid_0_96; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2415 = _GEN_15364 | valid_0_97; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2416 = _GEN_15365 | valid_0_98; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2417 = _GEN_15366 | valid_0_99; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2418 = _GEN_15367 | valid_0_100; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2419 = _GEN_15368 | valid_0_101; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2420 = _GEN_15369 | valid_0_102; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2421 = _GEN_15370 | valid_0_103; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2422 = _GEN_15371 | valid_0_104; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2423 = _GEN_15372 | valid_0_105; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2424 = _GEN_15373 | valid_0_106; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2425 = _GEN_15374 | valid_0_107; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2426 = _GEN_15375 | valid_0_108; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2427 = _GEN_15376 | valid_0_109; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2428 = _GEN_15377 | valid_0_110; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2429 = _GEN_15378 | valid_0_111; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2430 = _GEN_15379 | valid_0_112; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2431 = _GEN_15380 | valid_0_113; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2432 = _GEN_15381 | valid_0_114; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2433 = _GEN_15382 | valid_0_115; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2434 = _GEN_15383 | valid_0_116; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2435 = _GEN_15384 | valid_0_117; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2436 = _GEN_15385 | valid_0_118; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2437 = _GEN_15386 | valid_0_119; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2438 = _GEN_15387 | valid_0_120; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2439 = _GEN_15388 | valid_0_121; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2440 = _GEN_15389 | valid_0_122; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2441 = _GEN_15390 | valid_0_123; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2442 = _GEN_15391 | valid_0_124; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2443 = _GEN_15392 | valid_0_125; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2444 = _GEN_15393 | valid_0_126; // @[d_cache.scala 123:{32,32} 22:26]
  wire  _GEN_2445 = _GEN_15394 | valid_0_127; // @[d_cache.scala 123:{32,32} 22:26]
  wire [63:0] _GEN_2446 = 7'h0 == index ? receive_data : ram_1_0; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2447 = 7'h1 == index ? receive_data : ram_1_1; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2448 = 7'h2 == index ? receive_data : ram_1_2; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2449 = 7'h3 == index ? receive_data : ram_1_3; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2450 = 7'h4 == index ? receive_data : ram_1_4; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2451 = 7'h5 == index ? receive_data : ram_1_5; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2452 = 7'h6 == index ? receive_data : ram_1_6; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2453 = 7'h7 == index ? receive_data : ram_1_7; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2454 = 7'h8 == index ? receive_data : ram_1_8; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2455 = 7'h9 == index ? receive_data : ram_1_9; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2456 = 7'ha == index ? receive_data : ram_1_10; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2457 = 7'hb == index ? receive_data : ram_1_11; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2458 = 7'hc == index ? receive_data : ram_1_12; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2459 = 7'hd == index ? receive_data : ram_1_13; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2460 = 7'he == index ? receive_data : ram_1_14; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2461 = 7'hf == index ? receive_data : ram_1_15; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2462 = 7'h10 == index ? receive_data : ram_1_16; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2463 = 7'h11 == index ? receive_data : ram_1_17; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2464 = 7'h12 == index ? receive_data : ram_1_18; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2465 = 7'h13 == index ? receive_data : ram_1_19; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2466 = 7'h14 == index ? receive_data : ram_1_20; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2467 = 7'h15 == index ? receive_data : ram_1_21; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2468 = 7'h16 == index ? receive_data : ram_1_22; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2469 = 7'h17 == index ? receive_data : ram_1_23; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2470 = 7'h18 == index ? receive_data : ram_1_24; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2471 = 7'h19 == index ? receive_data : ram_1_25; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2472 = 7'h1a == index ? receive_data : ram_1_26; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2473 = 7'h1b == index ? receive_data : ram_1_27; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2474 = 7'h1c == index ? receive_data : ram_1_28; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2475 = 7'h1d == index ? receive_data : ram_1_29; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2476 = 7'h1e == index ? receive_data : ram_1_30; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2477 = 7'h1f == index ? receive_data : ram_1_31; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2478 = 7'h20 == index ? receive_data : ram_1_32; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2479 = 7'h21 == index ? receive_data : ram_1_33; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2480 = 7'h22 == index ? receive_data : ram_1_34; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2481 = 7'h23 == index ? receive_data : ram_1_35; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2482 = 7'h24 == index ? receive_data : ram_1_36; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2483 = 7'h25 == index ? receive_data : ram_1_37; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2484 = 7'h26 == index ? receive_data : ram_1_38; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2485 = 7'h27 == index ? receive_data : ram_1_39; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2486 = 7'h28 == index ? receive_data : ram_1_40; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2487 = 7'h29 == index ? receive_data : ram_1_41; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2488 = 7'h2a == index ? receive_data : ram_1_42; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2489 = 7'h2b == index ? receive_data : ram_1_43; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2490 = 7'h2c == index ? receive_data : ram_1_44; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2491 = 7'h2d == index ? receive_data : ram_1_45; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2492 = 7'h2e == index ? receive_data : ram_1_46; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2493 = 7'h2f == index ? receive_data : ram_1_47; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2494 = 7'h30 == index ? receive_data : ram_1_48; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2495 = 7'h31 == index ? receive_data : ram_1_49; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2496 = 7'h32 == index ? receive_data : ram_1_50; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2497 = 7'h33 == index ? receive_data : ram_1_51; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2498 = 7'h34 == index ? receive_data : ram_1_52; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2499 = 7'h35 == index ? receive_data : ram_1_53; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2500 = 7'h36 == index ? receive_data : ram_1_54; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2501 = 7'h37 == index ? receive_data : ram_1_55; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2502 = 7'h38 == index ? receive_data : ram_1_56; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2503 = 7'h39 == index ? receive_data : ram_1_57; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2504 = 7'h3a == index ? receive_data : ram_1_58; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2505 = 7'h3b == index ? receive_data : ram_1_59; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2506 = 7'h3c == index ? receive_data : ram_1_60; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2507 = 7'h3d == index ? receive_data : ram_1_61; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2508 = 7'h3e == index ? receive_data : ram_1_62; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2509 = 7'h3f == index ? receive_data : ram_1_63; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2510 = 7'h40 == index ? receive_data : ram_1_64; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2511 = 7'h41 == index ? receive_data : ram_1_65; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2512 = 7'h42 == index ? receive_data : ram_1_66; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2513 = 7'h43 == index ? receive_data : ram_1_67; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2514 = 7'h44 == index ? receive_data : ram_1_68; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2515 = 7'h45 == index ? receive_data : ram_1_69; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2516 = 7'h46 == index ? receive_data : ram_1_70; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2517 = 7'h47 == index ? receive_data : ram_1_71; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2518 = 7'h48 == index ? receive_data : ram_1_72; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2519 = 7'h49 == index ? receive_data : ram_1_73; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2520 = 7'h4a == index ? receive_data : ram_1_74; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2521 = 7'h4b == index ? receive_data : ram_1_75; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2522 = 7'h4c == index ? receive_data : ram_1_76; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2523 = 7'h4d == index ? receive_data : ram_1_77; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2524 = 7'h4e == index ? receive_data : ram_1_78; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2525 = 7'h4f == index ? receive_data : ram_1_79; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2526 = 7'h50 == index ? receive_data : ram_1_80; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2527 = 7'h51 == index ? receive_data : ram_1_81; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2528 = 7'h52 == index ? receive_data : ram_1_82; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2529 = 7'h53 == index ? receive_data : ram_1_83; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2530 = 7'h54 == index ? receive_data : ram_1_84; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2531 = 7'h55 == index ? receive_data : ram_1_85; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2532 = 7'h56 == index ? receive_data : ram_1_86; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2533 = 7'h57 == index ? receive_data : ram_1_87; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2534 = 7'h58 == index ? receive_data : ram_1_88; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2535 = 7'h59 == index ? receive_data : ram_1_89; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2536 = 7'h5a == index ? receive_data : ram_1_90; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2537 = 7'h5b == index ? receive_data : ram_1_91; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2538 = 7'h5c == index ? receive_data : ram_1_92; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2539 = 7'h5d == index ? receive_data : ram_1_93; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2540 = 7'h5e == index ? receive_data : ram_1_94; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2541 = 7'h5f == index ? receive_data : ram_1_95; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2542 = 7'h60 == index ? receive_data : ram_1_96; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2543 = 7'h61 == index ? receive_data : ram_1_97; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2544 = 7'h62 == index ? receive_data : ram_1_98; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2545 = 7'h63 == index ? receive_data : ram_1_99; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2546 = 7'h64 == index ? receive_data : ram_1_100; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2547 = 7'h65 == index ? receive_data : ram_1_101; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2548 = 7'h66 == index ? receive_data : ram_1_102; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2549 = 7'h67 == index ? receive_data : ram_1_103; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2550 = 7'h68 == index ? receive_data : ram_1_104; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2551 = 7'h69 == index ? receive_data : ram_1_105; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2552 = 7'h6a == index ? receive_data : ram_1_106; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2553 = 7'h6b == index ? receive_data : ram_1_107; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2554 = 7'h6c == index ? receive_data : ram_1_108; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2555 = 7'h6d == index ? receive_data : ram_1_109; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2556 = 7'h6e == index ? receive_data : ram_1_110; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2557 = 7'h6f == index ? receive_data : ram_1_111; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2558 = 7'h70 == index ? receive_data : ram_1_112; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2559 = 7'h71 == index ? receive_data : ram_1_113; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2560 = 7'h72 == index ? receive_data : ram_1_114; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2561 = 7'h73 == index ? receive_data : ram_1_115; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2562 = 7'h74 == index ? receive_data : ram_1_116; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2563 = 7'h75 == index ? receive_data : ram_1_117; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2564 = 7'h76 == index ? receive_data : ram_1_118; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2565 = 7'h77 == index ? receive_data : ram_1_119; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2566 = 7'h78 == index ? receive_data : ram_1_120; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2567 = 7'h79 == index ? receive_data : ram_1_121; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2568 = 7'h7a == index ? receive_data : ram_1_122; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2569 = 7'h7b == index ? receive_data : ram_1_123; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2570 = 7'h7c == index ? receive_data : ram_1_124; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2571 = 7'h7d == index ? receive_data : ram_1_125; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2572 = 7'h7e == index ? receive_data : ram_1_126; // @[d_cache.scala 127:{30,30} 19:24]
  wire [63:0] _GEN_2573 = 7'h7f == index ? receive_data : ram_1_127; // @[d_cache.scala 127:{30,30} 19:24]
  wire [31:0] _GEN_2574 = 7'h0 == index ? _GEN_15265 : tag_1_0; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2575 = 7'h1 == index ? _GEN_15265 : tag_1_1; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2576 = 7'h2 == index ? _GEN_15265 : tag_1_2; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2577 = 7'h3 == index ? _GEN_15265 : tag_1_3; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2578 = 7'h4 == index ? _GEN_15265 : tag_1_4; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2579 = 7'h5 == index ? _GEN_15265 : tag_1_5; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2580 = 7'h6 == index ? _GEN_15265 : tag_1_6; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2581 = 7'h7 == index ? _GEN_15265 : tag_1_7; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2582 = 7'h8 == index ? _GEN_15265 : tag_1_8; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2583 = 7'h9 == index ? _GEN_15265 : tag_1_9; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2584 = 7'ha == index ? _GEN_15265 : tag_1_10; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2585 = 7'hb == index ? _GEN_15265 : tag_1_11; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2586 = 7'hc == index ? _GEN_15265 : tag_1_12; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2587 = 7'hd == index ? _GEN_15265 : tag_1_13; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2588 = 7'he == index ? _GEN_15265 : tag_1_14; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2589 = 7'hf == index ? _GEN_15265 : tag_1_15; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2590 = 7'h10 == index ? _GEN_15265 : tag_1_16; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2591 = 7'h11 == index ? _GEN_15265 : tag_1_17; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2592 = 7'h12 == index ? _GEN_15265 : tag_1_18; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2593 = 7'h13 == index ? _GEN_15265 : tag_1_19; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2594 = 7'h14 == index ? _GEN_15265 : tag_1_20; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2595 = 7'h15 == index ? _GEN_15265 : tag_1_21; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2596 = 7'h16 == index ? _GEN_15265 : tag_1_22; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2597 = 7'h17 == index ? _GEN_15265 : tag_1_23; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2598 = 7'h18 == index ? _GEN_15265 : tag_1_24; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2599 = 7'h19 == index ? _GEN_15265 : tag_1_25; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2600 = 7'h1a == index ? _GEN_15265 : tag_1_26; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2601 = 7'h1b == index ? _GEN_15265 : tag_1_27; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2602 = 7'h1c == index ? _GEN_15265 : tag_1_28; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2603 = 7'h1d == index ? _GEN_15265 : tag_1_29; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2604 = 7'h1e == index ? _GEN_15265 : tag_1_30; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2605 = 7'h1f == index ? _GEN_15265 : tag_1_31; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2606 = 7'h20 == index ? _GEN_15265 : tag_1_32; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2607 = 7'h21 == index ? _GEN_15265 : tag_1_33; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2608 = 7'h22 == index ? _GEN_15265 : tag_1_34; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2609 = 7'h23 == index ? _GEN_15265 : tag_1_35; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2610 = 7'h24 == index ? _GEN_15265 : tag_1_36; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2611 = 7'h25 == index ? _GEN_15265 : tag_1_37; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2612 = 7'h26 == index ? _GEN_15265 : tag_1_38; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2613 = 7'h27 == index ? _GEN_15265 : tag_1_39; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2614 = 7'h28 == index ? _GEN_15265 : tag_1_40; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2615 = 7'h29 == index ? _GEN_15265 : tag_1_41; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2616 = 7'h2a == index ? _GEN_15265 : tag_1_42; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2617 = 7'h2b == index ? _GEN_15265 : tag_1_43; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2618 = 7'h2c == index ? _GEN_15265 : tag_1_44; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2619 = 7'h2d == index ? _GEN_15265 : tag_1_45; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2620 = 7'h2e == index ? _GEN_15265 : tag_1_46; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2621 = 7'h2f == index ? _GEN_15265 : tag_1_47; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2622 = 7'h30 == index ? _GEN_15265 : tag_1_48; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2623 = 7'h31 == index ? _GEN_15265 : tag_1_49; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2624 = 7'h32 == index ? _GEN_15265 : tag_1_50; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2625 = 7'h33 == index ? _GEN_15265 : tag_1_51; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2626 = 7'h34 == index ? _GEN_15265 : tag_1_52; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2627 = 7'h35 == index ? _GEN_15265 : tag_1_53; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2628 = 7'h36 == index ? _GEN_15265 : tag_1_54; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2629 = 7'h37 == index ? _GEN_15265 : tag_1_55; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2630 = 7'h38 == index ? _GEN_15265 : tag_1_56; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2631 = 7'h39 == index ? _GEN_15265 : tag_1_57; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2632 = 7'h3a == index ? _GEN_15265 : tag_1_58; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2633 = 7'h3b == index ? _GEN_15265 : tag_1_59; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2634 = 7'h3c == index ? _GEN_15265 : tag_1_60; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2635 = 7'h3d == index ? _GEN_15265 : tag_1_61; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2636 = 7'h3e == index ? _GEN_15265 : tag_1_62; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2637 = 7'h3f == index ? _GEN_15265 : tag_1_63; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2638 = 7'h40 == index ? _GEN_15265 : tag_1_64; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2639 = 7'h41 == index ? _GEN_15265 : tag_1_65; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2640 = 7'h42 == index ? _GEN_15265 : tag_1_66; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2641 = 7'h43 == index ? _GEN_15265 : tag_1_67; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2642 = 7'h44 == index ? _GEN_15265 : tag_1_68; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2643 = 7'h45 == index ? _GEN_15265 : tag_1_69; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2644 = 7'h46 == index ? _GEN_15265 : tag_1_70; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2645 = 7'h47 == index ? _GEN_15265 : tag_1_71; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2646 = 7'h48 == index ? _GEN_15265 : tag_1_72; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2647 = 7'h49 == index ? _GEN_15265 : tag_1_73; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2648 = 7'h4a == index ? _GEN_15265 : tag_1_74; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2649 = 7'h4b == index ? _GEN_15265 : tag_1_75; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2650 = 7'h4c == index ? _GEN_15265 : tag_1_76; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2651 = 7'h4d == index ? _GEN_15265 : tag_1_77; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2652 = 7'h4e == index ? _GEN_15265 : tag_1_78; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2653 = 7'h4f == index ? _GEN_15265 : tag_1_79; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2654 = 7'h50 == index ? _GEN_15265 : tag_1_80; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2655 = 7'h51 == index ? _GEN_15265 : tag_1_81; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2656 = 7'h52 == index ? _GEN_15265 : tag_1_82; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2657 = 7'h53 == index ? _GEN_15265 : tag_1_83; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2658 = 7'h54 == index ? _GEN_15265 : tag_1_84; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2659 = 7'h55 == index ? _GEN_15265 : tag_1_85; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2660 = 7'h56 == index ? _GEN_15265 : tag_1_86; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2661 = 7'h57 == index ? _GEN_15265 : tag_1_87; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2662 = 7'h58 == index ? _GEN_15265 : tag_1_88; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2663 = 7'h59 == index ? _GEN_15265 : tag_1_89; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2664 = 7'h5a == index ? _GEN_15265 : tag_1_90; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2665 = 7'h5b == index ? _GEN_15265 : tag_1_91; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2666 = 7'h5c == index ? _GEN_15265 : tag_1_92; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2667 = 7'h5d == index ? _GEN_15265 : tag_1_93; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2668 = 7'h5e == index ? _GEN_15265 : tag_1_94; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2669 = 7'h5f == index ? _GEN_15265 : tag_1_95; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2670 = 7'h60 == index ? _GEN_15265 : tag_1_96; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2671 = 7'h61 == index ? _GEN_15265 : tag_1_97; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2672 = 7'h62 == index ? _GEN_15265 : tag_1_98; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2673 = 7'h63 == index ? _GEN_15265 : tag_1_99; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2674 = 7'h64 == index ? _GEN_15265 : tag_1_100; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2675 = 7'h65 == index ? _GEN_15265 : tag_1_101; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2676 = 7'h66 == index ? _GEN_15265 : tag_1_102; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2677 = 7'h67 == index ? _GEN_15265 : tag_1_103; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2678 = 7'h68 == index ? _GEN_15265 : tag_1_104; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2679 = 7'h69 == index ? _GEN_15265 : tag_1_105; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2680 = 7'h6a == index ? _GEN_15265 : tag_1_106; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2681 = 7'h6b == index ? _GEN_15265 : tag_1_107; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2682 = 7'h6c == index ? _GEN_15265 : tag_1_108; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2683 = 7'h6d == index ? _GEN_15265 : tag_1_109; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2684 = 7'h6e == index ? _GEN_15265 : tag_1_110; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2685 = 7'h6f == index ? _GEN_15265 : tag_1_111; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2686 = 7'h70 == index ? _GEN_15265 : tag_1_112; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2687 = 7'h71 == index ? _GEN_15265 : tag_1_113; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2688 = 7'h72 == index ? _GEN_15265 : tag_1_114; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2689 = 7'h73 == index ? _GEN_15265 : tag_1_115; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2690 = 7'h74 == index ? _GEN_15265 : tag_1_116; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2691 = 7'h75 == index ? _GEN_15265 : tag_1_117; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2692 = 7'h76 == index ? _GEN_15265 : tag_1_118; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2693 = 7'h77 == index ? _GEN_15265 : tag_1_119; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2694 = 7'h78 == index ? _GEN_15265 : tag_1_120; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2695 = 7'h79 == index ? _GEN_15265 : tag_1_121; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2696 = 7'h7a == index ? _GEN_15265 : tag_1_122; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2697 = 7'h7b == index ? _GEN_15265 : tag_1_123; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2698 = 7'h7c == index ? _GEN_15265 : tag_1_124; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2699 = 7'h7d == index ? _GEN_15265 : tag_1_125; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2700 = 7'h7e == index ? _GEN_15265 : tag_1_126; // @[d_cache.scala 128:{30,30} 21:24]
  wire [31:0] _GEN_2701 = 7'h7f == index ? _GEN_15265 : tag_1_127; // @[d_cache.scala 128:{30,30} 21:24]
  wire  _GEN_2702 = _GEN_15267 | valid_1_0; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2703 = _GEN_15268 | valid_1_1; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2704 = _GEN_15269 | valid_1_2; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2705 = _GEN_15270 | valid_1_3; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2706 = _GEN_15271 | valid_1_4; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2707 = _GEN_15272 | valid_1_5; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2708 = _GEN_15273 | valid_1_6; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2709 = _GEN_15274 | valid_1_7; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2710 = _GEN_15275 | valid_1_8; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2711 = _GEN_15276 | valid_1_9; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2712 = _GEN_15277 | valid_1_10; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2713 = _GEN_15278 | valid_1_11; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2714 = _GEN_15279 | valid_1_12; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2715 = _GEN_15280 | valid_1_13; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2716 = _GEN_15281 | valid_1_14; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2717 = _GEN_15282 | valid_1_15; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2718 = _GEN_15283 | valid_1_16; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2719 = _GEN_15284 | valid_1_17; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2720 = _GEN_15285 | valid_1_18; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2721 = _GEN_15286 | valid_1_19; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2722 = _GEN_15287 | valid_1_20; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2723 = _GEN_15288 | valid_1_21; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2724 = _GEN_15289 | valid_1_22; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2725 = _GEN_15290 | valid_1_23; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2726 = _GEN_15291 | valid_1_24; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2727 = _GEN_15292 | valid_1_25; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2728 = _GEN_15293 | valid_1_26; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2729 = _GEN_15294 | valid_1_27; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2730 = _GEN_15295 | valid_1_28; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2731 = _GEN_15296 | valid_1_29; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2732 = _GEN_15297 | valid_1_30; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2733 = _GEN_15298 | valid_1_31; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2734 = _GEN_15299 | valid_1_32; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2735 = _GEN_15300 | valid_1_33; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2736 = _GEN_15301 | valid_1_34; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2737 = _GEN_15302 | valid_1_35; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2738 = _GEN_15303 | valid_1_36; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2739 = _GEN_15304 | valid_1_37; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2740 = _GEN_15305 | valid_1_38; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2741 = _GEN_15306 | valid_1_39; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2742 = _GEN_15307 | valid_1_40; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2743 = _GEN_15308 | valid_1_41; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2744 = _GEN_15309 | valid_1_42; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2745 = _GEN_15310 | valid_1_43; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2746 = _GEN_15311 | valid_1_44; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2747 = _GEN_15312 | valid_1_45; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2748 = _GEN_15313 | valid_1_46; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2749 = _GEN_15314 | valid_1_47; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2750 = _GEN_15315 | valid_1_48; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2751 = _GEN_15316 | valid_1_49; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2752 = _GEN_15317 | valid_1_50; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2753 = _GEN_15318 | valid_1_51; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2754 = _GEN_15319 | valid_1_52; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2755 = _GEN_15320 | valid_1_53; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2756 = _GEN_15321 | valid_1_54; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2757 = _GEN_15322 | valid_1_55; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2758 = _GEN_15323 | valid_1_56; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2759 = _GEN_15324 | valid_1_57; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2760 = _GEN_15325 | valid_1_58; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2761 = _GEN_15326 | valid_1_59; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2762 = _GEN_15327 | valid_1_60; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2763 = _GEN_15328 | valid_1_61; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2764 = _GEN_15329 | valid_1_62; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2765 = _GEN_15330 | valid_1_63; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2766 = _GEN_15331 | valid_1_64; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2767 = _GEN_15332 | valid_1_65; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2768 = _GEN_15333 | valid_1_66; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2769 = _GEN_15334 | valid_1_67; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2770 = _GEN_15335 | valid_1_68; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2771 = _GEN_15336 | valid_1_69; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2772 = _GEN_15337 | valid_1_70; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2773 = _GEN_15338 | valid_1_71; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2774 = _GEN_15339 | valid_1_72; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2775 = _GEN_15340 | valid_1_73; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2776 = _GEN_15341 | valid_1_74; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2777 = _GEN_15342 | valid_1_75; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2778 = _GEN_15343 | valid_1_76; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2779 = _GEN_15344 | valid_1_77; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2780 = _GEN_15345 | valid_1_78; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2781 = _GEN_15346 | valid_1_79; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2782 = _GEN_15347 | valid_1_80; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2783 = _GEN_15348 | valid_1_81; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2784 = _GEN_15349 | valid_1_82; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2785 = _GEN_15350 | valid_1_83; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2786 = _GEN_15351 | valid_1_84; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2787 = _GEN_15352 | valid_1_85; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2788 = _GEN_15353 | valid_1_86; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2789 = _GEN_15354 | valid_1_87; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2790 = _GEN_15355 | valid_1_88; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2791 = _GEN_15356 | valid_1_89; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2792 = _GEN_15357 | valid_1_90; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2793 = _GEN_15358 | valid_1_91; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2794 = _GEN_15359 | valid_1_92; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2795 = _GEN_15360 | valid_1_93; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2796 = _GEN_15361 | valid_1_94; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2797 = _GEN_15362 | valid_1_95; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2798 = _GEN_15363 | valid_1_96; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2799 = _GEN_15364 | valid_1_97; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2800 = _GEN_15365 | valid_1_98; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2801 = _GEN_15366 | valid_1_99; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2802 = _GEN_15367 | valid_1_100; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2803 = _GEN_15368 | valid_1_101; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2804 = _GEN_15369 | valid_1_102; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2805 = _GEN_15370 | valid_1_103; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2806 = _GEN_15371 | valid_1_104; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2807 = _GEN_15372 | valid_1_105; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2808 = _GEN_15373 | valid_1_106; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2809 = _GEN_15374 | valid_1_107; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2810 = _GEN_15375 | valid_1_108; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2811 = _GEN_15376 | valid_1_109; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2812 = _GEN_15377 | valid_1_110; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2813 = _GEN_15378 | valid_1_111; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2814 = _GEN_15379 | valid_1_112; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2815 = _GEN_15380 | valid_1_113; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2816 = _GEN_15381 | valid_1_114; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2817 = _GEN_15382 | valid_1_115; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2818 = _GEN_15383 | valid_1_116; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2819 = _GEN_15384 | valid_1_117; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2820 = _GEN_15385 | valid_1_118; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2821 = _GEN_15386 | valid_1_119; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2822 = _GEN_15387 | valid_1_120; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2823 = _GEN_15388 | valid_1_121; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2824 = _GEN_15389 | valid_1_122; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2825 = _GEN_15390 | valid_1_123; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2826 = _GEN_15391 | valid_1_124; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2827 = _GEN_15392 | valid_1_125; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2828 = _GEN_15393 | valid_1_126; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _GEN_2829 = _GEN_15394 | valid_1_127; // @[d_cache.scala 129:{32,32} 23:26]
  wire  _T_28 = ~quene; // @[d_cache.scala 132:27]
  wire [63:0] _GEN_2831 = 7'h1 == index ? ram_0_1 : ram_0_0; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2832 = 7'h2 == index ? ram_0_2 : _GEN_2831; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2833 = 7'h3 == index ? ram_0_3 : _GEN_2832; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2834 = 7'h4 == index ? ram_0_4 : _GEN_2833; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2835 = 7'h5 == index ? ram_0_5 : _GEN_2834; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2836 = 7'h6 == index ? ram_0_6 : _GEN_2835; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2837 = 7'h7 == index ? ram_0_7 : _GEN_2836; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2838 = 7'h8 == index ? ram_0_8 : _GEN_2837; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2839 = 7'h9 == index ? ram_0_9 : _GEN_2838; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2840 = 7'ha == index ? ram_0_10 : _GEN_2839; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2841 = 7'hb == index ? ram_0_11 : _GEN_2840; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2842 = 7'hc == index ? ram_0_12 : _GEN_2841; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2843 = 7'hd == index ? ram_0_13 : _GEN_2842; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2844 = 7'he == index ? ram_0_14 : _GEN_2843; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2845 = 7'hf == index ? ram_0_15 : _GEN_2844; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2846 = 7'h10 == index ? ram_0_16 : _GEN_2845; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2847 = 7'h11 == index ? ram_0_17 : _GEN_2846; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2848 = 7'h12 == index ? ram_0_18 : _GEN_2847; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2849 = 7'h13 == index ? ram_0_19 : _GEN_2848; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2850 = 7'h14 == index ? ram_0_20 : _GEN_2849; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2851 = 7'h15 == index ? ram_0_21 : _GEN_2850; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2852 = 7'h16 == index ? ram_0_22 : _GEN_2851; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2853 = 7'h17 == index ? ram_0_23 : _GEN_2852; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2854 = 7'h18 == index ? ram_0_24 : _GEN_2853; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2855 = 7'h19 == index ? ram_0_25 : _GEN_2854; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2856 = 7'h1a == index ? ram_0_26 : _GEN_2855; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2857 = 7'h1b == index ? ram_0_27 : _GEN_2856; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2858 = 7'h1c == index ? ram_0_28 : _GEN_2857; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2859 = 7'h1d == index ? ram_0_29 : _GEN_2858; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2860 = 7'h1e == index ? ram_0_30 : _GEN_2859; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2861 = 7'h1f == index ? ram_0_31 : _GEN_2860; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2862 = 7'h20 == index ? ram_0_32 : _GEN_2861; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2863 = 7'h21 == index ? ram_0_33 : _GEN_2862; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2864 = 7'h22 == index ? ram_0_34 : _GEN_2863; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2865 = 7'h23 == index ? ram_0_35 : _GEN_2864; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2866 = 7'h24 == index ? ram_0_36 : _GEN_2865; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2867 = 7'h25 == index ? ram_0_37 : _GEN_2866; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2868 = 7'h26 == index ? ram_0_38 : _GEN_2867; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2869 = 7'h27 == index ? ram_0_39 : _GEN_2868; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2870 = 7'h28 == index ? ram_0_40 : _GEN_2869; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2871 = 7'h29 == index ? ram_0_41 : _GEN_2870; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2872 = 7'h2a == index ? ram_0_42 : _GEN_2871; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2873 = 7'h2b == index ? ram_0_43 : _GEN_2872; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2874 = 7'h2c == index ? ram_0_44 : _GEN_2873; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2875 = 7'h2d == index ? ram_0_45 : _GEN_2874; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2876 = 7'h2e == index ? ram_0_46 : _GEN_2875; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2877 = 7'h2f == index ? ram_0_47 : _GEN_2876; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2878 = 7'h30 == index ? ram_0_48 : _GEN_2877; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2879 = 7'h31 == index ? ram_0_49 : _GEN_2878; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2880 = 7'h32 == index ? ram_0_50 : _GEN_2879; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2881 = 7'h33 == index ? ram_0_51 : _GEN_2880; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2882 = 7'h34 == index ? ram_0_52 : _GEN_2881; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2883 = 7'h35 == index ? ram_0_53 : _GEN_2882; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2884 = 7'h36 == index ? ram_0_54 : _GEN_2883; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2885 = 7'h37 == index ? ram_0_55 : _GEN_2884; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2886 = 7'h38 == index ? ram_0_56 : _GEN_2885; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2887 = 7'h39 == index ? ram_0_57 : _GEN_2886; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2888 = 7'h3a == index ? ram_0_58 : _GEN_2887; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2889 = 7'h3b == index ? ram_0_59 : _GEN_2888; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2890 = 7'h3c == index ? ram_0_60 : _GEN_2889; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2891 = 7'h3d == index ? ram_0_61 : _GEN_2890; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2892 = 7'h3e == index ? ram_0_62 : _GEN_2891; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2893 = 7'h3f == index ? ram_0_63 : _GEN_2892; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2894 = 7'h40 == index ? ram_0_64 : _GEN_2893; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2895 = 7'h41 == index ? ram_0_65 : _GEN_2894; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2896 = 7'h42 == index ? ram_0_66 : _GEN_2895; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2897 = 7'h43 == index ? ram_0_67 : _GEN_2896; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2898 = 7'h44 == index ? ram_0_68 : _GEN_2897; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2899 = 7'h45 == index ? ram_0_69 : _GEN_2898; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2900 = 7'h46 == index ? ram_0_70 : _GEN_2899; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2901 = 7'h47 == index ? ram_0_71 : _GEN_2900; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2902 = 7'h48 == index ? ram_0_72 : _GEN_2901; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2903 = 7'h49 == index ? ram_0_73 : _GEN_2902; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2904 = 7'h4a == index ? ram_0_74 : _GEN_2903; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2905 = 7'h4b == index ? ram_0_75 : _GEN_2904; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2906 = 7'h4c == index ? ram_0_76 : _GEN_2905; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2907 = 7'h4d == index ? ram_0_77 : _GEN_2906; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2908 = 7'h4e == index ? ram_0_78 : _GEN_2907; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2909 = 7'h4f == index ? ram_0_79 : _GEN_2908; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2910 = 7'h50 == index ? ram_0_80 : _GEN_2909; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2911 = 7'h51 == index ? ram_0_81 : _GEN_2910; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2912 = 7'h52 == index ? ram_0_82 : _GEN_2911; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2913 = 7'h53 == index ? ram_0_83 : _GEN_2912; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2914 = 7'h54 == index ? ram_0_84 : _GEN_2913; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2915 = 7'h55 == index ? ram_0_85 : _GEN_2914; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2916 = 7'h56 == index ? ram_0_86 : _GEN_2915; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2917 = 7'h57 == index ? ram_0_87 : _GEN_2916; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2918 = 7'h58 == index ? ram_0_88 : _GEN_2917; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2919 = 7'h59 == index ? ram_0_89 : _GEN_2918; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2920 = 7'h5a == index ? ram_0_90 : _GEN_2919; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2921 = 7'h5b == index ? ram_0_91 : _GEN_2920; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2922 = 7'h5c == index ? ram_0_92 : _GEN_2921; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2923 = 7'h5d == index ? ram_0_93 : _GEN_2922; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2924 = 7'h5e == index ? ram_0_94 : _GEN_2923; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2925 = 7'h5f == index ? ram_0_95 : _GEN_2924; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2926 = 7'h60 == index ? ram_0_96 : _GEN_2925; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2927 = 7'h61 == index ? ram_0_97 : _GEN_2926; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2928 = 7'h62 == index ? ram_0_98 : _GEN_2927; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2929 = 7'h63 == index ? ram_0_99 : _GEN_2928; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2930 = 7'h64 == index ? ram_0_100 : _GEN_2929; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2931 = 7'h65 == index ? ram_0_101 : _GEN_2930; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2932 = 7'h66 == index ? ram_0_102 : _GEN_2931; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2933 = 7'h67 == index ? ram_0_103 : _GEN_2932; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2934 = 7'h68 == index ? ram_0_104 : _GEN_2933; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2935 = 7'h69 == index ? ram_0_105 : _GEN_2934; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2936 = 7'h6a == index ? ram_0_106 : _GEN_2935; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2937 = 7'h6b == index ? ram_0_107 : _GEN_2936; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2938 = 7'h6c == index ? ram_0_108 : _GEN_2937; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2939 = 7'h6d == index ? ram_0_109 : _GEN_2938; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2940 = 7'h6e == index ? ram_0_110 : _GEN_2939; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2941 = 7'h6f == index ? ram_0_111 : _GEN_2940; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2942 = 7'h70 == index ? ram_0_112 : _GEN_2941; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2943 = 7'h71 == index ? ram_0_113 : _GEN_2942; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2944 = 7'h72 == index ? ram_0_114 : _GEN_2943; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2945 = 7'h73 == index ? ram_0_115 : _GEN_2944; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2946 = 7'h74 == index ? ram_0_116 : _GEN_2945; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2947 = 7'h75 == index ? ram_0_117 : _GEN_2946; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2948 = 7'h76 == index ? ram_0_118 : _GEN_2947; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2949 = 7'h77 == index ? ram_0_119 : _GEN_2948; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2950 = 7'h78 == index ? ram_0_120 : _GEN_2949; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2951 = 7'h79 == index ? ram_0_121 : _GEN_2950; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2952 = 7'h7a == index ? ram_0_122 : _GEN_2951; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2953 = 7'h7b == index ? ram_0_123 : _GEN_2952; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2954 = 7'h7c == index ? ram_0_124 : _GEN_2953; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2955 = 7'h7d == index ? ram_0_125 : _GEN_2954; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2956 = 7'h7e == index ? ram_0_126 : _GEN_2955; // @[d_cache.scala 135:{41,41}]
  wire [63:0] _GEN_2957 = 7'h7f == index ? ram_0_127 : _GEN_2956; // @[d_cache.scala 135:{41,41}]
  wire [38:0] _write_back_addr_T = {_GEN_127, 7'h0}; // @[d_cache.scala 136:57]
  wire [38:0] _GEN_15779 = {{32'd0}, index}; // @[d_cache.scala 136:62]
  wire [38:0] _write_back_addr_T_1 = _write_back_addr_T | _GEN_15779; // @[d_cache.scala 136:62]
  wire  _GEN_3214 = 7'h0 == index ? 1'h0 : dirty_0_0; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3215 = 7'h1 == index ? 1'h0 : dirty_0_1; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3216 = 7'h2 == index ? 1'h0 : dirty_0_2; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3217 = 7'h3 == index ? 1'h0 : dirty_0_3; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3218 = 7'h4 == index ? 1'h0 : dirty_0_4; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3219 = 7'h5 == index ? 1'h0 : dirty_0_5; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3220 = 7'h6 == index ? 1'h0 : dirty_0_6; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3221 = 7'h7 == index ? 1'h0 : dirty_0_7; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3222 = 7'h8 == index ? 1'h0 : dirty_0_8; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3223 = 7'h9 == index ? 1'h0 : dirty_0_9; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3224 = 7'ha == index ? 1'h0 : dirty_0_10; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3225 = 7'hb == index ? 1'h0 : dirty_0_11; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3226 = 7'hc == index ? 1'h0 : dirty_0_12; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3227 = 7'hd == index ? 1'h0 : dirty_0_13; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3228 = 7'he == index ? 1'h0 : dirty_0_14; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3229 = 7'hf == index ? 1'h0 : dirty_0_15; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3230 = 7'h10 == index ? 1'h0 : dirty_0_16; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3231 = 7'h11 == index ? 1'h0 : dirty_0_17; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3232 = 7'h12 == index ? 1'h0 : dirty_0_18; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3233 = 7'h13 == index ? 1'h0 : dirty_0_19; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3234 = 7'h14 == index ? 1'h0 : dirty_0_20; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3235 = 7'h15 == index ? 1'h0 : dirty_0_21; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3236 = 7'h16 == index ? 1'h0 : dirty_0_22; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3237 = 7'h17 == index ? 1'h0 : dirty_0_23; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3238 = 7'h18 == index ? 1'h0 : dirty_0_24; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3239 = 7'h19 == index ? 1'h0 : dirty_0_25; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3240 = 7'h1a == index ? 1'h0 : dirty_0_26; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3241 = 7'h1b == index ? 1'h0 : dirty_0_27; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3242 = 7'h1c == index ? 1'h0 : dirty_0_28; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3243 = 7'h1d == index ? 1'h0 : dirty_0_29; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3244 = 7'h1e == index ? 1'h0 : dirty_0_30; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3245 = 7'h1f == index ? 1'h0 : dirty_0_31; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3246 = 7'h20 == index ? 1'h0 : dirty_0_32; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3247 = 7'h21 == index ? 1'h0 : dirty_0_33; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3248 = 7'h22 == index ? 1'h0 : dirty_0_34; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3249 = 7'h23 == index ? 1'h0 : dirty_0_35; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3250 = 7'h24 == index ? 1'h0 : dirty_0_36; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3251 = 7'h25 == index ? 1'h0 : dirty_0_37; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3252 = 7'h26 == index ? 1'h0 : dirty_0_38; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3253 = 7'h27 == index ? 1'h0 : dirty_0_39; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3254 = 7'h28 == index ? 1'h0 : dirty_0_40; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3255 = 7'h29 == index ? 1'h0 : dirty_0_41; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3256 = 7'h2a == index ? 1'h0 : dirty_0_42; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3257 = 7'h2b == index ? 1'h0 : dirty_0_43; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3258 = 7'h2c == index ? 1'h0 : dirty_0_44; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3259 = 7'h2d == index ? 1'h0 : dirty_0_45; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3260 = 7'h2e == index ? 1'h0 : dirty_0_46; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3261 = 7'h2f == index ? 1'h0 : dirty_0_47; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3262 = 7'h30 == index ? 1'h0 : dirty_0_48; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3263 = 7'h31 == index ? 1'h0 : dirty_0_49; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3264 = 7'h32 == index ? 1'h0 : dirty_0_50; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3265 = 7'h33 == index ? 1'h0 : dirty_0_51; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3266 = 7'h34 == index ? 1'h0 : dirty_0_52; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3267 = 7'h35 == index ? 1'h0 : dirty_0_53; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3268 = 7'h36 == index ? 1'h0 : dirty_0_54; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3269 = 7'h37 == index ? 1'h0 : dirty_0_55; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3270 = 7'h38 == index ? 1'h0 : dirty_0_56; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3271 = 7'h39 == index ? 1'h0 : dirty_0_57; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3272 = 7'h3a == index ? 1'h0 : dirty_0_58; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3273 = 7'h3b == index ? 1'h0 : dirty_0_59; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3274 = 7'h3c == index ? 1'h0 : dirty_0_60; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3275 = 7'h3d == index ? 1'h0 : dirty_0_61; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3276 = 7'h3e == index ? 1'h0 : dirty_0_62; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3277 = 7'h3f == index ? 1'h0 : dirty_0_63; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3278 = 7'h40 == index ? 1'h0 : dirty_0_64; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3279 = 7'h41 == index ? 1'h0 : dirty_0_65; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3280 = 7'h42 == index ? 1'h0 : dirty_0_66; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3281 = 7'h43 == index ? 1'h0 : dirty_0_67; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3282 = 7'h44 == index ? 1'h0 : dirty_0_68; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3283 = 7'h45 == index ? 1'h0 : dirty_0_69; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3284 = 7'h46 == index ? 1'h0 : dirty_0_70; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3285 = 7'h47 == index ? 1'h0 : dirty_0_71; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3286 = 7'h48 == index ? 1'h0 : dirty_0_72; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3287 = 7'h49 == index ? 1'h0 : dirty_0_73; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3288 = 7'h4a == index ? 1'h0 : dirty_0_74; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3289 = 7'h4b == index ? 1'h0 : dirty_0_75; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3290 = 7'h4c == index ? 1'h0 : dirty_0_76; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3291 = 7'h4d == index ? 1'h0 : dirty_0_77; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3292 = 7'h4e == index ? 1'h0 : dirty_0_78; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3293 = 7'h4f == index ? 1'h0 : dirty_0_79; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3294 = 7'h50 == index ? 1'h0 : dirty_0_80; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3295 = 7'h51 == index ? 1'h0 : dirty_0_81; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3296 = 7'h52 == index ? 1'h0 : dirty_0_82; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3297 = 7'h53 == index ? 1'h0 : dirty_0_83; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3298 = 7'h54 == index ? 1'h0 : dirty_0_84; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3299 = 7'h55 == index ? 1'h0 : dirty_0_85; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3300 = 7'h56 == index ? 1'h0 : dirty_0_86; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3301 = 7'h57 == index ? 1'h0 : dirty_0_87; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3302 = 7'h58 == index ? 1'h0 : dirty_0_88; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3303 = 7'h59 == index ? 1'h0 : dirty_0_89; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3304 = 7'h5a == index ? 1'h0 : dirty_0_90; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3305 = 7'h5b == index ? 1'h0 : dirty_0_91; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3306 = 7'h5c == index ? 1'h0 : dirty_0_92; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3307 = 7'h5d == index ? 1'h0 : dirty_0_93; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3308 = 7'h5e == index ? 1'h0 : dirty_0_94; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3309 = 7'h5f == index ? 1'h0 : dirty_0_95; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3310 = 7'h60 == index ? 1'h0 : dirty_0_96; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3311 = 7'h61 == index ? 1'h0 : dirty_0_97; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3312 = 7'h62 == index ? 1'h0 : dirty_0_98; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3313 = 7'h63 == index ? 1'h0 : dirty_0_99; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3314 = 7'h64 == index ? 1'h0 : dirty_0_100; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3315 = 7'h65 == index ? 1'h0 : dirty_0_101; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3316 = 7'h66 == index ? 1'h0 : dirty_0_102; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3317 = 7'h67 == index ? 1'h0 : dirty_0_103; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3318 = 7'h68 == index ? 1'h0 : dirty_0_104; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3319 = 7'h69 == index ? 1'h0 : dirty_0_105; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3320 = 7'h6a == index ? 1'h0 : dirty_0_106; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3321 = 7'h6b == index ? 1'h0 : dirty_0_107; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3322 = 7'h6c == index ? 1'h0 : dirty_0_108; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3323 = 7'h6d == index ? 1'h0 : dirty_0_109; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3324 = 7'h6e == index ? 1'h0 : dirty_0_110; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3325 = 7'h6f == index ? 1'h0 : dirty_0_111; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3326 = 7'h70 == index ? 1'h0 : dirty_0_112; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3327 = 7'h71 == index ? 1'h0 : dirty_0_113; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3328 = 7'h72 == index ? 1'h0 : dirty_0_114; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3329 = 7'h73 == index ? 1'h0 : dirty_0_115; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3330 = 7'h74 == index ? 1'h0 : dirty_0_116; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3331 = 7'h75 == index ? 1'h0 : dirty_0_117; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3332 = 7'h76 == index ? 1'h0 : dirty_0_118; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3333 = 7'h77 == index ? 1'h0 : dirty_0_119; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3334 = 7'h78 == index ? 1'h0 : dirty_0_120; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3335 = 7'h79 == index ? 1'h0 : dirty_0_121; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3336 = 7'h7a == index ? 1'h0 : dirty_0_122; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3337 = 7'h7b == index ? 1'h0 : dirty_0_123; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3338 = 7'h7c == index ? 1'h0 : dirty_0_124; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3339 = 7'h7d == index ? 1'h0 : dirty_0_125; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3340 = 7'h7e == index ? 1'h0 : dirty_0_126; // @[d_cache.scala 139:{40,40} 24:26]
  wire  _GEN_3341 = 7'h7f == index ? 1'h0 : dirty_0_127; // @[d_cache.scala 139:{40,40} 24:26]
  wire [63:0] _GEN_3854 = _GEN_645 ? _GEN_2957 : write_back_data; // @[d_cache.scala 134:47 135:41 29:34]
  wire [38:0] _GEN_3855 = _GEN_645 ? _write_back_addr_T_1 : {{7'd0}, write_back_addr}; // @[d_cache.scala 134:47 136:41 30:34]
  wire [63:0] _GEN_3856 = _GEN_645 ? _GEN_2062 : _GEN_2062; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3857 = _GEN_645 ? _GEN_2063 : _GEN_2063; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3858 = _GEN_645 ? _GEN_2064 : _GEN_2064; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3859 = _GEN_645 ? _GEN_2065 : _GEN_2065; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3860 = _GEN_645 ? _GEN_2066 : _GEN_2066; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3861 = _GEN_645 ? _GEN_2067 : _GEN_2067; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3862 = _GEN_645 ? _GEN_2068 : _GEN_2068; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3863 = _GEN_645 ? _GEN_2069 : _GEN_2069; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3864 = _GEN_645 ? _GEN_2070 : _GEN_2070; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3865 = _GEN_645 ? _GEN_2071 : _GEN_2071; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3866 = _GEN_645 ? _GEN_2072 : _GEN_2072; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3867 = _GEN_645 ? _GEN_2073 : _GEN_2073; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3868 = _GEN_645 ? _GEN_2074 : _GEN_2074; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3869 = _GEN_645 ? _GEN_2075 : _GEN_2075; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3870 = _GEN_645 ? _GEN_2076 : _GEN_2076; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3871 = _GEN_645 ? _GEN_2077 : _GEN_2077; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3872 = _GEN_645 ? _GEN_2078 : _GEN_2078; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3873 = _GEN_645 ? _GEN_2079 : _GEN_2079; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3874 = _GEN_645 ? _GEN_2080 : _GEN_2080; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3875 = _GEN_645 ? _GEN_2081 : _GEN_2081; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3876 = _GEN_645 ? _GEN_2082 : _GEN_2082; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3877 = _GEN_645 ? _GEN_2083 : _GEN_2083; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3878 = _GEN_645 ? _GEN_2084 : _GEN_2084; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3879 = _GEN_645 ? _GEN_2085 : _GEN_2085; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3880 = _GEN_645 ? _GEN_2086 : _GEN_2086; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3881 = _GEN_645 ? _GEN_2087 : _GEN_2087; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3882 = _GEN_645 ? _GEN_2088 : _GEN_2088; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3883 = _GEN_645 ? _GEN_2089 : _GEN_2089; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3884 = _GEN_645 ? _GEN_2090 : _GEN_2090; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3885 = _GEN_645 ? _GEN_2091 : _GEN_2091; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3886 = _GEN_645 ? _GEN_2092 : _GEN_2092; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3887 = _GEN_645 ? _GEN_2093 : _GEN_2093; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3888 = _GEN_645 ? _GEN_2094 : _GEN_2094; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3889 = _GEN_645 ? _GEN_2095 : _GEN_2095; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3890 = _GEN_645 ? _GEN_2096 : _GEN_2096; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3891 = _GEN_645 ? _GEN_2097 : _GEN_2097; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3892 = _GEN_645 ? _GEN_2098 : _GEN_2098; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3893 = _GEN_645 ? _GEN_2099 : _GEN_2099; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3894 = _GEN_645 ? _GEN_2100 : _GEN_2100; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3895 = _GEN_645 ? _GEN_2101 : _GEN_2101; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3896 = _GEN_645 ? _GEN_2102 : _GEN_2102; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3897 = _GEN_645 ? _GEN_2103 : _GEN_2103; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3898 = _GEN_645 ? _GEN_2104 : _GEN_2104; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3899 = _GEN_645 ? _GEN_2105 : _GEN_2105; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3900 = _GEN_645 ? _GEN_2106 : _GEN_2106; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3901 = _GEN_645 ? _GEN_2107 : _GEN_2107; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3902 = _GEN_645 ? _GEN_2108 : _GEN_2108; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3903 = _GEN_645 ? _GEN_2109 : _GEN_2109; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3904 = _GEN_645 ? _GEN_2110 : _GEN_2110; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3905 = _GEN_645 ? _GEN_2111 : _GEN_2111; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3906 = _GEN_645 ? _GEN_2112 : _GEN_2112; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3907 = _GEN_645 ? _GEN_2113 : _GEN_2113; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3908 = _GEN_645 ? _GEN_2114 : _GEN_2114; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3909 = _GEN_645 ? _GEN_2115 : _GEN_2115; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3910 = _GEN_645 ? _GEN_2116 : _GEN_2116; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3911 = _GEN_645 ? _GEN_2117 : _GEN_2117; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3912 = _GEN_645 ? _GEN_2118 : _GEN_2118; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3913 = _GEN_645 ? _GEN_2119 : _GEN_2119; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3914 = _GEN_645 ? _GEN_2120 : _GEN_2120; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3915 = _GEN_645 ? _GEN_2121 : _GEN_2121; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3916 = _GEN_645 ? _GEN_2122 : _GEN_2122; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3917 = _GEN_645 ? _GEN_2123 : _GEN_2123; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3918 = _GEN_645 ? _GEN_2124 : _GEN_2124; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3919 = _GEN_645 ? _GEN_2125 : _GEN_2125; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3920 = _GEN_645 ? _GEN_2126 : _GEN_2126; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3921 = _GEN_645 ? _GEN_2127 : _GEN_2127; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3922 = _GEN_645 ? _GEN_2128 : _GEN_2128; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3923 = _GEN_645 ? _GEN_2129 : _GEN_2129; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3924 = _GEN_645 ? _GEN_2130 : _GEN_2130; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3925 = _GEN_645 ? _GEN_2131 : _GEN_2131; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3926 = _GEN_645 ? _GEN_2132 : _GEN_2132; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3927 = _GEN_645 ? _GEN_2133 : _GEN_2133; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3928 = _GEN_645 ? _GEN_2134 : _GEN_2134; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3929 = _GEN_645 ? _GEN_2135 : _GEN_2135; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3930 = _GEN_645 ? _GEN_2136 : _GEN_2136; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3931 = _GEN_645 ? _GEN_2137 : _GEN_2137; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3932 = _GEN_645 ? _GEN_2138 : _GEN_2138; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3933 = _GEN_645 ? _GEN_2139 : _GEN_2139; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3934 = _GEN_645 ? _GEN_2140 : _GEN_2140; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3935 = _GEN_645 ? _GEN_2141 : _GEN_2141; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3936 = _GEN_645 ? _GEN_2142 : _GEN_2142; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3937 = _GEN_645 ? _GEN_2143 : _GEN_2143; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3938 = _GEN_645 ? _GEN_2144 : _GEN_2144; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3939 = _GEN_645 ? _GEN_2145 : _GEN_2145; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3940 = _GEN_645 ? _GEN_2146 : _GEN_2146; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3941 = _GEN_645 ? _GEN_2147 : _GEN_2147; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3942 = _GEN_645 ? _GEN_2148 : _GEN_2148; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3943 = _GEN_645 ? _GEN_2149 : _GEN_2149; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3944 = _GEN_645 ? _GEN_2150 : _GEN_2150; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3945 = _GEN_645 ? _GEN_2151 : _GEN_2151; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3946 = _GEN_645 ? _GEN_2152 : _GEN_2152; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3947 = _GEN_645 ? _GEN_2153 : _GEN_2153; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3948 = _GEN_645 ? _GEN_2154 : _GEN_2154; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3949 = _GEN_645 ? _GEN_2155 : _GEN_2155; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3950 = _GEN_645 ? _GEN_2156 : _GEN_2156; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3951 = _GEN_645 ? _GEN_2157 : _GEN_2157; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3952 = _GEN_645 ? _GEN_2158 : _GEN_2158; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3953 = _GEN_645 ? _GEN_2159 : _GEN_2159; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3954 = _GEN_645 ? _GEN_2160 : _GEN_2160; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3955 = _GEN_645 ? _GEN_2161 : _GEN_2161; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3956 = _GEN_645 ? _GEN_2162 : _GEN_2162; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3957 = _GEN_645 ? _GEN_2163 : _GEN_2163; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3958 = _GEN_645 ? _GEN_2164 : _GEN_2164; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3959 = _GEN_645 ? _GEN_2165 : _GEN_2165; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3960 = _GEN_645 ? _GEN_2166 : _GEN_2166; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3961 = _GEN_645 ? _GEN_2167 : _GEN_2167; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3962 = _GEN_645 ? _GEN_2168 : _GEN_2168; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3963 = _GEN_645 ? _GEN_2169 : _GEN_2169; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3964 = _GEN_645 ? _GEN_2170 : _GEN_2170; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3965 = _GEN_645 ? _GEN_2171 : _GEN_2171; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3966 = _GEN_645 ? _GEN_2172 : _GEN_2172; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3967 = _GEN_645 ? _GEN_2173 : _GEN_2173; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3968 = _GEN_645 ? _GEN_2174 : _GEN_2174; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3969 = _GEN_645 ? _GEN_2175 : _GEN_2175; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3970 = _GEN_645 ? _GEN_2176 : _GEN_2176; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3971 = _GEN_645 ? _GEN_2177 : _GEN_2177; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3972 = _GEN_645 ? _GEN_2178 : _GEN_2178; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3973 = _GEN_645 ? _GEN_2179 : _GEN_2179; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3974 = _GEN_645 ? _GEN_2180 : _GEN_2180; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3975 = _GEN_645 ? _GEN_2181 : _GEN_2181; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3976 = _GEN_645 ? _GEN_2182 : _GEN_2182; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3977 = _GEN_645 ? _GEN_2183 : _GEN_2183; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3978 = _GEN_645 ? _GEN_2184 : _GEN_2184; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3979 = _GEN_645 ? _GEN_2185 : _GEN_2185; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3980 = _GEN_645 ? _GEN_2186 : _GEN_2186; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3981 = _GEN_645 ? _GEN_2187 : _GEN_2187; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3982 = _GEN_645 ? _GEN_2188 : _GEN_2188; // @[d_cache.scala 134:47]
  wire [63:0] _GEN_3983 = _GEN_645 ? _GEN_2189 : _GEN_2189; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3984 = _GEN_645 ? _GEN_2190 : _GEN_2190; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3985 = _GEN_645 ? _GEN_2191 : _GEN_2191; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3986 = _GEN_645 ? _GEN_2192 : _GEN_2192; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3987 = _GEN_645 ? _GEN_2193 : _GEN_2193; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3988 = _GEN_645 ? _GEN_2194 : _GEN_2194; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3989 = _GEN_645 ? _GEN_2195 : _GEN_2195; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3990 = _GEN_645 ? _GEN_2196 : _GEN_2196; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3991 = _GEN_645 ? _GEN_2197 : _GEN_2197; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3992 = _GEN_645 ? _GEN_2198 : _GEN_2198; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3993 = _GEN_645 ? _GEN_2199 : _GEN_2199; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3994 = _GEN_645 ? _GEN_2200 : _GEN_2200; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3995 = _GEN_645 ? _GEN_2201 : _GEN_2201; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3996 = _GEN_645 ? _GEN_2202 : _GEN_2202; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3997 = _GEN_645 ? _GEN_2203 : _GEN_2203; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3998 = _GEN_645 ? _GEN_2204 : _GEN_2204; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_3999 = _GEN_645 ? _GEN_2205 : _GEN_2205; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4000 = _GEN_645 ? _GEN_2206 : _GEN_2206; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4001 = _GEN_645 ? _GEN_2207 : _GEN_2207; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4002 = _GEN_645 ? _GEN_2208 : _GEN_2208; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4003 = _GEN_645 ? _GEN_2209 : _GEN_2209; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4004 = _GEN_645 ? _GEN_2210 : _GEN_2210; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4005 = _GEN_645 ? _GEN_2211 : _GEN_2211; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4006 = _GEN_645 ? _GEN_2212 : _GEN_2212; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4007 = _GEN_645 ? _GEN_2213 : _GEN_2213; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4008 = _GEN_645 ? _GEN_2214 : _GEN_2214; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4009 = _GEN_645 ? _GEN_2215 : _GEN_2215; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4010 = _GEN_645 ? _GEN_2216 : _GEN_2216; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4011 = _GEN_645 ? _GEN_2217 : _GEN_2217; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4012 = _GEN_645 ? _GEN_2218 : _GEN_2218; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4013 = _GEN_645 ? _GEN_2219 : _GEN_2219; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4014 = _GEN_645 ? _GEN_2220 : _GEN_2220; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4015 = _GEN_645 ? _GEN_2221 : _GEN_2221; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4016 = _GEN_645 ? _GEN_2222 : _GEN_2222; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4017 = _GEN_645 ? _GEN_2223 : _GEN_2223; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4018 = _GEN_645 ? _GEN_2224 : _GEN_2224; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4019 = _GEN_645 ? _GEN_2225 : _GEN_2225; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4020 = _GEN_645 ? _GEN_2226 : _GEN_2226; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4021 = _GEN_645 ? _GEN_2227 : _GEN_2227; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4022 = _GEN_645 ? _GEN_2228 : _GEN_2228; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4023 = _GEN_645 ? _GEN_2229 : _GEN_2229; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4024 = _GEN_645 ? _GEN_2230 : _GEN_2230; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4025 = _GEN_645 ? _GEN_2231 : _GEN_2231; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4026 = _GEN_645 ? _GEN_2232 : _GEN_2232; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4027 = _GEN_645 ? _GEN_2233 : _GEN_2233; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4028 = _GEN_645 ? _GEN_2234 : _GEN_2234; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4029 = _GEN_645 ? _GEN_2235 : _GEN_2235; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4030 = _GEN_645 ? _GEN_2236 : _GEN_2236; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4031 = _GEN_645 ? _GEN_2237 : _GEN_2237; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4032 = _GEN_645 ? _GEN_2238 : _GEN_2238; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4033 = _GEN_645 ? _GEN_2239 : _GEN_2239; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4034 = _GEN_645 ? _GEN_2240 : _GEN_2240; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4035 = _GEN_645 ? _GEN_2241 : _GEN_2241; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4036 = _GEN_645 ? _GEN_2242 : _GEN_2242; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4037 = _GEN_645 ? _GEN_2243 : _GEN_2243; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4038 = _GEN_645 ? _GEN_2244 : _GEN_2244; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4039 = _GEN_645 ? _GEN_2245 : _GEN_2245; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4040 = _GEN_645 ? _GEN_2246 : _GEN_2246; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4041 = _GEN_645 ? _GEN_2247 : _GEN_2247; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4042 = _GEN_645 ? _GEN_2248 : _GEN_2248; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4043 = _GEN_645 ? _GEN_2249 : _GEN_2249; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4044 = _GEN_645 ? _GEN_2250 : _GEN_2250; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4045 = _GEN_645 ? _GEN_2251 : _GEN_2251; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4046 = _GEN_645 ? _GEN_2252 : _GEN_2252; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4047 = _GEN_645 ? _GEN_2253 : _GEN_2253; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4048 = _GEN_645 ? _GEN_2254 : _GEN_2254; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4049 = _GEN_645 ? _GEN_2255 : _GEN_2255; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4050 = _GEN_645 ? _GEN_2256 : _GEN_2256; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4051 = _GEN_645 ? _GEN_2257 : _GEN_2257; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4052 = _GEN_645 ? _GEN_2258 : _GEN_2258; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4053 = _GEN_645 ? _GEN_2259 : _GEN_2259; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4054 = _GEN_645 ? _GEN_2260 : _GEN_2260; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4055 = _GEN_645 ? _GEN_2261 : _GEN_2261; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4056 = _GEN_645 ? _GEN_2262 : _GEN_2262; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4057 = _GEN_645 ? _GEN_2263 : _GEN_2263; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4058 = _GEN_645 ? _GEN_2264 : _GEN_2264; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4059 = _GEN_645 ? _GEN_2265 : _GEN_2265; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4060 = _GEN_645 ? _GEN_2266 : _GEN_2266; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4061 = _GEN_645 ? _GEN_2267 : _GEN_2267; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4062 = _GEN_645 ? _GEN_2268 : _GEN_2268; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4063 = _GEN_645 ? _GEN_2269 : _GEN_2269; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4064 = _GEN_645 ? _GEN_2270 : _GEN_2270; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4065 = _GEN_645 ? _GEN_2271 : _GEN_2271; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4066 = _GEN_645 ? _GEN_2272 : _GEN_2272; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4067 = _GEN_645 ? _GEN_2273 : _GEN_2273; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4068 = _GEN_645 ? _GEN_2274 : _GEN_2274; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4069 = _GEN_645 ? _GEN_2275 : _GEN_2275; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4070 = _GEN_645 ? _GEN_2276 : _GEN_2276; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4071 = _GEN_645 ? _GEN_2277 : _GEN_2277; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4072 = _GEN_645 ? _GEN_2278 : _GEN_2278; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4073 = _GEN_645 ? _GEN_2279 : _GEN_2279; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4074 = _GEN_645 ? _GEN_2280 : _GEN_2280; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4075 = _GEN_645 ? _GEN_2281 : _GEN_2281; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4076 = _GEN_645 ? _GEN_2282 : _GEN_2282; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4077 = _GEN_645 ? _GEN_2283 : _GEN_2283; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4078 = _GEN_645 ? _GEN_2284 : _GEN_2284; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4079 = _GEN_645 ? _GEN_2285 : _GEN_2285; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4080 = _GEN_645 ? _GEN_2286 : _GEN_2286; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4081 = _GEN_645 ? _GEN_2287 : _GEN_2287; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4082 = _GEN_645 ? _GEN_2288 : _GEN_2288; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4083 = _GEN_645 ? _GEN_2289 : _GEN_2289; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4084 = _GEN_645 ? _GEN_2290 : _GEN_2290; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4085 = _GEN_645 ? _GEN_2291 : _GEN_2291; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4086 = _GEN_645 ? _GEN_2292 : _GEN_2292; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4087 = _GEN_645 ? _GEN_2293 : _GEN_2293; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4088 = _GEN_645 ? _GEN_2294 : _GEN_2294; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4089 = _GEN_645 ? _GEN_2295 : _GEN_2295; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4090 = _GEN_645 ? _GEN_2296 : _GEN_2296; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4091 = _GEN_645 ? _GEN_2297 : _GEN_2297; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4092 = _GEN_645 ? _GEN_2298 : _GEN_2298; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4093 = _GEN_645 ? _GEN_2299 : _GEN_2299; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4094 = _GEN_645 ? _GEN_2300 : _GEN_2300; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4095 = _GEN_645 ? _GEN_2301 : _GEN_2301; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4096 = _GEN_645 ? _GEN_2302 : _GEN_2302; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4097 = _GEN_645 ? _GEN_2303 : _GEN_2303; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4098 = _GEN_645 ? _GEN_2304 : _GEN_2304; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4099 = _GEN_645 ? _GEN_2305 : _GEN_2305; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4100 = _GEN_645 ? _GEN_2306 : _GEN_2306; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4101 = _GEN_645 ? _GEN_2307 : _GEN_2307; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4102 = _GEN_645 ? _GEN_2308 : _GEN_2308; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4103 = _GEN_645 ? _GEN_2309 : _GEN_2309; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4104 = _GEN_645 ? _GEN_2310 : _GEN_2310; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4105 = _GEN_645 ? _GEN_2311 : _GEN_2311; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4106 = _GEN_645 ? _GEN_2312 : _GEN_2312; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4107 = _GEN_645 ? _GEN_2313 : _GEN_2313; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4108 = _GEN_645 ? _GEN_2314 : _GEN_2314; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4109 = _GEN_645 ? _GEN_2315 : _GEN_2315; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4110 = _GEN_645 ? _GEN_2316 : _GEN_2316; // @[d_cache.scala 134:47]
  wire [31:0] _GEN_4111 = _GEN_645 ? _GEN_2317 : _GEN_2317; // @[d_cache.scala 134:47]
  wire  _GEN_4112 = _GEN_645 ? _GEN_3214 : dirty_0_0; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4113 = _GEN_645 ? _GEN_3215 : dirty_0_1; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4114 = _GEN_645 ? _GEN_3216 : dirty_0_2; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4115 = _GEN_645 ? _GEN_3217 : dirty_0_3; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4116 = _GEN_645 ? _GEN_3218 : dirty_0_4; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4117 = _GEN_645 ? _GEN_3219 : dirty_0_5; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4118 = _GEN_645 ? _GEN_3220 : dirty_0_6; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4119 = _GEN_645 ? _GEN_3221 : dirty_0_7; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4120 = _GEN_645 ? _GEN_3222 : dirty_0_8; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4121 = _GEN_645 ? _GEN_3223 : dirty_0_9; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4122 = _GEN_645 ? _GEN_3224 : dirty_0_10; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4123 = _GEN_645 ? _GEN_3225 : dirty_0_11; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4124 = _GEN_645 ? _GEN_3226 : dirty_0_12; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4125 = _GEN_645 ? _GEN_3227 : dirty_0_13; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4126 = _GEN_645 ? _GEN_3228 : dirty_0_14; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4127 = _GEN_645 ? _GEN_3229 : dirty_0_15; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4128 = _GEN_645 ? _GEN_3230 : dirty_0_16; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4129 = _GEN_645 ? _GEN_3231 : dirty_0_17; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4130 = _GEN_645 ? _GEN_3232 : dirty_0_18; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4131 = _GEN_645 ? _GEN_3233 : dirty_0_19; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4132 = _GEN_645 ? _GEN_3234 : dirty_0_20; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4133 = _GEN_645 ? _GEN_3235 : dirty_0_21; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4134 = _GEN_645 ? _GEN_3236 : dirty_0_22; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4135 = _GEN_645 ? _GEN_3237 : dirty_0_23; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4136 = _GEN_645 ? _GEN_3238 : dirty_0_24; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4137 = _GEN_645 ? _GEN_3239 : dirty_0_25; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4138 = _GEN_645 ? _GEN_3240 : dirty_0_26; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4139 = _GEN_645 ? _GEN_3241 : dirty_0_27; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4140 = _GEN_645 ? _GEN_3242 : dirty_0_28; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4141 = _GEN_645 ? _GEN_3243 : dirty_0_29; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4142 = _GEN_645 ? _GEN_3244 : dirty_0_30; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4143 = _GEN_645 ? _GEN_3245 : dirty_0_31; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4144 = _GEN_645 ? _GEN_3246 : dirty_0_32; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4145 = _GEN_645 ? _GEN_3247 : dirty_0_33; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4146 = _GEN_645 ? _GEN_3248 : dirty_0_34; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4147 = _GEN_645 ? _GEN_3249 : dirty_0_35; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4148 = _GEN_645 ? _GEN_3250 : dirty_0_36; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4149 = _GEN_645 ? _GEN_3251 : dirty_0_37; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4150 = _GEN_645 ? _GEN_3252 : dirty_0_38; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4151 = _GEN_645 ? _GEN_3253 : dirty_0_39; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4152 = _GEN_645 ? _GEN_3254 : dirty_0_40; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4153 = _GEN_645 ? _GEN_3255 : dirty_0_41; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4154 = _GEN_645 ? _GEN_3256 : dirty_0_42; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4155 = _GEN_645 ? _GEN_3257 : dirty_0_43; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4156 = _GEN_645 ? _GEN_3258 : dirty_0_44; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4157 = _GEN_645 ? _GEN_3259 : dirty_0_45; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4158 = _GEN_645 ? _GEN_3260 : dirty_0_46; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4159 = _GEN_645 ? _GEN_3261 : dirty_0_47; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4160 = _GEN_645 ? _GEN_3262 : dirty_0_48; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4161 = _GEN_645 ? _GEN_3263 : dirty_0_49; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4162 = _GEN_645 ? _GEN_3264 : dirty_0_50; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4163 = _GEN_645 ? _GEN_3265 : dirty_0_51; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4164 = _GEN_645 ? _GEN_3266 : dirty_0_52; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4165 = _GEN_645 ? _GEN_3267 : dirty_0_53; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4166 = _GEN_645 ? _GEN_3268 : dirty_0_54; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4167 = _GEN_645 ? _GEN_3269 : dirty_0_55; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4168 = _GEN_645 ? _GEN_3270 : dirty_0_56; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4169 = _GEN_645 ? _GEN_3271 : dirty_0_57; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4170 = _GEN_645 ? _GEN_3272 : dirty_0_58; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4171 = _GEN_645 ? _GEN_3273 : dirty_0_59; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4172 = _GEN_645 ? _GEN_3274 : dirty_0_60; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4173 = _GEN_645 ? _GEN_3275 : dirty_0_61; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4174 = _GEN_645 ? _GEN_3276 : dirty_0_62; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4175 = _GEN_645 ? _GEN_3277 : dirty_0_63; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4176 = _GEN_645 ? _GEN_3278 : dirty_0_64; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4177 = _GEN_645 ? _GEN_3279 : dirty_0_65; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4178 = _GEN_645 ? _GEN_3280 : dirty_0_66; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4179 = _GEN_645 ? _GEN_3281 : dirty_0_67; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4180 = _GEN_645 ? _GEN_3282 : dirty_0_68; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4181 = _GEN_645 ? _GEN_3283 : dirty_0_69; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4182 = _GEN_645 ? _GEN_3284 : dirty_0_70; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4183 = _GEN_645 ? _GEN_3285 : dirty_0_71; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4184 = _GEN_645 ? _GEN_3286 : dirty_0_72; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4185 = _GEN_645 ? _GEN_3287 : dirty_0_73; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4186 = _GEN_645 ? _GEN_3288 : dirty_0_74; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4187 = _GEN_645 ? _GEN_3289 : dirty_0_75; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4188 = _GEN_645 ? _GEN_3290 : dirty_0_76; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4189 = _GEN_645 ? _GEN_3291 : dirty_0_77; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4190 = _GEN_645 ? _GEN_3292 : dirty_0_78; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4191 = _GEN_645 ? _GEN_3293 : dirty_0_79; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4192 = _GEN_645 ? _GEN_3294 : dirty_0_80; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4193 = _GEN_645 ? _GEN_3295 : dirty_0_81; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4194 = _GEN_645 ? _GEN_3296 : dirty_0_82; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4195 = _GEN_645 ? _GEN_3297 : dirty_0_83; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4196 = _GEN_645 ? _GEN_3298 : dirty_0_84; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4197 = _GEN_645 ? _GEN_3299 : dirty_0_85; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4198 = _GEN_645 ? _GEN_3300 : dirty_0_86; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4199 = _GEN_645 ? _GEN_3301 : dirty_0_87; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4200 = _GEN_645 ? _GEN_3302 : dirty_0_88; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4201 = _GEN_645 ? _GEN_3303 : dirty_0_89; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4202 = _GEN_645 ? _GEN_3304 : dirty_0_90; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4203 = _GEN_645 ? _GEN_3305 : dirty_0_91; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4204 = _GEN_645 ? _GEN_3306 : dirty_0_92; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4205 = _GEN_645 ? _GEN_3307 : dirty_0_93; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4206 = _GEN_645 ? _GEN_3308 : dirty_0_94; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4207 = _GEN_645 ? _GEN_3309 : dirty_0_95; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4208 = _GEN_645 ? _GEN_3310 : dirty_0_96; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4209 = _GEN_645 ? _GEN_3311 : dirty_0_97; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4210 = _GEN_645 ? _GEN_3312 : dirty_0_98; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4211 = _GEN_645 ? _GEN_3313 : dirty_0_99; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4212 = _GEN_645 ? _GEN_3314 : dirty_0_100; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4213 = _GEN_645 ? _GEN_3315 : dirty_0_101; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4214 = _GEN_645 ? _GEN_3316 : dirty_0_102; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4215 = _GEN_645 ? _GEN_3317 : dirty_0_103; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4216 = _GEN_645 ? _GEN_3318 : dirty_0_104; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4217 = _GEN_645 ? _GEN_3319 : dirty_0_105; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4218 = _GEN_645 ? _GEN_3320 : dirty_0_106; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4219 = _GEN_645 ? _GEN_3321 : dirty_0_107; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4220 = _GEN_645 ? _GEN_3322 : dirty_0_108; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4221 = _GEN_645 ? _GEN_3323 : dirty_0_109; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4222 = _GEN_645 ? _GEN_3324 : dirty_0_110; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4223 = _GEN_645 ? _GEN_3325 : dirty_0_111; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4224 = _GEN_645 ? _GEN_3326 : dirty_0_112; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4225 = _GEN_645 ? _GEN_3327 : dirty_0_113; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4226 = _GEN_645 ? _GEN_3328 : dirty_0_114; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4227 = _GEN_645 ? _GEN_3329 : dirty_0_115; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4228 = _GEN_645 ? _GEN_3330 : dirty_0_116; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4229 = _GEN_645 ? _GEN_3331 : dirty_0_117; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4230 = _GEN_645 ? _GEN_3332 : dirty_0_118; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4231 = _GEN_645 ? _GEN_3333 : dirty_0_119; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4232 = _GEN_645 ? _GEN_3334 : dirty_0_120; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4233 = _GEN_645 ? _GEN_3335 : dirty_0_121; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4234 = _GEN_645 ? _GEN_3336 : dirty_0_122; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4235 = _GEN_645 ? _GEN_3337 : dirty_0_123; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4236 = _GEN_645 ? _GEN_3338 : dirty_0_124; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4237 = _GEN_645 ? _GEN_3339 : dirty_0_125; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4238 = _GEN_645 ? _GEN_3340 : dirty_0_126; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4239 = _GEN_645 ? _GEN_3341 : dirty_0_127; // @[d_cache.scala 134:47 24:26]
  wire  _GEN_4240 = _GEN_645 ? _GEN_2318 : _GEN_2318; // @[d_cache.scala 134:47]
  wire  _GEN_4241 = _GEN_645 ? _GEN_2319 : _GEN_2319; // @[d_cache.scala 134:47]
  wire  _GEN_4242 = _GEN_645 ? _GEN_2320 : _GEN_2320; // @[d_cache.scala 134:47]
  wire  _GEN_4243 = _GEN_645 ? _GEN_2321 : _GEN_2321; // @[d_cache.scala 134:47]
  wire  _GEN_4244 = _GEN_645 ? _GEN_2322 : _GEN_2322; // @[d_cache.scala 134:47]
  wire  _GEN_4245 = _GEN_645 ? _GEN_2323 : _GEN_2323; // @[d_cache.scala 134:47]
  wire  _GEN_4246 = _GEN_645 ? _GEN_2324 : _GEN_2324; // @[d_cache.scala 134:47]
  wire  _GEN_4247 = _GEN_645 ? _GEN_2325 : _GEN_2325; // @[d_cache.scala 134:47]
  wire  _GEN_4248 = _GEN_645 ? _GEN_2326 : _GEN_2326; // @[d_cache.scala 134:47]
  wire  _GEN_4249 = _GEN_645 ? _GEN_2327 : _GEN_2327; // @[d_cache.scala 134:47]
  wire  _GEN_4250 = _GEN_645 ? _GEN_2328 : _GEN_2328; // @[d_cache.scala 134:47]
  wire  _GEN_4251 = _GEN_645 ? _GEN_2329 : _GEN_2329; // @[d_cache.scala 134:47]
  wire  _GEN_4252 = _GEN_645 ? _GEN_2330 : _GEN_2330; // @[d_cache.scala 134:47]
  wire  _GEN_4253 = _GEN_645 ? _GEN_2331 : _GEN_2331; // @[d_cache.scala 134:47]
  wire  _GEN_4254 = _GEN_645 ? _GEN_2332 : _GEN_2332; // @[d_cache.scala 134:47]
  wire  _GEN_4255 = _GEN_645 ? _GEN_2333 : _GEN_2333; // @[d_cache.scala 134:47]
  wire  _GEN_4256 = _GEN_645 ? _GEN_2334 : _GEN_2334; // @[d_cache.scala 134:47]
  wire  _GEN_4257 = _GEN_645 ? _GEN_2335 : _GEN_2335; // @[d_cache.scala 134:47]
  wire  _GEN_4258 = _GEN_645 ? _GEN_2336 : _GEN_2336; // @[d_cache.scala 134:47]
  wire  _GEN_4259 = _GEN_645 ? _GEN_2337 : _GEN_2337; // @[d_cache.scala 134:47]
  wire  _GEN_4260 = _GEN_645 ? _GEN_2338 : _GEN_2338; // @[d_cache.scala 134:47]
  wire  _GEN_4261 = _GEN_645 ? _GEN_2339 : _GEN_2339; // @[d_cache.scala 134:47]
  wire  _GEN_4262 = _GEN_645 ? _GEN_2340 : _GEN_2340; // @[d_cache.scala 134:47]
  wire  _GEN_4263 = _GEN_645 ? _GEN_2341 : _GEN_2341; // @[d_cache.scala 134:47]
  wire  _GEN_4264 = _GEN_645 ? _GEN_2342 : _GEN_2342; // @[d_cache.scala 134:47]
  wire  _GEN_4265 = _GEN_645 ? _GEN_2343 : _GEN_2343; // @[d_cache.scala 134:47]
  wire  _GEN_4266 = _GEN_645 ? _GEN_2344 : _GEN_2344; // @[d_cache.scala 134:47]
  wire  _GEN_4267 = _GEN_645 ? _GEN_2345 : _GEN_2345; // @[d_cache.scala 134:47]
  wire  _GEN_4268 = _GEN_645 ? _GEN_2346 : _GEN_2346; // @[d_cache.scala 134:47]
  wire  _GEN_4269 = _GEN_645 ? _GEN_2347 : _GEN_2347; // @[d_cache.scala 134:47]
  wire  _GEN_4270 = _GEN_645 ? _GEN_2348 : _GEN_2348; // @[d_cache.scala 134:47]
  wire  _GEN_4271 = _GEN_645 ? _GEN_2349 : _GEN_2349; // @[d_cache.scala 134:47]
  wire  _GEN_4272 = _GEN_645 ? _GEN_2350 : _GEN_2350; // @[d_cache.scala 134:47]
  wire  _GEN_4273 = _GEN_645 ? _GEN_2351 : _GEN_2351; // @[d_cache.scala 134:47]
  wire  _GEN_4274 = _GEN_645 ? _GEN_2352 : _GEN_2352; // @[d_cache.scala 134:47]
  wire  _GEN_4275 = _GEN_645 ? _GEN_2353 : _GEN_2353; // @[d_cache.scala 134:47]
  wire  _GEN_4276 = _GEN_645 ? _GEN_2354 : _GEN_2354; // @[d_cache.scala 134:47]
  wire  _GEN_4277 = _GEN_645 ? _GEN_2355 : _GEN_2355; // @[d_cache.scala 134:47]
  wire  _GEN_4278 = _GEN_645 ? _GEN_2356 : _GEN_2356; // @[d_cache.scala 134:47]
  wire  _GEN_4279 = _GEN_645 ? _GEN_2357 : _GEN_2357; // @[d_cache.scala 134:47]
  wire  _GEN_4280 = _GEN_645 ? _GEN_2358 : _GEN_2358; // @[d_cache.scala 134:47]
  wire  _GEN_4281 = _GEN_645 ? _GEN_2359 : _GEN_2359; // @[d_cache.scala 134:47]
  wire  _GEN_4282 = _GEN_645 ? _GEN_2360 : _GEN_2360; // @[d_cache.scala 134:47]
  wire  _GEN_4283 = _GEN_645 ? _GEN_2361 : _GEN_2361; // @[d_cache.scala 134:47]
  wire  _GEN_4284 = _GEN_645 ? _GEN_2362 : _GEN_2362; // @[d_cache.scala 134:47]
  wire  _GEN_4285 = _GEN_645 ? _GEN_2363 : _GEN_2363; // @[d_cache.scala 134:47]
  wire  _GEN_4286 = _GEN_645 ? _GEN_2364 : _GEN_2364; // @[d_cache.scala 134:47]
  wire  _GEN_4287 = _GEN_645 ? _GEN_2365 : _GEN_2365; // @[d_cache.scala 134:47]
  wire  _GEN_4288 = _GEN_645 ? _GEN_2366 : _GEN_2366; // @[d_cache.scala 134:47]
  wire  _GEN_4289 = _GEN_645 ? _GEN_2367 : _GEN_2367; // @[d_cache.scala 134:47]
  wire  _GEN_4290 = _GEN_645 ? _GEN_2368 : _GEN_2368; // @[d_cache.scala 134:47]
  wire  _GEN_4291 = _GEN_645 ? _GEN_2369 : _GEN_2369; // @[d_cache.scala 134:47]
  wire  _GEN_4292 = _GEN_645 ? _GEN_2370 : _GEN_2370; // @[d_cache.scala 134:47]
  wire  _GEN_4293 = _GEN_645 ? _GEN_2371 : _GEN_2371; // @[d_cache.scala 134:47]
  wire  _GEN_4294 = _GEN_645 ? _GEN_2372 : _GEN_2372; // @[d_cache.scala 134:47]
  wire  _GEN_4295 = _GEN_645 ? _GEN_2373 : _GEN_2373; // @[d_cache.scala 134:47]
  wire  _GEN_4296 = _GEN_645 ? _GEN_2374 : _GEN_2374; // @[d_cache.scala 134:47]
  wire  _GEN_4297 = _GEN_645 ? _GEN_2375 : _GEN_2375; // @[d_cache.scala 134:47]
  wire  _GEN_4298 = _GEN_645 ? _GEN_2376 : _GEN_2376; // @[d_cache.scala 134:47]
  wire  _GEN_4299 = _GEN_645 ? _GEN_2377 : _GEN_2377; // @[d_cache.scala 134:47]
  wire  _GEN_4300 = _GEN_645 ? _GEN_2378 : _GEN_2378; // @[d_cache.scala 134:47]
  wire  _GEN_4301 = _GEN_645 ? _GEN_2379 : _GEN_2379; // @[d_cache.scala 134:47]
  wire  _GEN_4302 = _GEN_645 ? _GEN_2380 : _GEN_2380; // @[d_cache.scala 134:47]
  wire  _GEN_4303 = _GEN_645 ? _GEN_2381 : _GEN_2381; // @[d_cache.scala 134:47]
  wire  _GEN_4304 = _GEN_645 ? _GEN_2382 : _GEN_2382; // @[d_cache.scala 134:47]
  wire  _GEN_4305 = _GEN_645 ? _GEN_2383 : _GEN_2383; // @[d_cache.scala 134:47]
  wire  _GEN_4306 = _GEN_645 ? _GEN_2384 : _GEN_2384; // @[d_cache.scala 134:47]
  wire  _GEN_4307 = _GEN_645 ? _GEN_2385 : _GEN_2385; // @[d_cache.scala 134:47]
  wire  _GEN_4308 = _GEN_645 ? _GEN_2386 : _GEN_2386; // @[d_cache.scala 134:47]
  wire  _GEN_4309 = _GEN_645 ? _GEN_2387 : _GEN_2387; // @[d_cache.scala 134:47]
  wire  _GEN_4310 = _GEN_645 ? _GEN_2388 : _GEN_2388; // @[d_cache.scala 134:47]
  wire  _GEN_4311 = _GEN_645 ? _GEN_2389 : _GEN_2389; // @[d_cache.scala 134:47]
  wire  _GEN_4312 = _GEN_645 ? _GEN_2390 : _GEN_2390; // @[d_cache.scala 134:47]
  wire  _GEN_4313 = _GEN_645 ? _GEN_2391 : _GEN_2391; // @[d_cache.scala 134:47]
  wire  _GEN_4314 = _GEN_645 ? _GEN_2392 : _GEN_2392; // @[d_cache.scala 134:47]
  wire  _GEN_4315 = _GEN_645 ? _GEN_2393 : _GEN_2393; // @[d_cache.scala 134:47]
  wire  _GEN_4316 = _GEN_645 ? _GEN_2394 : _GEN_2394; // @[d_cache.scala 134:47]
  wire  _GEN_4317 = _GEN_645 ? _GEN_2395 : _GEN_2395; // @[d_cache.scala 134:47]
  wire  _GEN_4318 = _GEN_645 ? _GEN_2396 : _GEN_2396; // @[d_cache.scala 134:47]
  wire  _GEN_4319 = _GEN_645 ? _GEN_2397 : _GEN_2397; // @[d_cache.scala 134:47]
  wire  _GEN_4320 = _GEN_645 ? _GEN_2398 : _GEN_2398; // @[d_cache.scala 134:47]
  wire  _GEN_4321 = _GEN_645 ? _GEN_2399 : _GEN_2399; // @[d_cache.scala 134:47]
  wire  _GEN_4322 = _GEN_645 ? _GEN_2400 : _GEN_2400; // @[d_cache.scala 134:47]
  wire  _GEN_4323 = _GEN_645 ? _GEN_2401 : _GEN_2401; // @[d_cache.scala 134:47]
  wire  _GEN_4324 = _GEN_645 ? _GEN_2402 : _GEN_2402; // @[d_cache.scala 134:47]
  wire  _GEN_4325 = _GEN_645 ? _GEN_2403 : _GEN_2403; // @[d_cache.scala 134:47]
  wire  _GEN_4326 = _GEN_645 ? _GEN_2404 : _GEN_2404; // @[d_cache.scala 134:47]
  wire  _GEN_4327 = _GEN_645 ? _GEN_2405 : _GEN_2405; // @[d_cache.scala 134:47]
  wire  _GEN_4328 = _GEN_645 ? _GEN_2406 : _GEN_2406; // @[d_cache.scala 134:47]
  wire  _GEN_4329 = _GEN_645 ? _GEN_2407 : _GEN_2407; // @[d_cache.scala 134:47]
  wire  _GEN_4330 = _GEN_645 ? _GEN_2408 : _GEN_2408; // @[d_cache.scala 134:47]
  wire  _GEN_4331 = _GEN_645 ? _GEN_2409 : _GEN_2409; // @[d_cache.scala 134:47]
  wire  _GEN_4332 = _GEN_645 ? _GEN_2410 : _GEN_2410; // @[d_cache.scala 134:47]
  wire  _GEN_4333 = _GEN_645 ? _GEN_2411 : _GEN_2411; // @[d_cache.scala 134:47]
  wire  _GEN_4334 = _GEN_645 ? _GEN_2412 : _GEN_2412; // @[d_cache.scala 134:47]
  wire  _GEN_4335 = _GEN_645 ? _GEN_2413 : _GEN_2413; // @[d_cache.scala 134:47]
  wire  _GEN_4336 = _GEN_645 ? _GEN_2414 : _GEN_2414; // @[d_cache.scala 134:47]
  wire  _GEN_4337 = _GEN_645 ? _GEN_2415 : _GEN_2415; // @[d_cache.scala 134:47]
  wire  _GEN_4338 = _GEN_645 ? _GEN_2416 : _GEN_2416; // @[d_cache.scala 134:47]
  wire  _GEN_4339 = _GEN_645 ? _GEN_2417 : _GEN_2417; // @[d_cache.scala 134:47]
  wire  _GEN_4340 = _GEN_645 ? _GEN_2418 : _GEN_2418; // @[d_cache.scala 134:47]
  wire  _GEN_4341 = _GEN_645 ? _GEN_2419 : _GEN_2419; // @[d_cache.scala 134:47]
  wire  _GEN_4342 = _GEN_645 ? _GEN_2420 : _GEN_2420; // @[d_cache.scala 134:47]
  wire  _GEN_4343 = _GEN_645 ? _GEN_2421 : _GEN_2421; // @[d_cache.scala 134:47]
  wire  _GEN_4344 = _GEN_645 ? _GEN_2422 : _GEN_2422; // @[d_cache.scala 134:47]
  wire  _GEN_4345 = _GEN_645 ? _GEN_2423 : _GEN_2423; // @[d_cache.scala 134:47]
  wire  _GEN_4346 = _GEN_645 ? _GEN_2424 : _GEN_2424; // @[d_cache.scala 134:47]
  wire  _GEN_4347 = _GEN_645 ? _GEN_2425 : _GEN_2425; // @[d_cache.scala 134:47]
  wire  _GEN_4348 = _GEN_645 ? _GEN_2426 : _GEN_2426; // @[d_cache.scala 134:47]
  wire  _GEN_4349 = _GEN_645 ? _GEN_2427 : _GEN_2427; // @[d_cache.scala 134:47]
  wire  _GEN_4350 = _GEN_645 ? _GEN_2428 : _GEN_2428; // @[d_cache.scala 134:47]
  wire  _GEN_4351 = _GEN_645 ? _GEN_2429 : _GEN_2429; // @[d_cache.scala 134:47]
  wire  _GEN_4352 = _GEN_645 ? _GEN_2430 : _GEN_2430; // @[d_cache.scala 134:47]
  wire  _GEN_4353 = _GEN_645 ? _GEN_2431 : _GEN_2431; // @[d_cache.scala 134:47]
  wire  _GEN_4354 = _GEN_645 ? _GEN_2432 : _GEN_2432; // @[d_cache.scala 134:47]
  wire  _GEN_4355 = _GEN_645 ? _GEN_2433 : _GEN_2433; // @[d_cache.scala 134:47]
  wire  _GEN_4356 = _GEN_645 ? _GEN_2434 : _GEN_2434; // @[d_cache.scala 134:47]
  wire  _GEN_4357 = _GEN_645 ? _GEN_2435 : _GEN_2435; // @[d_cache.scala 134:47]
  wire  _GEN_4358 = _GEN_645 ? _GEN_2436 : _GEN_2436; // @[d_cache.scala 134:47]
  wire  _GEN_4359 = _GEN_645 ? _GEN_2437 : _GEN_2437; // @[d_cache.scala 134:47]
  wire  _GEN_4360 = _GEN_645 ? _GEN_2438 : _GEN_2438; // @[d_cache.scala 134:47]
  wire  _GEN_4361 = _GEN_645 ? _GEN_2439 : _GEN_2439; // @[d_cache.scala 134:47]
  wire  _GEN_4362 = _GEN_645 ? _GEN_2440 : _GEN_2440; // @[d_cache.scala 134:47]
  wire  _GEN_4363 = _GEN_645 ? _GEN_2441 : _GEN_2441; // @[d_cache.scala 134:47]
  wire  _GEN_4364 = _GEN_645 ? _GEN_2442 : _GEN_2442; // @[d_cache.scala 134:47]
  wire  _GEN_4365 = _GEN_645 ? _GEN_2443 : _GEN_2443; // @[d_cache.scala 134:47]
  wire  _GEN_4366 = _GEN_645 ? _GEN_2444 : _GEN_2444; // @[d_cache.scala 134:47]
  wire  _GEN_4367 = _GEN_645 ? _GEN_2445 : _GEN_2445; // @[d_cache.scala 134:47]
  wire [2:0] _GEN_4368 = _GEN_645 ? 3'h6 : 3'h7; // @[d_cache.scala 134:47 141:31 144:31]
  wire [63:0] _GEN_4371 = 7'h1 == index ? ram_1_1 : ram_1_0; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4372 = 7'h2 == index ? ram_1_2 : _GEN_4371; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4373 = 7'h3 == index ? ram_1_3 : _GEN_4372; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4374 = 7'h4 == index ? ram_1_4 : _GEN_4373; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4375 = 7'h5 == index ? ram_1_5 : _GEN_4374; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4376 = 7'h6 == index ? ram_1_6 : _GEN_4375; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4377 = 7'h7 == index ? ram_1_7 : _GEN_4376; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4378 = 7'h8 == index ? ram_1_8 : _GEN_4377; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4379 = 7'h9 == index ? ram_1_9 : _GEN_4378; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4380 = 7'ha == index ? ram_1_10 : _GEN_4379; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4381 = 7'hb == index ? ram_1_11 : _GEN_4380; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4382 = 7'hc == index ? ram_1_12 : _GEN_4381; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4383 = 7'hd == index ? ram_1_13 : _GEN_4382; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4384 = 7'he == index ? ram_1_14 : _GEN_4383; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4385 = 7'hf == index ? ram_1_15 : _GEN_4384; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4386 = 7'h10 == index ? ram_1_16 : _GEN_4385; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4387 = 7'h11 == index ? ram_1_17 : _GEN_4386; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4388 = 7'h12 == index ? ram_1_18 : _GEN_4387; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4389 = 7'h13 == index ? ram_1_19 : _GEN_4388; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4390 = 7'h14 == index ? ram_1_20 : _GEN_4389; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4391 = 7'h15 == index ? ram_1_21 : _GEN_4390; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4392 = 7'h16 == index ? ram_1_22 : _GEN_4391; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4393 = 7'h17 == index ? ram_1_23 : _GEN_4392; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4394 = 7'h18 == index ? ram_1_24 : _GEN_4393; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4395 = 7'h19 == index ? ram_1_25 : _GEN_4394; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4396 = 7'h1a == index ? ram_1_26 : _GEN_4395; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4397 = 7'h1b == index ? ram_1_27 : _GEN_4396; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4398 = 7'h1c == index ? ram_1_28 : _GEN_4397; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4399 = 7'h1d == index ? ram_1_29 : _GEN_4398; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4400 = 7'h1e == index ? ram_1_30 : _GEN_4399; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4401 = 7'h1f == index ? ram_1_31 : _GEN_4400; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4402 = 7'h20 == index ? ram_1_32 : _GEN_4401; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4403 = 7'h21 == index ? ram_1_33 : _GEN_4402; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4404 = 7'h22 == index ? ram_1_34 : _GEN_4403; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4405 = 7'h23 == index ? ram_1_35 : _GEN_4404; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4406 = 7'h24 == index ? ram_1_36 : _GEN_4405; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4407 = 7'h25 == index ? ram_1_37 : _GEN_4406; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4408 = 7'h26 == index ? ram_1_38 : _GEN_4407; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4409 = 7'h27 == index ? ram_1_39 : _GEN_4408; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4410 = 7'h28 == index ? ram_1_40 : _GEN_4409; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4411 = 7'h29 == index ? ram_1_41 : _GEN_4410; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4412 = 7'h2a == index ? ram_1_42 : _GEN_4411; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4413 = 7'h2b == index ? ram_1_43 : _GEN_4412; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4414 = 7'h2c == index ? ram_1_44 : _GEN_4413; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4415 = 7'h2d == index ? ram_1_45 : _GEN_4414; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4416 = 7'h2e == index ? ram_1_46 : _GEN_4415; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4417 = 7'h2f == index ? ram_1_47 : _GEN_4416; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4418 = 7'h30 == index ? ram_1_48 : _GEN_4417; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4419 = 7'h31 == index ? ram_1_49 : _GEN_4418; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4420 = 7'h32 == index ? ram_1_50 : _GEN_4419; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4421 = 7'h33 == index ? ram_1_51 : _GEN_4420; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4422 = 7'h34 == index ? ram_1_52 : _GEN_4421; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4423 = 7'h35 == index ? ram_1_53 : _GEN_4422; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4424 = 7'h36 == index ? ram_1_54 : _GEN_4423; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4425 = 7'h37 == index ? ram_1_55 : _GEN_4424; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4426 = 7'h38 == index ? ram_1_56 : _GEN_4425; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4427 = 7'h39 == index ? ram_1_57 : _GEN_4426; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4428 = 7'h3a == index ? ram_1_58 : _GEN_4427; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4429 = 7'h3b == index ? ram_1_59 : _GEN_4428; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4430 = 7'h3c == index ? ram_1_60 : _GEN_4429; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4431 = 7'h3d == index ? ram_1_61 : _GEN_4430; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4432 = 7'h3e == index ? ram_1_62 : _GEN_4431; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4433 = 7'h3f == index ? ram_1_63 : _GEN_4432; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4434 = 7'h40 == index ? ram_1_64 : _GEN_4433; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4435 = 7'h41 == index ? ram_1_65 : _GEN_4434; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4436 = 7'h42 == index ? ram_1_66 : _GEN_4435; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4437 = 7'h43 == index ? ram_1_67 : _GEN_4436; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4438 = 7'h44 == index ? ram_1_68 : _GEN_4437; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4439 = 7'h45 == index ? ram_1_69 : _GEN_4438; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4440 = 7'h46 == index ? ram_1_70 : _GEN_4439; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4441 = 7'h47 == index ? ram_1_71 : _GEN_4440; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4442 = 7'h48 == index ? ram_1_72 : _GEN_4441; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4443 = 7'h49 == index ? ram_1_73 : _GEN_4442; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4444 = 7'h4a == index ? ram_1_74 : _GEN_4443; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4445 = 7'h4b == index ? ram_1_75 : _GEN_4444; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4446 = 7'h4c == index ? ram_1_76 : _GEN_4445; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4447 = 7'h4d == index ? ram_1_77 : _GEN_4446; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4448 = 7'h4e == index ? ram_1_78 : _GEN_4447; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4449 = 7'h4f == index ? ram_1_79 : _GEN_4448; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4450 = 7'h50 == index ? ram_1_80 : _GEN_4449; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4451 = 7'h51 == index ? ram_1_81 : _GEN_4450; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4452 = 7'h52 == index ? ram_1_82 : _GEN_4451; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4453 = 7'h53 == index ? ram_1_83 : _GEN_4452; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4454 = 7'h54 == index ? ram_1_84 : _GEN_4453; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4455 = 7'h55 == index ? ram_1_85 : _GEN_4454; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4456 = 7'h56 == index ? ram_1_86 : _GEN_4455; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4457 = 7'h57 == index ? ram_1_87 : _GEN_4456; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4458 = 7'h58 == index ? ram_1_88 : _GEN_4457; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4459 = 7'h59 == index ? ram_1_89 : _GEN_4458; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4460 = 7'h5a == index ? ram_1_90 : _GEN_4459; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4461 = 7'h5b == index ? ram_1_91 : _GEN_4460; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4462 = 7'h5c == index ? ram_1_92 : _GEN_4461; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4463 = 7'h5d == index ? ram_1_93 : _GEN_4462; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4464 = 7'h5e == index ? ram_1_94 : _GEN_4463; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4465 = 7'h5f == index ? ram_1_95 : _GEN_4464; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4466 = 7'h60 == index ? ram_1_96 : _GEN_4465; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4467 = 7'h61 == index ? ram_1_97 : _GEN_4466; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4468 = 7'h62 == index ? ram_1_98 : _GEN_4467; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4469 = 7'h63 == index ? ram_1_99 : _GEN_4468; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4470 = 7'h64 == index ? ram_1_100 : _GEN_4469; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4471 = 7'h65 == index ? ram_1_101 : _GEN_4470; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4472 = 7'h66 == index ? ram_1_102 : _GEN_4471; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4473 = 7'h67 == index ? ram_1_103 : _GEN_4472; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4474 = 7'h68 == index ? ram_1_104 : _GEN_4473; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4475 = 7'h69 == index ? ram_1_105 : _GEN_4474; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4476 = 7'h6a == index ? ram_1_106 : _GEN_4475; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4477 = 7'h6b == index ? ram_1_107 : _GEN_4476; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4478 = 7'h6c == index ? ram_1_108 : _GEN_4477; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4479 = 7'h6d == index ? ram_1_109 : _GEN_4478; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4480 = 7'h6e == index ? ram_1_110 : _GEN_4479; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4481 = 7'h6f == index ? ram_1_111 : _GEN_4480; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4482 = 7'h70 == index ? ram_1_112 : _GEN_4481; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4483 = 7'h71 == index ? ram_1_113 : _GEN_4482; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4484 = 7'h72 == index ? ram_1_114 : _GEN_4483; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4485 = 7'h73 == index ? ram_1_115 : _GEN_4484; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4486 = 7'h74 == index ? ram_1_116 : _GEN_4485; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4487 = 7'h75 == index ? ram_1_117 : _GEN_4486; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4488 = 7'h76 == index ? ram_1_118 : _GEN_4487; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4489 = 7'h77 == index ? ram_1_119 : _GEN_4488; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4490 = 7'h78 == index ? ram_1_120 : _GEN_4489; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4491 = 7'h79 == index ? ram_1_121 : _GEN_4490; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4492 = 7'h7a == index ? ram_1_122 : _GEN_4491; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4493 = 7'h7b == index ? ram_1_123 : _GEN_4492; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4494 = 7'h7c == index ? ram_1_124 : _GEN_4493; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4495 = 7'h7d == index ? ram_1_125 : _GEN_4494; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4496 = 7'h7e == index ? ram_1_126 : _GEN_4495; // @[d_cache.scala 152:{41,41}]
  wire [63:0] _GEN_4497 = 7'h7f == index ? ram_1_127 : _GEN_4496; // @[d_cache.scala 152:{41,41}]
  wire [38:0] _write_back_addr_T_2 = {_GEN_384, 7'h0}; // @[d_cache.scala 153:57]
  wire [38:0] _write_back_addr_T_3 = _write_back_addr_T_2 | _GEN_15779; // @[d_cache.scala 153:62]
  wire  _GEN_4754 = 7'h0 == index ? 1'h0 : dirty_1_0; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4755 = 7'h1 == index ? 1'h0 : dirty_1_1; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4756 = 7'h2 == index ? 1'h0 : dirty_1_2; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4757 = 7'h3 == index ? 1'h0 : dirty_1_3; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4758 = 7'h4 == index ? 1'h0 : dirty_1_4; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4759 = 7'h5 == index ? 1'h0 : dirty_1_5; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4760 = 7'h6 == index ? 1'h0 : dirty_1_6; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4761 = 7'h7 == index ? 1'h0 : dirty_1_7; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4762 = 7'h8 == index ? 1'h0 : dirty_1_8; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4763 = 7'h9 == index ? 1'h0 : dirty_1_9; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4764 = 7'ha == index ? 1'h0 : dirty_1_10; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4765 = 7'hb == index ? 1'h0 : dirty_1_11; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4766 = 7'hc == index ? 1'h0 : dirty_1_12; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4767 = 7'hd == index ? 1'h0 : dirty_1_13; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4768 = 7'he == index ? 1'h0 : dirty_1_14; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4769 = 7'hf == index ? 1'h0 : dirty_1_15; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4770 = 7'h10 == index ? 1'h0 : dirty_1_16; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4771 = 7'h11 == index ? 1'h0 : dirty_1_17; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4772 = 7'h12 == index ? 1'h0 : dirty_1_18; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4773 = 7'h13 == index ? 1'h0 : dirty_1_19; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4774 = 7'h14 == index ? 1'h0 : dirty_1_20; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4775 = 7'h15 == index ? 1'h0 : dirty_1_21; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4776 = 7'h16 == index ? 1'h0 : dirty_1_22; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4777 = 7'h17 == index ? 1'h0 : dirty_1_23; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4778 = 7'h18 == index ? 1'h0 : dirty_1_24; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4779 = 7'h19 == index ? 1'h0 : dirty_1_25; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4780 = 7'h1a == index ? 1'h0 : dirty_1_26; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4781 = 7'h1b == index ? 1'h0 : dirty_1_27; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4782 = 7'h1c == index ? 1'h0 : dirty_1_28; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4783 = 7'h1d == index ? 1'h0 : dirty_1_29; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4784 = 7'h1e == index ? 1'h0 : dirty_1_30; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4785 = 7'h1f == index ? 1'h0 : dirty_1_31; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4786 = 7'h20 == index ? 1'h0 : dirty_1_32; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4787 = 7'h21 == index ? 1'h0 : dirty_1_33; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4788 = 7'h22 == index ? 1'h0 : dirty_1_34; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4789 = 7'h23 == index ? 1'h0 : dirty_1_35; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4790 = 7'h24 == index ? 1'h0 : dirty_1_36; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4791 = 7'h25 == index ? 1'h0 : dirty_1_37; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4792 = 7'h26 == index ? 1'h0 : dirty_1_38; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4793 = 7'h27 == index ? 1'h0 : dirty_1_39; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4794 = 7'h28 == index ? 1'h0 : dirty_1_40; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4795 = 7'h29 == index ? 1'h0 : dirty_1_41; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4796 = 7'h2a == index ? 1'h0 : dirty_1_42; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4797 = 7'h2b == index ? 1'h0 : dirty_1_43; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4798 = 7'h2c == index ? 1'h0 : dirty_1_44; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4799 = 7'h2d == index ? 1'h0 : dirty_1_45; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4800 = 7'h2e == index ? 1'h0 : dirty_1_46; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4801 = 7'h2f == index ? 1'h0 : dirty_1_47; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4802 = 7'h30 == index ? 1'h0 : dirty_1_48; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4803 = 7'h31 == index ? 1'h0 : dirty_1_49; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4804 = 7'h32 == index ? 1'h0 : dirty_1_50; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4805 = 7'h33 == index ? 1'h0 : dirty_1_51; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4806 = 7'h34 == index ? 1'h0 : dirty_1_52; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4807 = 7'h35 == index ? 1'h0 : dirty_1_53; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4808 = 7'h36 == index ? 1'h0 : dirty_1_54; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4809 = 7'h37 == index ? 1'h0 : dirty_1_55; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4810 = 7'h38 == index ? 1'h0 : dirty_1_56; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4811 = 7'h39 == index ? 1'h0 : dirty_1_57; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4812 = 7'h3a == index ? 1'h0 : dirty_1_58; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4813 = 7'h3b == index ? 1'h0 : dirty_1_59; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4814 = 7'h3c == index ? 1'h0 : dirty_1_60; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4815 = 7'h3d == index ? 1'h0 : dirty_1_61; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4816 = 7'h3e == index ? 1'h0 : dirty_1_62; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4817 = 7'h3f == index ? 1'h0 : dirty_1_63; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4818 = 7'h40 == index ? 1'h0 : dirty_1_64; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4819 = 7'h41 == index ? 1'h0 : dirty_1_65; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4820 = 7'h42 == index ? 1'h0 : dirty_1_66; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4821 = 7'h43 == index ? 1'h0 : dirty_1_67; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4822 = 7'h44 == index ? 1'h0 : dirty_1_68; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4823 = 7'h45 == index ? 1'h0 : dirty_1_69; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4824 = 7'h46 == index ? 1'h0 : dirty_1_70; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4825 = 7'h47 == index ? 1'h0 : dirty_1_71; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4826 = 7'h48 == index ? 1'h0 : dirty_1_72; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4827 = 7'h49 == index ? 1'h0 : dirty_1_73; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4828 = 7'h4a == index ? 1'h0 : dirty_1_74; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4829 = 7'h4b == index ? 1'h0 : dirty_1_75; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4830 = 7'h4c == index ? 1'h0 : dirty_1_76; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4831 = 7'h4d == index ? 1'h0 : dirty_1_77; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4832 = 7'h4e == index ? 1'h0 : dirty_1_78; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4833 = 7'h4f == index ? 1'h0 : dirty_1_79; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4834 = 7'h50 == index ? 1'h0 : dirty_1_80; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4835 = 7'h51 == index ? 1'h0 : dirty_1_81; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4836 = 7'h52 == index ? 1'h0 : dirty_1_82; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4837 = 7'h53 == index ? 1'h0 : dirty_1_83; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4838 = 7'h54 == index ? 1'h0 : dirty_1_84; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4839 = 7'h55 == index ? 1'h0 : dirty_1_85; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4840 = 7'h56 == index ? 1'h0 : dirty_1_86; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4841 = 7'h57 == index ? 1'h0 : dirty_1_87; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4842 = 7'h58 == index ? 1'h0 : dirty_1_88; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4843 = 7'h59 == index ? 1'h0 : dirty_1_89; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4844 = 7'h5a == index ? 1'h0 : dirty_1_90; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4845 = 7'h5b == index ? 1'h0 : dirty_1_91; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4846 = 7'h5c == index ? 1'h0 : dirty_1_92; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4847 = 7'h5d == index ? 1'h0 : dirty_1_93; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4848 = 7'h5e == index ? 1'h0 : dirty_1_94; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4849 = 7'h5f == index ? 1'h0 : dirty_1_95; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4850 = 7'h60 == index ? 1'h0 : dirty_1_96; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4851 = 7'h61 == index ? 1'h0 : dirty_1_97; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4852 = 7'h62 == index ? 1'h0 : dirty_1_98; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4853 = 7'h63 == index ? 1'h0 : dirty_1_99; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4854 = 7'h64 == index ? 1'h0 : dirty_1_100; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4855 = 7'h65 == index ? 1'h0 : dirty_1_101; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4856 = 7'h66 == index ? 1'h0 : dirty_1_102; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4857 = 7'h67 == index ? 1'h0 : dirty_1_103; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4858 = 7'h68 == index ? 1'h0 : dirty_1_104; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4859 = 7'h69 == index ? 1'h0 : dirty_1_105; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4860 = 7'h6a == index ? 1'h0 : dirty_1_106; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4861 = 7'h6b == index ? 1'h0 : dirty_1_107; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4862 = 7'h6c == index ? 1'h0 : dirty_1_108; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4863 = 7'h6d == index ? 1'h0 : dirty_1_109; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4864 = 7'h6e == index ? 1'h0 : dirty_1_110; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4865 = 7'h6f == index ? 1'h0 : dirty_1_111; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4866 = 7'h70 == index ? 1'h0 : dirty_1_112; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4867 = 7'h71 == index ? 1'h0 : dirty_1_113; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4868 = 7'h72 == index ? 1'h0 : dirty_1_114; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4869 = 7'h73 == index ? 1'h0 : dirty_1_115; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4870 = 7'h74 == index ? 1'h0 : dirty_1_116; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4871 = 7'h75 == index ? 1'h0 : dirty_1_117; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4872 = 7'h76 == index ? 1'h0 : dirty_1_118; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4873 = 7'h77 == index ? 1'h0 : dirty_1_119; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4874 = 7'h78 == index ? 1'h0 : dirty_1_120; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4875 = 7'h79 == index ? 1'h0 : dirty_1_121; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4876 = 7'h7a == index ? 1'h0 : dirty_1_122; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4877 = 7'h7b == index ? 1'h0 : dirty_1_123; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4878 = 7'h7c == index ? 1'h0 : dirty_1_124; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4879 = 7'h7d == index ? 1'h0 : dirty_1_125; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4880 = 7'h7e == index ? 1'h0 : dirty_1_126; // @[d_cache.scala 156:{40,40} 25:26]
  wire  _GEN_4881 = 7'h7f == index ? 1'h0 : dirty_1_127; // @[d_cache.scala 156:{40,40} 25:26]
  wire [63:0] _GEN_5394 = _GEN_774 ? _GEN_4497 : write_back_data; // @[d_cache.scala 151:47 152:41 29:34]
  wire [38:0] _GEN_5395 = _GEN_774 ? _write_back_addr_T_3 : {{7'd0}, write_back_addr}; // @[d_cache.scala 151:47 153:41 30:34]
  wire [63:0] _GEN_5396 = _GEN_774 ? _GEN_2446 : _GEN_2446; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5397 = _GEN_774 ? _GEN_2447 : _GEN_2447; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5398 = _GEN_774 ? _GEN_2448 : _GEN_2448; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5399 = _GEN_774 ? _GEN_2449 : _GEN_2449; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5400 = _GEN_774 ? _GEN_2450 : _GEN_2450; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5401 = _GEN_774 ? _GEN_2451 : _GEN_2451; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5402 = _GEN_774 ? _GEN_2452 : _GEN_2452; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5403 = _GEN_774 ? _GEN_2453 : _GEN_2453; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5404 = _GEN_774 ? _GEN_2454 : _GEN_2454; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5405 = _GEN_774 ? _GEN_2455 : _GEN_2455; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5406 = _GEN_774 ? _GEN_2456 : _GEN_2456; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5407 = _GEN_774 ? _GEN_2457 : _GEN_2457; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5408 = _GEN_774 ? _GEN_2458 : _GEN_2458; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5409 = _GEN_774 ? _GEN_2459 : _GEN_2459; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5410 = _GEN_774 ? _GEN_2460 : _GEN_2460; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5411 = _GEN_774 ? _GEN_2461 : _GEN_2461; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5412 = _GEN_774 ? _GEN_2462 : _GEN_2462; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5413 = _GEN_774 ? _GEN_2463 : _GEN_2463; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5414 = _GEN_774 ? _GEN_2464 : _GEN_2464; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5415 = _GEN_774 ? _GEN_2465 : _GEN_2465; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5416 = _GEN_774 ? _GEN_2466 : _GEN_2466; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5417 = _GEN_774 ? _GEN_2467 : _GEN_2467; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5418 = _GEN_774 ? _GEN_2468 : _GEN_2468; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5419 = _GEN_774 ? _GEN_2469 : _GEN_2469; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5420 = _GEN_774 ? _GEN_2470 : _GEN_2470; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5421 = _GEN_774 ? _GEN_2471 : _GEN_2471; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5422 = _GEN_774 ? _GEN_2472 : _GEN_2472; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5423 = _GEN_774 ? _GEN_2473 : _GEN_2473; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5424 = _GEN_774 ? _GEN_2474 : _GEN_2474; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5425 = _GEN_774 ? _GEN_2475 : _GEN_2475; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5426 = _GEN_774 ? _GEN_2476 : _GEN_2476; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5427 = _GEN_774 ? _GEN_2477 : _GEN_2477; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5428 = _GEN_774 ? _GEN_2478 : _GEN_2478; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5429 = _GEN_774 ? _GEN_2479 : _GEN_2479; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5430 = _GEN_774 ? _GEN_2480 : _GEN_2480; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5431 = _GEN_774 ? _GEN_2481 : _GEN_2481; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5432 = _GEN_774 ? _GEN_2482 : _GEN_2482; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5433 = _GEN_774 ? _GEN_2483 : _GEN_2483; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5434 = _GEN_774 ? _GEN_2484 : _GEN_2484; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5435 = _GEN_774 ? _GEN_2485 : _GEN_2485; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5436 = _GEN_774 ? _GEN_2486 : _GEN_2486; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5437 = _GEN_774 ? _GEN_2487 : _GEN_2487; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5438 = _GEN_774 ? _GEN_2488 : _GEN_2488; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5439 = _GEN_774 ? _GEN_2489 : _GEN_2489; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5440 = _GEN_774 ? _GEN_2490 : _GEN_2490; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5441 = _GEN_774 ? _GEN_2491 : _GEN_2491; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5442 = _GEN_774 ? _GEN_2492 : _GEN_2492; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5443 = _GEN_774 ? _GEN_2493 : _GEN_2493; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5444 = _GEN_774 ? _GEN_2494 : _GEN_2494; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5445 = _GEN_774 ? _GEN_2495 : _GEN_2495; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5446 = _GEN_774 ? _GEN_2496 : _GEN_2496; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5447 = _GEN_774 ? _GEN_2497 : _GEN_2497; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5448 = _GEN_774 ? _GEN_2498 : _GEN_2498; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5449 = _GEN_774 ? _GEN_2499 : _GEN_2499; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5450 = _GEN_774 ? _GEN_2500 : _GEN_2500; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5451 = _GEN_774 ? _GEN_2501 : _GEN_2501; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5452 = _GEN_774 ? _GEN_2502 : _GEN_2502; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5453 = _GEN_774 ? _GEN_2503 : _GEN_2503; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5454 = _GEN_774 ? _GEN_2504 : _GEN_2504; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5455 = _GEN_774 ? _GEN_2505 : _GEN_2505; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5456 = _GEN_774 ? _GEN_2506 : _GEN_2506; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5457 = _GEN_774 ? _GEN_2507 : _GEN_2507; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5458 = _GEN_774 ? _GEN_2508 : _GEN_2508; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5459 = _GEN_774 ? _GEN_2509 : _GEN_2509; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5460 = _GEN_774 ? _GEN_2510 : _GEN_2510; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5461 = _GEN_774 ? _GEN_2511 : _GEN_2511; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5462 = _GEN_774 ? _GEN_2512 : _GEN_2512; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5463 = _GEN_774 ? _GEN_2513 : _GEN_2513; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5464 = _GEN_774 ? _GEN_2514 : _GEN_2514; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5465 = _GEN_774 ? _GEN_2515 : _GEN_2515; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5466 = _GEN_774 ? _GEN_2516 : _GEN_2516; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5467 = _GEN_774 ? _GEN_2517 : _GEN_2517; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5468 = _GEN_774 ? _GEN_2518 : _GEN_2518; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5469 = _GEN_774 ? _GEN_2519 : _GEN_2519; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5470 = _GEN_774 ? _GEN_2520 : _GEN_2520; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5471 = _GEN_774 ? _GEN_2521 : _GEN_2521; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5472 = _GEN_774 ? _GEN_2522 : _GEN_2522; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5473 = _GEN_774 ? _GEN_2523 : _GEN_2523; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5474 = _GEN_774 ? _GEN_2524 : _GEN_2524; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5475 = _GEN_774 ? _GEN_2525 : _GEN_2525; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5476 = _GEN_774 ? _GEN_2526 : _GEN_2526; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5477 = _GEN_774 ? _GEN_2527 : _GEN_2527; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5478 = _GEN_774 ? _GEN_2528 : _GEN_2528; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5479 = _GEN_774 ? _GEN_2529 : _GEN_2529; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5480 = _GEN_774 ? _GEN_2530 : _GEN_2530; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5481 = _GEN_774 ? _GEN_2531 : _GEN_2531; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5482 = _GEN_774 ? _GEN_2532 : _GEN_2532; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5483 = _GEN_774 ? _GEN_2533 : _GEN_2533; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5484 = _GEN_774 ? _GEN_2534 : _GEN_2534; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5485 = _GEN_774 ? _GEN_2535 : _GEN_2535; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5486 = _GEN_774 ? _GEN_2536 : _GEN_2536; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5487 = _GEN_774 ? _GEN_2537 : _GEN_2537; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5488 = _GEN_774 ? _GEN_2538 : _GEN_2538; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5489 = _GEN_774 ? _GEN_2539 : _GEN_2539; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5490 = _GEN_774 ? _GEN_2540 : _GEN_2540; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5491 = _GEN_774 ? _GEN_2541 : _GEN_2541; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5492 = _GEN_774 ? _GEN_2542 : _GEN_2542; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5493 = _GEN_774 ? _GEN_2543 : _GEN_2543; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5494 = _GEN_774 ? _GEN_2544 : _GEN_2544; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5495 = _GEN_774 ? _GEN_2545 : _GEN_2545; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5496 = _GEN_774 ? _GEN_2546 : _GEN_2546; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5497 = _GEN_774 ? _GEN_2547 : _GEN_2547; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5498 = _GEN_774 ? _GEN_2548 : _GEN_2548; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5499 = _GEN_774 ? _GEN_2549 : _GEN_2549; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5500 = _GEN_774 ? _GEN_2550 : _GEN_2550; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5501 = _GEN_774 ? _GEN_2551 : _GEN_2551; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5502 = _GEN_774 ? _GEN_2552 : _GEN_2552; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5503 = _GEN_774 ? _GEN_2553 : _GEN_2553; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5504 = _GEN_774 ? _GEN_2554 : _GEN_2554; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5505 = _GEN_774 ? _GEN_2555 : _GEN_2555; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5506 = _GEN_774 ? _GEN_2556 : _GEN_2556; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5507 = _GEN_774 ? _GEN_2557 : _GEN_2557; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5508 = _GEN_774 ? _GEN_2558 : _GEN_2558; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5509 = _GEN_774 ? _GEN_2559 : _GEN_2559; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5510 = _GEN_774 ? _GEN_2560 : _GEN_2560; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5511 = _GEN_774 ? _GEN_2561 : _GEN_2561; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5512 = _GEN_774 ? _GEN_2562 : _GEN_2562; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5513 = _GEN_774 ? _GEN_2563 : _GEN_2563; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5514 = _GEN_774 ? _GEN_2564 : _GEN_2564; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5515 = _GEN_774 ? _GEN_2565 : _GEN_2565; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5516 = _GEN_774 ? _GEN_2566 : _GEN_2566; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5517 = _GEN_774 ? _GEN_2567 : _GEN_2567; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5518 = _GEN_774 ? _GEN_2568 : _GEN_2568; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5519 = _GEN_774 ? _GEN_2569 : _GEN_2569; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5520 = _GEN_774 ? _GEN_2570 : _GEN_2570; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5521 = _GEN_774 ? _GEN_2571 : _GEN_2571; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5522 = _GEN_774 ? _GEN_2572 : _GEN_2572; // @[d_cache.scala 151:47]
  wire [63:0] _GEN_5523 = _GEN_774 ? _GEN_2573 : _GEN_2573; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5524 = _GEN_774 ? _GEN_2574 : _GEN_2574; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5525 = _GEN_774 ? _GEN_2575 : _GEN_2575; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5526 = _GEN_774 ? _GEN_2576 : _GEN_2576; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5527 = _GEN_774 ? _GEN_2577 : _GEN_2577; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5528 = _GEN_774 ? _GEN_2578 : _GEN_2578; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5529 = _GEN_774 ? _GEN_2579 : _GEN_2579; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5530 = _GEN_774 ? _GEN_2580 : _GEN_2580; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5531 = _GEN_774 ? _GEN_2581 : _GEN_2581; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5532 = _GEN_774 ? _GEN_2582 : _GEN_2582; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5533 = _GEN_774 ? _GEN_2583 : _GEN_2583; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5534 = _GEN_774 ? _GEN_2584 : _GEN_2584; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5535 = _GEN_774 ? _GEN_2585 : _GEN_2585; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5536 = _GEN_774 ? _GEN_2586 : _GEN_2586; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5537 = _GEN_774 ? _GEN_2587 : _GEN_2587; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5538 = _GEN_774 ? _GEN_2588 : _GEN_2588; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5539 = _GEN_774 ? _GEN_2589 : _GEN_2589; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5540 = _GEN_774 ? _GEN_2590 : _GEN_2590; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5541 = _GEN_774 ? _GEN_2591 : _GEN_2591; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5542 = _GEN_774 ? _GEN_2592 : _GEN_2592; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5543 = _GEN_774 ? _GEN_2593 : _GEN_2593; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5544 = _GEN_774 ? _GEN_2594 : _GEN_2594; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5545 = _GEN_774 ? _GEN_2595 : _GEN_2595; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5546 = _GEN_774 ? _GEN_2596 : _GEN_2596; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5547 = _GEN_774 ? _GEN_2597 : _GEN_2597; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5548 = _GEN_774 ? _GEN_2598 : _GEN_2598; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5549 = _GEN_774 ? _GEN_2599 : _GEN_2599; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5550 = _GEN_774 ? _GEN_2600 : _GEN_2600; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5551 = _GEN_774 ? _GEN_2601 : _GEN_2601; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5552 = _GEN_774 ? _GEN_2602 : _GEN_2602; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5553 = _GEN_774 ? _GEN_2603 : _GEN_2603; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5554 = _GEN_774 ? _GEN_2604 : _GEN_2604; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5555 = _GEN_774 ? _GEN_2605 : _GEN_2605; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5556 = _GEN_774 ? _GEN_2606 : _GEN_2606; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5557 = _GEN_774 ? _GEN_2607 : _GEN_2607; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5558 = _GEN_774 ? _GEN_2608 : _GEN_2608; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5559 = _GEN_774 ? _GEN_2609 : _GEN_2609; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5560 = _GEN_774 ? _GEN_2610 : _GEN_2610; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5561 = _GEN_774 ? _GEN_2611 : _GEN_2611; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5562 = _GEN_774 ? _GEN_2612 : _GEN_2612; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5563 = _GEN_774 ? _GEN_2613 : _GEN_2613; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5564 = _GEN_774 ? _GEN_2614 : _GEN_2614; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5565 = _GEN_774 ? _GEN_2615 : _GEN_2615; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5566 = _GEN_774 ? _GEN_2616 : _GEN_2616; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5567 = _GEN_774 ? _GEN_2617 : _GEN_2617; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5568 = _GEN_774 ? _GEN_2618 : _GEN_2618; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5569 = _GEN_774 ? _GEN_2619 : _GEN_2619; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5570 = _GEN_774 ? _GEN_2620 : _GEN_2620; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5571 = _GEN_774 ? _GEN_2621 : _GEN_2621; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5572 = _GEN_774 ? _GEN_2622 : _GEN_2622; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5573 = _GEN_774 ? _GEN_2623 : _GEN_2623; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5574 = _GEN_774 ? _GEN_2624 : _GEN_2624; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5575 = _GEN_774 ? _GEN_2625 : _GEN_2625; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5576 = _GEN_774 ? _GEN_2626 : _GEN_2626; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5577 = _GEN_774 ? _GEN_2627 : _GEN_2627; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5578 = _GEN_774 ? _GEN_2628 : _GEN_2628; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5579 = _GEN_774 ? _GEN_2629 : _GEN_2629; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5580 = _GEN_774 ? _GEN_2630 : _GEN_2630; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5581 = _GEN_774 ? _GEN_2631 : _GEN_2631; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5582 = _GEN_774 ? _GEN_2632 : _GEN_2632; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5583 = _GEN_774 ? _GEN_2633 : _GEN_2633; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5584 = _GEN_774 ? _GEN_2634 : _GEN_2634; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5585 = _GEN_774 ? _GEN_2635 : _GEN_2635; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5586 = _GEN_774 ? _GEN_2636 : _GEN_2636; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5587 = _GEN_774 ? _GEN_2637 : _GEN_2637; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5588 = _GEN_774 ? _GEN_2638 : _GEN_2638; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5589 = _GEN_774 ? _GEN_2639 : _GEN_2639; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5590 = _GEN_774 ? _GEN_2640 : _GEN_2640; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5591 = _GEN_774 ? _GEN_2641 : _GEN_2641; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5592 = _GEN_774 ? _GEN_2642 : _GEN_2642; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5593 = _GEN_774 ? _GEN_2643 : _GEN_2643; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5594 = _GEN_774 ? _GEN_2644 : _GEN_2644; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5595 = _GEN_774 ? _GEN_2645 : _GEN_2645; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5596 = _GEN_774 ? _GEN_2646 : _GEN_2646; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5597 = _GEN_774 ? _GEN_2647 : _GEN_2647; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5598 = _GEN_774 ? _GEN_2648 : _GEN_2648; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5599 = _GEN_774 ? _GEN_2649 : _GEN_2649; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5600 = _GEN_774 ? _GEN_2650 : _GEN_2650; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5601 = _GEN_774 ? _GEN_2651 : _GEN_2651; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5602 = _GEN_774 ? _GEN_2652 : _GEN_2652; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5603 = _GEN_774 ? _GEN_2653 : _GEN_2653; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5604 = _GEN_774 ? _GEN_2654 : _GEN_2654; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5605 = _GEN_774 ? _GEN_2655 : _GEN_2655; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5606 = _GEN_774 ? _GEN_2656 : _GEN_2656; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5607 = _GEN_774 ? _GEN_2657 : _GEN_2657; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5608 = _GEN_774 ? _GEN_2658 : _GEN_2658; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5609 = _GEN_774 ? _GEN_2659 : _GEN_2659; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5610 = _GEN_774 ? _GEN_2660 : _GEN_2660; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5611 = _GEN_774 ? _GEN_2661 : _GEN_2661; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5612 = _GEN_774 ? _GEN_2662 : _GEN_2662; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5613 = _GEN_774 ? _GEN_2663 : _GEN_2663; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5614 = _GEN_774 ? _GEN_2664 : _GEN_2664; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5615 = _GEN_774 ? _GEN_2665 : _GEN_2665; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5616 = _GEN_774 ? _GEN_2666 : _GEN_2666; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5617 = _GEN_774 ? _GEN_2667 : _GEN_2667; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5618 = _GEN_774 ? _GEN_2668 : _GEN_2668; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5619 = _GEN_774 ? _GEN_2669 : _GEN_2669; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5620 = _GEN_774 ? _GEN_2670 : _GEN_2670; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5621 = _GEN_774 ? _GEN_2671 : _GEN_2671; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5622 = _GEN_774 ? _GEN_2672 : _GEN_2672; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5623 = _GEN_774 ? _GEN_2673 : _GEN_2673; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5624 = _GEN_774 ? _GEN_2674 : _GEN_2674; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5625 = _GEN_774 ? _GEN_2675 : _GEN_2675; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5626 = _GEN_774 ? _GEN_2676 : _GEN_2676; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5627 = _GEN_774 ? _GEN_2677 : _GEN_2677; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5628 = _GEN_774 ? _GEN_2678 : _GEN_2678; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5629 = _GEN_774 ? _GEN_2679 : _GEN_2679; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5630 = _GEN_774 ? _GEN_2680 : _GEN_2680; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5631 = _GEN_774 ? _GEN_2681 : _GEN_2681; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5632 = _GEN_774 ? _GEN_2682 : _GEN_2682; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5633 = _GEN_774 ? _GEN_2683 : _GEN_2683; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5634 = _GEN_774 ? _GEN_2684 : _GEN_2684; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5635 = _GEN_774 ? _GEN_2685 : _GEN_2685; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5636 = _GEN_774 ? _GEN_2686 : _GEN_2686; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5637 = _GEN_774 ? _GEN_2687 : _GEN_2687; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5638 = _GEN_774 ? _GEN_2688 : _GEN_2688; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5639 = _GEN_774 ? _GEN_2689 : _GEN_2689; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5640 = _GEN_774 ? _GEN_2690 : _GEN_2690; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5641 = _GEN_774 ? _GEN_2691 : _GEN_2691; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5642 = _GEN_774 ? _GEN_2692 : _GEN_2692; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5643 = _GEN_774 ? _GEN_2693 : _GEN_2693; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5644 = _GEN_774 ? _GEN_2694 : _GEN_2694; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5645 = _GEN_774 ? _GEN_2695 : _GEN_2695; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5646 = _GEN_774 ? _GEN_2696 : _GEN_2696; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5647 = _GEN_774 ? _GEN_2697 : _GEN_2697; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5648 = _GEN_774 ? _GEN_2698 : _GEN_2698; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5649 = _GEN_774 ? _GEN_2699 : _GEN_2699; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5650 = _GEN_774 ? _GEN_2700 : _GEN_2700; // @[d_cache.scala 151:47]
  wire [31:0] _GEN_5651 = _GEN_774 ? _GEN_2701 : _GEN_2701; // @[d_cache.scala 151:47]
  wire  _GEN_5652 = _GEN_774 ? _GEN_4754 : dirty_1_0; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5653 = _GEN_774 ? _GEN_4755 : dirty_1_1; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5654 = _GEN_774 ? _GEN_4756 : dirty_1_2; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5655 = _GEN_774 ? _GEN_4757 : dirty_1_3; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5656 = _GEN_774 ? _GEN_4758 : dirty_1_4; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5657 = _GEN_774 ? _GEN_4759 : dirty_1_5; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5658 = _GEN_774 ? _GEN_4760 : dirty_1_6; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5659 = _GEN_774 ? _GEN_4761 : dirty_1_7; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5660 = _GEN_774 ? _GEN_4762 : dirty_1_8; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5661 = _GEN_774 ? _GEN_4763 : dirty_1_9; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5662 = _GEN_774 ? _GEN_4764 : dirty_1_10; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5663 = _GEN_774 ? _GEN_4765 : dirty_1_11; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5664 = _GEN_774 ? _GEN_4766 : dirty_1_12; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5665 = _GEN_774 ? _GEN_4767 : dirty_1_13; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5666 = _GEN_774 ? _GEN_4768 : dirty_1_14; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5667 = _GEN_774 ? _GEN_4769 : dirty_1_15; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5668 = _GEN_774 ? _GEN_4770 : dirty_1_16; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5669 = _GEN_774 ? _GEN_4771 : dirty_1_17; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5670 = _GEN_774 ? _GEN_4772 : dirty_1_18; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5671 = _GEN_774 ? _GEN_4773 : dirty_1_19; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5672 = _GEN_774 ? _GEN_4774 : dirty_1_20; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5673 = _GEN_774 ? _GEN_4775 : dirty_1_21; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5674 = _GEN_774 ? _GEN_4776 : dirty_1_22; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5675 = _GEN_774 ? _GEN_4777 : dirty_1_23; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5676 = _GEN_774 ? _GEN_4778 : dirty_1_24; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5677 = _GEN_774 ? _GEN_4779 : dirty_1_25; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5678 = _GEN_774 ? _GEN_4780 : dirty_1_26; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5679 = _GEN_774 ? _GEN_4781 : dirty_1_27; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5680 = _GEN_774 ? _GEN_4782 : dirty_1_28; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5681 = _GEN_774 ? _GEN_4783 : dirty_1_29; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5682 = _GEN_774 ? _GEN_4784 : dirty_1_30; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5683 = _GEN_774 ? _GEN_4785 : dirty_1_31; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5684 = _GEN_774 ? _GEN_4786 : dirty_1_32; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5685 = _GEN_774 ? _GEN_4787 : dirty_1_33; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5686 = _GEN_774 ? _GEN_4788 : dirty_1_34; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5687 = _GEN_774 ? _GEN_4789 : dirty_1_35; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5688 = _GEN_774 ? _GEN_4790 : dirty_1_36; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5689 = _GEN_774 ? _GEN_4791 : dirty_1_37; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5690 = _GEN_774 ? _GEN_4792 : dirty_1_38; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5691 = _GEN_774 ? _GEN_4793 : dirty_1_39; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5692 = _GEN_774 ? _GEN_4794 : dirty_1_40; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5693 = _GEN_774 ? _GEN_4795 : dirty_1_41; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5694 = _GEN_774 ? _GEN_4796 : dirty_1_42; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5695 = _GEN_774 ? _GEN_4797 : dirty_1_43; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5696 = _GEN_774 ? _GEN_4798 : dirty_1_44; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5697 = _GEN_774 ? _GEN_4799 : dirty_1_45; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5698 = _GEN_774 ? _GEN_4800 : dirty_1_46; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5699 = _GEN_774 ? _GEN_4801 : dirty_1_47; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5700 = _GEN_774 ? _GEN_4802 : dirty_1_48; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5701 = _GEN_774 ? _GEN_4803 : dirty_1_49; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5702 = _GEN_774 ? _GEN_4804 : dirty_1_50; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5703 = _GEN_774 ? _GEN_4805 : dirty_1_51; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5704 = _GEN_774 ? _GEN_4806 : dirty_1_52; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5705 = _GEN_774 ? _GEN_4807 : dirty_1_53; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5706 = _GEN_774 ? _GEN_4808 : dirty_1_54; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5707 = _GEN_774 ? _GEN_4809 : dirty_1_55; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5708 = _GEN_774 ? _GEN_4810 : dirty_1_56; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5709 = _GEN_774 ? _GEN_4811 : dirty_1_57; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5710 = _GEN_774 ? _GEN_4812 : dirty_1_58; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5711 = _GEN_774 ? _GEN_4813 : dirty_1_59; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5712 = _GEN_774 ? _GEN_4814 : dirty_1_60; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5713 = _GEN_774 ? _GEN_4815 : dirty_1_61; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5714 = _GEN_774 ? _GEN_4816 : dirty_1_62; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5715 = _GEN_774 ? _GEN_4817 : dirty_1_63; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5716 = _GEN_774 ? _GEN_4818 : dirty_1_64; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5717 = _GEN_774 ? _GEN_4819 : dirty_1_65; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5718 = _GEN_774 ? _GEN_4820 : dirty_1_66; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5719 = _GEN_774 ? _GEN_4821 : dirty_1_67; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5720 = _GEN_774 ? _GEN_4822 : dirty_1_68; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5721 = _GEN_774 ? _GEN_4823 : dirty_1_69; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5722 = _GEN_774 ? _GEN_4824 : dirty_1_70; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5723 = _GEN_774 ? _GEN_4825 : dirty_1_71; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5724 = _GEN_774 ? _GEN_4826 : dirty_1_72; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5725 = _GEN_774 ? _GEN_4827 : dirty_1_73; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5726 = _GEN_774 ? _GEN_4828 : dirty_1_74; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5727 = _GEN_774 ? _GEN_4829 : dirty_1_75; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5728 = _GEN_774 ? _GEN_4830 : dirty_1_76; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5729 = _GEN_774 ? _GEN_4831 : dirty_1_77; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5730 = _GEN_774 ? _GEN_4832 : dirty_1_78; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5731 = _GEN_774 ? _GEN_4833 : dirty_1_79; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5732 = _GEN_774 ? _GEN_4834 : dirty_1_80; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5733 = _GEN_774 ? _GEN_4835 : dirty_1_81; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5734 = _GEN_774 ? _GEN_4836 : dirty_1_82; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5735 = _GEN_774 ? _GEN_4837 : dirty_1_83; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5736 = _GEN_774 ? _GEN_4838 : dirty_1_84; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5737 = _GEN_774 ? _GEN_4839 : dirty_1_85; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5738 = _GEN_774 ? _GEN_4840 : dirty_1_86; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5739 = _GEN_774 ? _GEN_4841 : dirty_1_87; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5740 = _GEN_774 ? _GEN_4842 : dirty_1_88; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5741 = _GEN_774 ? _GEN_4843 : dirty_1_89; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5742 = _GEN_774 ? _GEN_4844 : dirty_1_90; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5743 = _GEN_774 ? _GEN_4845 : dirty_1_91; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5744 = _GEN_774 ? _GEN_4846 : dirty_1_92; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5745 = _GEN_774 ? _GEN_4847 : dirty_1_93; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5746 = _GEN_774 ? _GEN_4848 : dirty_1_94; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5747 = _GEN_774 ? _GEN_4849 : dirty_1_95; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5748 = _GEN_774 ? _GEN_4850 : dirty_1_96; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5749 = _GEN_774 ? _GEN_4851 : dirty_1_97; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5750 = _GEN_774 ? _GEN_4852 : dirty_1_98; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5751 = _GEN_774 ? _GEN_4853 : dirty_1_99; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5752 = _GEN_774 ? _GEN_4854 : dirty_1_100; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5753 = _GEN_774 ? _GEN_4855 : dirty_1_101; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5754 = _GEN_774 ? _GEN_4856 : dirty_1_102; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5755 = _GEN_774 ? _GEN_4857 : dirty_1_103; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5756 = _GEN_774 ? _GEN_4858 : dirty_1_104; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5757 = _GEN_774 ? _GEN_4859 : dirty_1_105; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5758 = _GEN_774 ? _GEN_4860 : dirty_1_106; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5759 = _GEN_774 ? _GEN_4861 : dirty_1_107; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5760 = _GEN_774 ? _GEN_4862 : dirty_1_108; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5761 = _GEN_774 ? _GEN_4863 : dirty_1_109; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5762 = _GEN_774 ? _GEN_4864 : dirty_1_110; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5763 = _GEN_774 ? _GEN_4865 : dirty_1_111; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5764 = _GEN_774 ? _GEN_4866 : dirty_1_112; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5765 = _GEN_774 ? _GEN_4867 : dirty_1_113; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5766 = _GEN_774 ? _GEN_4868 : dirty_1_114; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5767 = _GEN_774 ? _GEN_4869 : dirty_1_115; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5768 = _GEN_774 ? _GEN_4870 : dirty_1_116; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5769 = _GEN_774 ? _GEN_4871 : dirty_1_117; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5770 = _GEN_774 ? _GEN_4872 : dirty_1_118; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5771 = _GEN_774 ? _GEN_4873 : dirty_1_119; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5772 = _GEN_774 ? _GEN_4874 : dirty_1_120; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5773 = _GEN_774 ? _GEN_4875 : dirty_1_121; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5774 = _GEN_774 ? _GEN_4876 : dirty_1_122; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5775 = _GEN_774 ? _GEN_4877 : dirty_1_123; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5776 = _GEN_774 ? _GEN_4878 : dirty_1_124; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5777 = _GEN_774 ? _GEN_4879 : dirty_1_125; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5778 = _GEN_774 ? _GEN_4880 : dirty_1_126; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5779 = _GEN_774 ? _GEN_4881 : dirty_1_127; // @[d_cache.scala 151:47 25:26]
  wire  _GEN_5780 = _GEN_774 ? _GEN_2702 : _GEN_2702; // @[d_cache.scala 151:47]
  wire  _GEN_5781 = _GEN_774 ? _GEN_2703 : _GEN_2703; // @[d_cache.scala 151:47]
  wire  _GEN_5782 = _GEN_774 ? _GEN_2704 : _GEN_2704; // @[d_cache.scala 151:47]
  wire  _GEN_5783 = _GEN_774 ? _GEN_2705 : _GEN_2705; // @[d_cache.scala 151:47]
  wire  _GEN_5784 = _GEN_774 ? _GEN_2706 : _GEN_2706; // @[d_cache.scala 151:47]
  wire  _GEN_5785 = _GEN_774 ? _GEN_2707 : _GEN_2707; // @[d_cache.scala 151:47]
  wire  _GEN_5786 = _GEN_774 ? _GEN_2708 : _GEN_2708; // @[d_cache.scala 151:47]
  wire  _GEN_5787 = _GEN_774 ? _GEN_2709 : _GEN_2709; // @[d_cache.scala 151:47]
  wire  _GEN_5788 = _GEN_774 ? _GEN_2710 : _GEN_2710; // @[d_cache.scala 151:47]
  wire  _GEN_5789 = _GEN_774 ? _GEN_2711 : _GEN_2711; // @[d_cache.scala 151:47]
  wire  _GEN_5790 = _GEN_774 ? _GEN_2712 : _GEN_2712; // @[d_cache.scala 151:47]
  wire  _GEN_5791 = _GEN_774 ? _GEN_2713 : _GEN_2713; // @[d_cache.scala 151:47]
  wire  _GEN_5792 = _GEN_774 ? _GEN_2714 : _GEN_2714; // @[d_cache.scala 151:47]
  wire  _GEN_5793 = _GEN_774 ? _GEN_2715 : _GEN_2715; // @[d_cache.scala 151:47]
  wire  _GEN_5794 = _GEN_774 ? _GEN_2716 : _GEN_2716; // @[d_cache.scala 151:47]
  wire  _GEN_5795 = _GEN_774 ? _GEN_2717 : _GEN_2717; // @[d_cache.scala 151:47]
  wire  _GEN_5796 = _GEN_774 ? _GEN_2718 : _GEN_2718; // @[d_cache.scala 151:47]
  wire  _GEN_5797 = _GEN_774 ? _GEN_2719 : _GEN_2719; // @[d_cache.scala 151:47]
  wire  _GEN_5798 = _GEN_774 ? _GEN_2720 : _GEN_2720; // @[d_cache.scala 151:47]
  wire  _GEN_5799 = _GEN_774 ? _GEN_2721 : _GEN_2721; // @[d_cache.scala 151:47]
  wire  _GEN_5800 = _GEN_774 ? _GEN_2722 : _GEN_2722; // @[d_cache.scala 151:47]
  wire  _GEN_5801 = _GEN_774 ? _GEN_2723 : _GEN_2723; // @[d_cache.scala 151:47]
  wire  _GEN_5802 = _GEN_774 ? _GEN_2724 : _GEN_2724; // @[d_cache.scala 151:47]
  wire  _GEN_5803 = _GEN_774 ? _GEN_2725 : _GEN_2725; // @[d_cache.scala 151:47]
  wire  _GEN_5804 = _GEN_774 ? _GEN_2726 : _GEN_2726; // @[d_cache.scala 151:47]
  wire  _GEN_5805 = _GEN_774 ? _GEN_2727 : _GEN_2727; // @[d_cache.scala 151:47]
  wire  _GEN_5806 = _GEN_774 ? _GEN_2728 : _GEN_2728; // @[d_cache.scala 151:47]
  wire  _GEN_5807 = _GEN_774 ? _GEN_2729 : _GEN_2729; // @[d_cache.scala 151:47]
  wire  _GEN_5808 = _GEN_774 ? _GEN_2730 : _GEN_2730; // @[d_cache.scala 151:47]
  wire  _GEN_5809 = _GEN_774 ? _GEN_2731 : _GEN_2731; // @[d_cache.scala 151:47]
  wire  _GEN_5810 = _GEN_774 ? _GEN_2732 : _GEN_2732; // @[d_cache.scala 151:47]
  wire  _GEN_5811 = _GEN_774 ? _GEN_2733 : _GEN_2733; // @[d_cache.scala 151:47]
  wire  _GEN_5812 = _GEN_774 ? _GEN_2734 : _GEN_2734; // @[d_cache.scala 151:47]
  wire  _GEN_5813 = _GEN_774 ? _GEN_2735 : _GEN_2735; // @[d_cache.scala 151:47]
  wire  _GEN_5814 = _GEN_774 ? _GEN_2736 : _GEN_2736; // @[d_cache.scala 151:47]
  wire  _GEN_5815 = _GEN_774 ? _GEN_2737 : _GEN_2737; // @[d_cache.scala 151:47]
  wire  _GEN_5816 = _GEN_774 ? _GEN_2738 : _GEN_2738; // @[d_cache.scala 151:47]
  wire  _GEN_5817 = _GEN_774 ? _GEN_2739 : _GEN_2739; // @[d_cache.scala 151:47]
  wire  _GEN_5818 = _GEN_774 ? _GEN_2740 : _GEN_2740; // @[d_cache.scala 151:47]
  wire  _GEN_5819 = _GEN_774 ? _GEN_2741 : _GEN_2741; // @[d_cache.scala 151:47]
  wire  _GEN_5820 = _GEN_774 ? _GEN_2742 : _GEN_2742; // @[d_cache.scala 151:47]
  wire  _GEN_5821 = _GEN_774 ? _GEN_2743 : _GEN_2743; // @[d_cache.scala 151:47]
  wire  _GEN_5822 = _GEN_774 ? _GEN_2744 : _GEN_2744; // @[d_cache.scala 151:47]
  wire  _GEN_5823 = _GEN_774 ? _GEN_2745 : _GEN_2745; // @[d_cache.scala 151:47]
  wire  _GEN_5824 = _GEN_774 ? _GEN_2746 : _GEN_2746; // @[d_cache.scala 151:47]
  wire  _GEN_5825 = _GEN_774 ? _GEN_2747 : _GEN_2747; // @[d_cache.scala 151:47]
  wire  _GEN_5826 = _GEN_774 ? _GEN_2748 : _GEN_2748; // @[d_cache.scala 151:47]
  wire  _GEN_5827 = _GEN_774 ? _GEN_2749 : _GEN_2749; // @[d_cache.scala 151:47]
  wire  _GEN_5828 = _GEN_774 ? _GEN_2750 : _GEN_2750; // @[d_cache.scala 151:47]
  wire  _GEN_5829 = _GEN_774 ? _GEN_2751 : _GEN_2751; // @[d_cache.scala 151:47]
  wire  _GEN_5830 = _GEN_774 ? _GEN_2752 : _GEN_2752; // @[d_cache.scala 151:47]
  wire  _GEN_5831 = _GEN_774 ? _GEN_2753 : _GEN_2753; // @[d_cache.scala 151:47]
  wire  _GEN_5832 = _GEN_774 ? _GEN_2754 : _GEN_2754; // @[d_cache.scala 151:47]
  wire  _GEN_5833 = _GEN_774 ? _GEN_2755 : _GEN_2755; // @[d_cache.scala 151:47]
  wire  _GEN_5834 = _GEN_774 ? _GEN_2756 : _GEN_2756; // @[d_cache.scala 151:47]
  wire  _GEN_5835 = _GEN_774 ? _GEN_2757 : _GEN_2757; // @[d_cache.scala 151:47]
  wire  _GEN_5836 = _GEN_774 ? _GEN_2758 : _GEN_2758; // @[d_cache.scala 151:47]
  wire  _GEN_5837 = _GEN_774 ? _GEN_2759 : _GEN_2759; // @[d_cache.scala 151:47]
  wire  _GEN_5838 = _GEN_774 ? _GEN_2760 : _GEN_2760; // @[d_cache.scala 151:47]
  wire  _GEN_5839 = _GEN_774 ? _GEN_2761 : _GEN_2761; // @[d_cache.scala 151:47]
  wire  _GEN_5840 = _GEN_774 ? _GEN_2762 : _GEN_2762; // @[d_cache.scala 151:47]
  wire  _GEN_5841 = _GEN_774 ? _GEN_2763 : _GEN_2763; // @[d_cache.scala 151:47]
  wire  _GEN_5842 = _GEN_774 ? _GEN_2764 : _GEN_2764; // @[d_cache.scala 151:47]
  wire  _GEN_5843 = _GEN_774 ? _GEN_2765 : _GEN_2765; // @[d_cache.scala 151:47]
  wire  _GEN_5844 = _GEN_774 ? _GEN_2766 : _GEN_2766; // @[d_cache.scala 151:47]
  wire  _GEN_5845 = _GEN_774 ? _GEN_2767 : _GEN_2767; // @[d_cache.scala 151:47]
  wire  _GEN_5846 = _GEN_774 ? _GEN_2768 : _GEN_2768; // @[d_cache.scala 151:47]
  wire  _GEN_5847 = _GEN_774 ? _GEN_2769 : _GEN_2769; // @[d_cache.scala 151:47]
  wire  _GEN_5848 = _GEN_774 ? _GEN_2770 : _GEN_2770; // @[d_cache.scala 151:47]
  wire  _GEN_5849 = _GEN_774 ? _GEN_2771 : _GEN_2771; // @[d_cache.scala 151:47]
  wire  _GEN_5850 = _GEN_774 ? _GEN_2772 : _GEN_2772; // @[d_cache.scala 151:47]
  wire  _GEN_5851 = _GEN_774 ? _GEN_2773 : _GEN_2773; // @[d_cache.scala 151:47]
  wire  _GEN_5852 = _GEN_774 ? _GEN_2774 : _GEN_2774; // @[d_cache.scala 151:47]
  wire  _GEN_5853 = _GEN_774 ? _GEN_2775 : _GEN_2775; // @[d_cache.scala 151:47]
  wire  _GEN_5854 = _GEN_774 ? _GEN_2776 : _GEN_2776; // @[d_cache.scala 151:47]
  wire  _GEN_5855 = _GEN_774 ? _GEN_2777 : _GEN_2777; // @[d_cache.scala 151:47]
  wire  _GEN_5856 = _GEN_774 ? _GEN_2778 : _GEN_2778; // @[d_cache.scala 151:47]
  wire  _GEN_5857 = _GEN_774 ? _GEN_2779 : _GEN_2779; // @[d_cache.scala 151:47]
  wire  _GEN_5858 = _GEN_774 ? _GEN_2780 : _GEN_2780; // @[d_cache.scala 151:47]
  wire  _GEN_5859 = _GEN_774 ? _GEN_2781 : _GEN_2781; // @[d_cache.scala 151:47]
  wire  _GEN_5860 = _GEN_774 ? _GEN_2782 : _GEN_2782; // @[d_cache.scala 151:47]
  wire  _GEN_5861 = _GEN_774 ? _GEN_2783 : _GEN_2783; // @[d_cache.scala 151:47]
  wire  _GEN_5862 = _GEN_774 ? _GEN_2784 : _GEN_2784; // @[d_cache.scala 151:47]
  wire  _GEN_5863 = _GEN_774 ? _GEN_2785 : _GEN_2785; // @[d_cache.scala 151:47]
  wire  _GEN_5864 = _GEN_774 ? _GEN_2786 : _GEN_2786; // @[d_cache.scala 151:47]
  wire  _GEN_5865 = _GEN_774 ? _GEN_2787 : _GEN_2787; // @[d_cache.scala 151:47]
  wire  _GEN_5866 = _GEN_774 ? _GEN_2788 : _GEN_2788; // @[d_cache.scala 151:47]
  wire  _GEN_5867 = _GEN_774 ? _GEN_2789 : _GEN_2789; // @[d_cache.scala 151:47]
  wire  _GEN_5868 = _GEN_774 ? _GEN_2790 : _GEN_2790; // @[d_cache.scala 151:47]
  wire  _GEN_5869 = _GEN_774 ? _GEN_2791 : _GEN_2791; // @[d_cache.scala 151:47]
  wire  _GEN_5870 = _GEN_774 ? _GEN_2792 : _GEN_2792; // @[d_cache.scala 151:47]
  wire  _GEN_5871 = _GEN_774 ? _GEN_2793 : _GEN_2793; // @[d_cache.scala 151:47]
  wire  _GEN_5872 = _GEN_774 ? _GEN_2794 : _GEN_2794; // @[d_cache.scala 151:47]
  wire  _GEN_5873 = _GEN_774 ? _GEN_2795 : _GEN_2795; // @[d_cache.scala 151:47]
  wire  _GEN_5874 = _GEN_774 ? _GEN_2796 : _GEN_2796; // @[d_cache.scala 151:47]
  wire  _GEN_5875 = _GEN_774 ? _GEN_2797 : _GEN_2797; // @[d_cache.scala 151:47]
  wire  _GEN_5876 = _GEN_774 ? _GEN_2798 : _GEN_2798; // @[d_cache.scala 151:47]
  wire  _GEN_5877 = _GEN_774 ? _GEN_2799 : _GEN_2799; // @[d_cache.scala 151:47]
  wire  _GEN_5878 = _GEN_774 ? _GEN_2800 : _GEN_2800; // @[d_cache.scala 151:47]
  wire  _GEN_5879 = _GEN_774 ? _GEN_2801 : _GEN_2801; // @[d_cache.scala 151:47]
  wire  _GEN_5880 = _GEN_774 ? _GEN_2802 : _GEN_2802; // @[d_cache.scala 151:47]
  wire  _GEN_5881 = _GEN_774 ? _GEN_2803 : _GEN_2803; // @[d_cache.scala 151:47]
  wire  _GEN_5882 = _GEN_774 ? _GEN_2804 : _GEN_2804; // @[d_cache.scala 151:47]
  wire  _GEN_5883 = _GEN_774 ? _GEN_2805 : _GEN_2805; // @[d_cache.scala 151:47]
  wire  _GEN_5884 = _GEN_774 ? _GEN_2806 : _GEN_2806; // @[d_cache.scala 151:47]
  wire  _GEN_5885 = _GEN_774 ? _GEN_2807 : _GEN_2807; // @[d_cache.scala 151:47]
  wire  _GEN_5886 = _GEN_774 ? _GEN_2808 : _GEN_2808; // @[d_cache.scala 151:47]
  wire  _GEN_5887 = _GEN_774 ? _GEN_2809 : _GEN_2809; // @[d_cache.scala 151:47]
  wire  _GEN_5888 = _GEN_774 ? _GEN_2810 : _GEN_2810; // @[d_cache.scala 151:47]
  wire  _GEN_5889 = _GEN_774 ? _GEN_2811 : _GEN_2811; // @[d_cache.scala 151:47]
  wire  _GEN_5890 = _GEN_774 ? _GEN_2812 : _GEN_2812; // @[d_cache.scala 151:47]
  wire  _GEN_5891 = _GEN_774 ? _GEN_2813 : _GEN_2813; // @[d_cache.scala 151:47]
  wire  _GEN_5892 = _GEN_774 ? _GEN_2814 : _GEN_2814; // @[d_cache.scala 151:47]
  wire  _GEN_5893 = _GEN_774 ? _GEN_2815 : _GEN_2815; // @[d_cache.scala 151:47]
  wire  _GEN_5894 = _GEN_774 ? _GEN_2816 : _GEN_2816; // @[d_cache.scala 151:47]
  wire  _GEN_5895 = _GEN_774 ? _GEN_2817 : _GEN_2817; // @[d_cache.scala 151:47]
  wire  _GEN_5896 = _GEN_774 ? _GEN_2818 : _GEN_2818; // @[d_cache.scala 151:47]
  wire  _GEN_5897 = _GEN_774 ? _GEN_2819 : _GEN_2819; // @[d_cache.scala 151:47]
  wire  _GEN_5898 = _GEN_774 ? _GEN_2820 : _GEN_2820; // @[d_cache.scala 151:47]
  wire  _GEN_5899 = _GEN_774 ? _GEN_2821 : _GEN_2821; // @[d_cache.scala 151:47]
  wire  _GEN_5900 = _GEN_774 ? _GEN_2822 : _GEN_2822; // @[d_cache.scala 151:47]
  wire  _GEN_5901 = _GEN_774 ? _GEN_2823 : _GEN_2823; // @[d_cache.scala 151:47]
  wire  _GEN_5902 = _GEN_774 ? _GEN_2824 : _GEN_2824; // @[d_cache.scala 151:47]
  wire  _GEN_5903 = _GEN_774 ? _GEN_2825 : _GEN_2825; // @[d_cache.scala 151:47]
  wire  _GEN_5904 = _GEN_774 ? _GEN_2826 : _GEN_2826; // @[d_cache.scala 151:47]
  wire  _GEN_5905 = _GEN_774 ? _GEN_2827 : _GEN_2827; // @[d_cache.scala 151:47]
  wire  _GEN_5906 = _GEN_774 ? _GEN_2828 : _GEN_2828; // @[d_cache.scala 151:47]
  wire  _GEN_5907 = _GEN_774 ? _GEN_2829 : _GEN_2829; // @[d_cache.scala 151:47]
  wire [2:0] _GEN_5908 = _GEN_774 ? 3'h6 : 3'h7; // @[d_cache.scala 151:47 158:31 161:31]
  wire [63:0] _GEN_5910 = ~quene ? _GEN_3854 : _GEN_5394; // @[d_cache.scala 132:34]
  wire [38:0] _GEN_5911 = ~quene ? _GEN_3855 : _GEN_5395; // @[d_cache.scala 132:34]
  wire [63:0] _GEN_5912 = ~quene ? _GEN_3856 : ram_0_0; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5913 = ~quene ? _GEN_3857 : ram_0_1; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5914 = ~quene ? _GEN_3858 : ram_0_2; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5915 = ~quene ? _GEN_3859 : ram_0_3; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5916 = ~quene ? _GEN_3860 : ram_0_4; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5917 = ~quene ? _GEN_3861 : ram_0_5; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5918 = ~quene ? _GEN_3862 : ram_0_6; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5919 = ~quene ? _GEN_3863 : ram_0_7; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5920 = ~quene ? _GEN_3864 : ram_0_8; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5921 = ~quene ? _GEN_3865 : ram_0_9; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5922 = ~quene ? _GEN_3866 : ram_0_10; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5923 = ~quene ? _GEN_3867 : ram_0_11; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5924 = ~quene ? _GEN_3868 : ram_0_12; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5925 = ~quene ? _GEN_3869 : ram_0_13; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5926 = ~quene ? _GEN_3870 : ram_0_14; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5927 = ~quene ? _GEN_3871 : ram_0_15; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5928 = ~quene ? _GEN_3872 : ram_0_16; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5929 = ~quene ? _GEN_3873 : ram_0_17; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5930 = ~quene ? _GEN_3874 : ram_0_18; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5931 = ~quene ? _GEN_3875 : ram_0_19; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5932 = ~quene ? _GEN_3876 : ram_0_20; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5933 = ~quene ? _GEN_3877 : ram_0_21; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5934 = ~quene ? _GEN_3878 : ram_0_22; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5935 = ~quene ? _GEN_3879 : ram_0_23; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5936 = ~quene ? _GEN_3880 : ram_0_24; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5937 = ~quene ? _GEN_3881 : ram_0_25; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5938 = ~quene ? _GEN_3882 : ram_0_26; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5939 = ~quene ? _GEN_3883 : ram_0_27; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5940 = ~quene ? _GEN_3884 : ram_0_28; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5941 = ~quene ? _GEN_3885 : ram_0_29; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5942 = ~quene ? _GEN_3886 : ram_0_30; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5943 = ~quene ? _GEN_3887 : ram_0_31; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5944 = ~quene ? _GEN_3888 : ram_0_32; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5945 = ~quene ? _GEN_3889 : ram_0_33; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5946 = ~quene ? _GEN_3890 : ram_0_34; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5947 = ~quene ? _GEN_3891 : ram_0_35; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5948 = ~quene ? _GEN_3892 : ram_0_36; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5949 = ~quene ? _GEN_3893 : ram_0_37; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5950 = ~quene ? _GEN_3894 : ram_0_38; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5951 = ~quene ? _GEN_3895 : ram_0_39; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5952 = ~quene ? _GEN_3896 : ram_0_40; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5953 = ~quene ? _GEN_3897 : ram_0_41; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5954 = ~quene ? _GEN_3898 : ram_0_42; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5955 = ~quene ? _GEN_3899 : ram_0_43; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5956 = ~quene ? _GEN_3900 : ram_0_44; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5957 = ~quene ? _GEN_3901 : ram_0_45; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5958 = ~quene ? _GEN_3902 : ram_0_46; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5959 = ~quene ? _GEN_3903 : ram_0_47; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5960 = ~quene ? _GEN_3904 : ram_0_48; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5961 = ~quene ? _GEN_3905 : ram_0_49; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5962 = ~quene ? _GEN_3906 : ram_0_50; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5963 = ~quene ? _GEN_3907 : ram_0_51; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5964 = ~quene ? _GEN_3908 : ram_0_52; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5965 = ~quene ? _GEN_3909 : ram_0_53; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5966 = ~quene ? _GEN_3910 : ram_0_54; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5967 = ~quene ? _GEN_3911 : ram_0_55; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5968 = ~quene ? _GEN_3912 : ram_0_56; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5969 = ~quene ? _GEN_3913 : ram_0_57; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5970 = ~quene ? _GEN_3914 : ram_0_58; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5971 = ~quene ? _GEN_3915 : ram_0_59; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5972 = ~quene ? _GEN_3916 : ram_0_60; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5973 = ~quene ? _GEN_3917 : ram_0_61; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5974 = ~quene ? _GEN_3918 : ram_0_62; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5975 = ~quene ? _GEN_3919 : ram_0_63; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5976 = ~quene ? _GEN_3920 : ram_0_64; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5977 = ~quene ? _GEN_3921 : ram_0_65; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5978 = ~quene ? _GEN_3922 : ram_0_66; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5979 = ~quene ? _GEN_3923 : ram_0_67; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5980 = ~quene ? _GEN_3924 : ram_0_68; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5981 = ~quene ? _GEN_3925 : ram_0_69; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5982 = ~quene ? _GEN_3926 : ram_0_70; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5983 = ~quene ? _GEN_3927 : ram_0_71; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5984 = ~quene ? _GEN_3928 : ram_0_72; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5985 = ~quene ? _GEN_3929 : ram_0_73; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5986 = ~quene ? _GEN_3930 : ram_0_74; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5987 = ~quene ? _GEN_3931 : ram_0_75; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5988 = ~quene ? _GEN_3932 : ram_0_76; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5989 = ~quene ? _GEN_3933 : ram_0_77; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5990 = ~quene ? _GEN_3934 : ram_0_78; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5991 = ~quene ? _GEN_3935 : ram_0_79; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5992 = ~quene ? _GEN_3936 : ram_0_80; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5993 = ~quene ? _GEN_3937 : ram_0_81; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5994 = ~quene ? _GEN_3938 : ram_0_82; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5995 = ~quene ? _GEN_3939 : ram_0_83; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5996 = ~quene ? _GEN_3940 : ram_0_84; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5997 = ~quene ? _GEN_3941 : ram_0_85; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5998 = ~quene ? _GEN_3942 : ram_0_86; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_5999 = ~quene ? _GEN_3943 : ram_0_87; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6000 = ~quene ? _GEN_3944 : ram_0_88; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6001 = ~quene ? _GEN_3945 : ram_0_89; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6002 = ~quene ? _GEN_3946 : ram_0_90; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6003 = ~quene ? _GEN_3947 : ram_0_91; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6004 = ~quene ? _GEN_3948 : ram_0_92; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6005 = ~quene ? _GEN_3949 : ram_0_93; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6006 = ~quene ? _GEN_3950 : ram_0_94; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6007 = ~quene ? _GEN_3951 : ram_0_95; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6008 = ~quene ? _GEN_3952 : ram_0_96; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6009 = ~quene ? _GEN_3953 : ram_0_97; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6010 = ~quene ? _GEN_3954 : ram_0_98; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6011 = ~quene ? _GEN_3955 : ram_0_99; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6012 = ~quene ? _GEN_3956 : ram_0_100; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6013 = ~quene ? _GEN_3957 : ram_0_101; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6014 = ~quene ? _GEN_3958 : ram_0_102; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6015 = ~quene ? _GEN_3959 : ram_0_103; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6016 = ~quene ? _GEN_3960 : ram_0_104; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6017 = ~quene ? _GEN_3961 : ram_0_105; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6018 = ~quene ? _GEN_3962 : ram_0_106; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6019 = ~quene ? _GEN_3963 : ram_0_107; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6020 = ~quene ? _GEN_3964 : ram_0_108; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6021 = ~quene ? _GEN_3965 : ram_0_109; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6022 = ~quene ? _GEN_3966 : ram_0_110; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6023 = ~quene ? _GEN_3967 : ram_0_111; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6024 = ~quene ? _GEN_3968 : ram_0_112; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6025 = ~quene ? _GEN_3969 : ram_0_113; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6026 = ~quene ? _GEN_3970 : ram_0_114; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6027 = ~quene ? _GEN_3971 : ram_0_115; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6028 = ~quene ? _GEN_3972 : ram_0_116; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6029 = ~quene ? _GEN_3973 : ram_0_117; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6030 = ~quene ? _GEN_3974 : ram_0_118; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6031 = ~quene ? _GEN_3975 : ram_0_119; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6032 = ~quene ? _GEN_3976 : ram_0_120; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6033 = ~quene ? _GEN_3977 : ram_0_121; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6034 = ~quene ? _GEN_3978 : ram_0_122; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6035 = ~quene ? _GEN_3979 : ram_0_123; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6036 = ~quene ? _GEN_3980 : ram_0_124; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6037 = ~quene ? _GEN_3981 : ram_0_125; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6038 = ~quene ? _GEN_3982 : ram_0_126; // @[d_cache.scala 132:34 18:24]
  wire [63:0] _GEN_6039 = ~quene ? _GEN_3983 : ram_0_127; // @[d_cache.scala 132:34 18:24]
  wire [31:0] _GEN_6040 = ~quene ? _GEN_3984 : tag_0_0; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6041 = ~quene ? _GEN_3985 : tag_0_1; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6042 = ~quene ? _GEN_3986 : tag_0_2; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6043 = ~quene ? _GEN_3987 : tag_0_3; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6044 = ~quene ? _GEN_3988 : tag_0_4; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6045 = ~quene ? _GEN_3989 : tag_0_5; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6046 = ~quene ? _GEN_3990 : tag_0_6; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6047 = ~quene ? _GEN_3991 : tag_0_7; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6048 = ~quene ? _GEN_3992 : tag_0_8; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6049 = ~quene ? _GEN_3993 : tag_0_9; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6050 = ~quene ? _GEN_3994 : tag_0_10; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6051 = ~quene ? _GEN_3995 : tag_0_11; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6052 = ~quene ? _GEN_3996 : tag_0_12; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6053 = ~quene ? _GEN_3997 : tag_0_13; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6054 = ~quene ? _GEN_3998 : tag_0_14; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6055 = ~quene ? _GEN_3999 : tag_0_15; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6056 = ~quene ? _GEN_4000 : tag_0_16; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6057 = ~quene ? _GEN_4001 : tag_0_17; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6058 = ~quene ? _GEN_4002 : tag_0_18; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6059 = ~quene ? _GEN_4003 : tag_0_19; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6060 = ~quene ? _GEN_4004 : tag_0_20; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6061 = ~quene ? _GEN_4005 : tag_0_21; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6062 = ~quene ? _GEN_4006 : tag_0_22; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6063 = ~quene ? _GEN_4007 : tag_0_23; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6064 = ~quene ? _GEN_4008 : tag_0_24; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6065 = ~quene ? _GEN_4009 : tag_0_25; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6066 = ~quene ? _GEN_4010 : tag_0_26; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6067 = ~quene ? _GEN_4011 : tag_0_27; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6068 = ~quene ? _GEN_4012 : tag_0_28; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6069 = ~quene ? _GEN_4013 : tag_0_29; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6070 = ~quene ? _GEN_4014 : tag_0_30; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6071 = ~quene ? _GEN_4015 : tag_0_31; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6072 = ~quene ? _GEN_4016 : tag_0_32; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6073 = ~quene ? _GEN_4017 : tag_0_33; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6074 = ~quene ? _GEN_4018 : tag_0_34; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6075 = ~quene ? _GEN_4019 : tag_0_35; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6076 = ~quene ? _GEN_4020 : tag_0_36; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6077 = ~quene ? _GEN_4021 : tag_0_37; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6078 = ~quene ? _GEN_4022 : tag_0_38; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6079 = ~quene ? _GEN_4023 : tag_0_39; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6080 = ~quene ? _GEN_4024 : tag_0_40; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6081 = ~quene ? _GEN_4025 : tag_0_41; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6082 = ~quene ? _GEN_4026 : tag_0_42; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6083 = ~quene ? _GEN_4027 : tag_0_43; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6084 = ~quene ? _GEN_4028 : tag_0_44; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6085 = ~quene ? _GEN_4029 : tag_0_45; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6086 = ~quene ? _GEN_4030 : tag_0_46; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6087 = ~quene ? _GEN_4031 : tag_0_47; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6088 = ~quene ? _GEN_4032 : tag_0_48; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6089 = ~quene ? _GEN_4033 : tag_0_49; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6090 = ~quene ? _GEN_4034 : tag_0_50; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6091 = ~quene ? _GEN_4035 : tag_0_51; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6092 = ~quene ? _GEN_4036 : tag_0_52; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6093 = ~quene ? _GEN_4037 : tag_0_53; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6094 = ~quene ? _GEN_4038 : tag_0_54; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6095 = ~quene ? _GEN_4039 : tag_0_55; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6096 = ~quene ? _GEN_4040 : tag_0_56; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6097 = ~quene ? _GEN_4041 : tag_0_57; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6098 = ~quene ? _GEN_4042 : tag_0_58; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6099 = ~quene ? _GEN_4043 : tag_0_59; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6100 = ~quene ? _GEN_4044 : tag_0_60; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6101 = ~quene ? _GEN_4045 : tag_0_61; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6102 = ~quene ? _GEN_4046 : tag_0_62; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6103 = ~quene ? _GEN_4047 : tag_0_63; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6104 = ~quene ? _GEN_4048 : tag_0_64; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6105 = ~quene ? _GEN_4049 : tag_0_65; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6106 = ~quene ? _GEN_4050 : tag_0_66; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6107 = ~quene ? _GEN_4051 : tag_0_67; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6108 = ~quene ? _GEN_4052 : tag_0_68; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6109 = ~quene ? _GEN_4053 : tag_0_69; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6110 = ~quene ? _GEN_4054 : tag_0_70; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6111 = ~quene ? _GEN_4055 : tag_0_71; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6112 = ~quene ? _GEN_4056 : tag_0_72; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6113 = ~quene ? _GEN_4057 : tag_0_73; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6114 = ~quene ? _GEN_4058 : tag_0_74; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6115 = ~quene ? _GEN_4059 : tag_0_75; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6116 = ~quene ? _GEN_4060 : tag_0_76; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6117 = ~quene ? _GEN_4061 : tag_0_77; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6118 = ~quene ? _GEN_4062 : tag_0_78; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6119 = ~quene ? _GEN_4063 : tag_0_79; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6120 = ~quene ? _GEN_4064 : tag_0_80; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6121 = ~quene ? _GEN_4065 : tag_0_81; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6122 = ~quene ? _GEN_4066 : tag_0_82; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6123 = ~quene ? _GEN_4067 : tag_0_83; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6124 = ~quene ? _GEN_4068 : tag_0_84; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6125 = ~quene ? _GEN_4069 : tag_0_85; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6126 = ~quene ? _GEN_4070 : tag_0_86; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6127 = ~quene ? _GEN_4071 : tag_0_87; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6128 = ~quene ? _GEN_4072 : tag_0_88; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6129 = ~quene ? _GEN_4073 : tag_0_89; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6130 = ~quene ? _GEN_4074 : tag_0_90; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6131 = ~quene ? _GEN_4075 : tag_0_91; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6132 = ~quene ? _GEN_4076 : tag_0_92; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6133 = ~quene ? _GEN_4077 : tag_0_93; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6134 = ~quene ? _GEN_4078 : tag_0_94; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6135 = ~quene ? _GEN_4079 : tag_0_95; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6136 = ~quene ? _GEN_4080 : tag_0_96; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6137 = ~quene ? _GEN_4081 : tag_0_97; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6138 = ~quene ? _GEN_4082 : tag_0_98; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6139 = ~quene ? _GEN_4083 : tag_0_99; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6140 = ~quene ? _GEN_4084 : tag_0_100; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6141 = ~quene ? _GEN_4085 : tag_0_101; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6142 = ~quene ? _GEN_4086 : tag_0_102; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6143 = ~quene ? _GEN_4087 : tag_0_103; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6144 = ~quene ? _GEN_4088 : tag_0_104; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6145 = ~quene ? _GEN_4089 : tag_0_105; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6146 = ~quene ? _GEN_4090 : tag_0_106; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6147 = ~quene ? _GEN_4091 : tag_0_107; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6148 = ~quene ? _GEN_4092 : tag_0_108; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6149 = ~quene ? _GEN_4093 : tag_0_109; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6150 = ~quene ? _GEN_4094 : tag_0_110; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6151 = ~quene ? _GEN_4095 : tag_0_111; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6152 = ~quene ? _GEN_4096 : tag_0_112; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6153 = ~quene ? _GEN_4097 : tag_0_113; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6154 = ~quene ? _GEN_4098 : tag_0_114; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6155 = ~quene ? _GEN_4099 : tag_0_115; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6156 = ~quene ? _GEN_4100 : tag_0_116; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6157 = ~quene ? _GEN_4101 : tag_0_117; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6158 = ~quene ? _GEN_4102 : tag_0_118; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6159 = ~quene ? _GEN_4103 : tag_0_119; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6160 = ~quene ? _GEN_4104 : tag_0_120; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6161 = ~quene ? _GEN_4105 : tag_0_121; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6162 = ~quene ? _GEN_4106 : tag_0_122; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6163 = ~quene ? _GEN_4107 : tag_0_123; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6164 = ~quene ? _GEN_4108 : tag_0_124; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6165 = ~quene ? _GEN_4109 : tag_0_125; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6166 = ~quene ? _GEN_4110 : tag_0_126; // @[d_cache.scala 132:34 20:24]
  wire [31:0] _GEN_6167 = ~quene ? _GEN_4111 : tag_0_127; // @[d_cache.scala 132:34 20:24]
  wire  _GEN_6168 = ~quene ? _GEN_4112 : dirty_0_0; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6169 = ~quene ? _GEN_4113 : dirty_0_1; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6170 = ~quene ? _GEN_4114 : dirty_0_2; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6171 = ~quene ? _GEN_4115 : dirty_0_3; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6172 = ~quene ? _GEN_4116 : dirty_0_4; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6173 = ~quene ? _GEN_4117 : dirty_0_5; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6174 = ~quene ? _GEN_4118 : dirty_0_6; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6175 = ~quene ? _GEN_4119 : dirty_0_7; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6176 = ~quene ? _GEN_4120 : dirty_0_8; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6177 = ~quene ? _GEN_4121 : dirty_0_9; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6178 = ~quene ? _GEN_4122 : dirty_0_10; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6179 = ~quene ? _GEN_4123 : dirty_0_11; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6180 = ~quene ? _GEN_4124 : dirty_0_12; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6181 = ~quene ? _GEN_4125 : dirty_0_13; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6182 = ~quene ? _GEN_4126 : dirty_0_14; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6183 = ~quene ? _GEN_4127 : dirty_0_15; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6184 = ~quene ? _GEN_4128 : dirty_0_16; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6185 = ~quene ? _GEN_4129 : dirty_0_17; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6186 = ~quene ? _GEN_4130 : dirty_0_18; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6187 = ~quene ? _GEN_4131 : dirty_0_19; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6188 = ~quene ? _GEN_4132 : dirty_0_20; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6189 = ~quene ? _GEN_4133 : dirty_0_21; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6190 = ~quene ? _GEN_4134 : dirty_0_22; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6191 = ~quene ? _GEN_4135 : dirty_0_23; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6192 = ~quene ? _GEN_4136 : dirty_0_24; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6193 = ~quene ? _GEN_4137 : dirty_0_25; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6194 = ~quene ? _GEN_4138 : dirty_0_26; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6195 = ~quene ? _GEN_4139 : dirty_0_27; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6196 = ~quene ? _GEN_4140 : dirty_0_28; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6197 = ~quene ? _GEN_4141 : dirty_0_29; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6198 = ~quene ? _GEN_4142 : dirty_0_30; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6199 = ~quene ? _GEN_4143 : dirty_0_31; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6200 = ~quene ? _GEN_4144 : dirty_0_32; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6201 = ~quene ? _GEN_4145 : dirty_0_33; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6202 = ~quene ? _GEN_4146 : dirty_0_34; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6203 = ~quene ? _GEN_4147 : dirty_0_35; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6204 = ~quene ? _GEN_4148 : dirty_0_36; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6205 = ~quene ? _GEN_4149 : dirty_0_37; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6206 = ~quene ? _GEN_4150 : dirty_0_38; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6207 = ~quene ? _GEN_4151 : dirty_0_39; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6208 = ~quene ? _GEN_4152 : dirty_0_40; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6209 = ~quene ? _GEN_4153 : dirty_0_41; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6210 = ~quene ? _GEN_4154 : dirty_0_42; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6211 = ~quene ? _GEN_4155 : dirty_0_43; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6212 = ~quene ? _GEN_4156 : dirty_0_44; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6213 = ~quene ? _GEN_4157 : dirty_0_45; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6214 = ~quene ? _GEN_4158 : dirty_0_46; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6215 = ~quene ? _GEN_4159 : dirty_0_47; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6216 = ~quene ? _GEN_4160 : dirty_0_48; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6217 = ~quene ? _GEN_4161 : dirty_0_49; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6218 = ~quene ? _GEN_4162 : dirty_0_50; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6219 = ~quene ? _GEN_4163 : dirty_0_51; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6220 = ~quene ? _GEN_4164 : dirty_0_52; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6221 = ~quene ? _GEN_4165 : dirty_0_53; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6222 = ~quene ? _GEN_4166 : dirty_0_54; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6223 = ~quene ? _GEN_4167 : dirty_0_55; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6224 = ~quene ? _GEN_4168 : dirty_0_56; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6225 = ~quene ? _GEN_4169 : dirty_0_57; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6226 = ~quene ? _GEN_4170 : dirty_0_58; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6227 = ~quene ? _GEN_4171 : dirty_0_59; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6228 = ~quene ? _GEN_4172 : dirty_0_60; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6229 = ~quene ? _GEN_4173 : dirty_0_61; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6230 = ~quene ? _GEN_4174 : dirty_0_62; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6231 = ~quene ? _GEN_4175 : dirty_0_63; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6232 = ~quene ? _GEN_4176 : dirty_0_64; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6233 = ~quene ? _GEN_4177 : dirty_0_65; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6234 = ~quene ? _GEN_4178 : dirty_0_66; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6235 = ~quene ? _GEN_4179 : dirty_0_67; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6236 = ~quene ? _GEN_4180 : dirty_0_68; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6237 = ~quene ? _GEN_4181 : dirty_0_69; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6238 = ~quene ? _GEN_4182 : dirty_0_70; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6239 = ~quene ? _GEN_4183 : dirty_0_71; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6240 = ~quene ? _GEN_4184 : dirty_0_72; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6241 = ~quene ? _GEN_4185 : dirty_0_73; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6242 = ~quene ? _GEN_4186 : dirty_0_74; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6243 = ~quene ? _GEN_4187 : dirty_0_75; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6244 = ~quene ? _GEN_4188 : dirty_0_76; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6245 = ~quene ? _GEN_4189 : dirty_0_77; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6246 = ~quene ? _GEN_4190 : dirty_0_78; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6247 = ~quene ? _GEN_4191 : dirty_0_79; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6248 = ~quene ? _GEN_4192 : dirty_0_80; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6249 = ~quene ? _GEN_4193 : dirty_0_81; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6250 = ~quene ? _GEN_4194 : dirty_0_82; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6251 = ~quene ? _GEN_4195 : dirty_0_83; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6252 = ~quene ? _GEN_4196 : dirty_0_84; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6253 = ~quene ? _GEN_4197 : dirty_0_85; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6254 = ~quene ? _GEN_4198 : dirty_0_86; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6255 = ~quene ? _GEN_4199 : dirty_0_87; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6256 = ~quene ? _GEN_4200 : dirty_0_88; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6257 = ~quene ? _GEN_4201 : dirty_0_89; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6258 = ~quene ? _GEN_4202 : dirty_0_90; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6259 = ~quene ? _GEN_4203 : dirty_0_91; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6260 = ~quene ? _GEN_4204 : dirty_0_92; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6261 = ~quene ? _GEN_4205 : dirty_0_93; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6262 = ~quene ? _GEN_4206 : dirty_0_94; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6263 = ~quene ? _GEN_4207 : dirty_0_95; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6264 = ~quene ? _GEN_4208 : dirty_0_96; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6265 = ~quene ? _GEN_4209 : dirty_0_97; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6266 = ~quene ? _GEN_4210 : dirty_0_98; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6267 = ~quene ? _GEN_4211 : dirty_0_99; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6268 = ~quene ? _GEN_4212 : dirty_0_100; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6269 = ~quene ? _GEN_4213 : dirty_0_101; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6270 = ~quene ? _GEN_4214 : dirty_0_102; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6271 = ~quene ? _GEN_4215 : dirty_0_103; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6272 = ~quene ? _GEN_4216 : dirty_0_104; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6273 = ~quene ? _GEN_4217 : dirty_0_105; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6274 = ~quene ? _GEN_4218 : dirty_0_106; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6275 = ~quene ? _GEN_4219 : dirty_0_107; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6276 = ~quene ? _GEN_4220 : dirty_0_108; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6277 = ~quene ? _GEN_4221 : dirty_0_109; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6278 = ~quene ? _GEN_4222 : dirty_0_110; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6279 = ~quene ? _GEN_4223 : dirty_0_111; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6280 = ~quene ? _GEN_4224 : dirty_0_112; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6281 = ~quene ? _GEN_4225 : dirty_0_113; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6282 = ~quene ? _GEN_4226 : dirty_0_114; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6283 = ~quene ? _GEN_4227 : dirty_0_115; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6284 = ~quene ? _GEN_4228 : dirty_0_116; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6285 = ~quene ? _GEN_4229 : dirty_0_117; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6286 = ~quene ? _GEN_4230 : dirty_0_118; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6287 = ~quene ? _GEN_4231 : dirty_0_119; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6288 = ~quene ? _GEN_4232 : dirty_0_120; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6289 = ~quene ? _GEN_4233 : dirty_0_121; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6290 = ~quene ? _GEN_4234 : dirty_0_122; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6291 = ~quene ? _GEN_4235 : dirty_0_123; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6292 = ~quene ? _GEN_4236 : dirty_0_124; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6293 = ~quene ? _GEN_4237 : dirty_0_125; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6294 = ~quene ? _GEN_4238 : dirty_0_126; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6295 = ~quene ? _GEN_4239 : dirty_0_127; // @[d_cache.scala 132:34 24:26]
  wire  _GEN_6296 = ~quene ? _GEN_4240 : valid_0_0; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6297 = ~quene ? _GEN_4241 : valid_0_1; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6298 = ~quene ? _GEN_4242 : valid_0_2; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6299 = ~quene ? _GEN_4243 : valid_0_3; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6300 = ~quene ? _GEN_4244 : valid_0_4; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6301 = ~quene ? _GEN_4245 : valid_0_5; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6302 = ~quene ? _GEN_4246 : valid_0_6; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6303 = ~quene ? _GEN_4247 : valid_0_7; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6304 = ~quene ? _GEN_4248 : valid_0_8; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6305 = ~quene ? _GEN_4249 : valid_0_9; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6306 = ~quene ? _GEN_4250 : valid_0_10; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6307 = ~quene ? _GEN_4251 : valid_0_11; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6308 = ~quene ? _GEN_4252 : valid_0_12; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6309 = ~quene ? _GEN_4253 : valid_0_13; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6310 = ~quene ? _GEN_4254 : valid_0_14; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6311 = ~quene ? _GEN_4255 : valid_0_15; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6312 = ~quene ? _GEN_4256 : valid_0_16; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6313 = ~quene ? _GEN_4257 : valid_0_17; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6314 = ~quene ? _GEN_4258 : valid_0_18; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6315 = ~quene ? _GEN_4259 : valid_0_19; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6316 = ~quene ? _GEN_4260 : valid_0_20; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6317 = ~quene ? _GEN_4261 : valid_0_21; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6318 = ~quene ? _GEN_4262 : valid_0_22; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6319 = ~quene ? _GEN_4263 : valid_0_23; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6320 = ~quene ? _GEN_4264 : valid_0_24; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6321 = ~quene ? _GEN_4265 : valid_0_25; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6322 = ~quene ? _GEN_4266 : valid_0_26; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6323 = ~quene ? _GEN_4267 : valid_0_27; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6324 = ~quene ? _GEN_4268 : valid_0_28; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6325 = ~quene ? _GEN_4269 : valid_0_29; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6326 = ~quene ? _GEN_4270 : valid_0_30; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6327 = ~quene ? _GEN_4271 : valid_0_31; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6328 = ~quene ? _GEN_4272 : valid_0_32; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6329 = ~quene ? _GEN_4273 : valid_0_33; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6330 = ~quene ? _GEN_4274 : valid_0_34; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6331 = ~quene ? _GEN_4275 : valid_0_35; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6332 = ~quene ? _GEN_4276 : valid_0_36; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6333 = ~quene ? _GEN_4277 : valid_0_37; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6334 = ~quene ? _GEN_4278 : valid_0_38; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6335 = ~quene ? _GEN_4279 : valid_0_39; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6336 = ~quene ? _GEN_4280 : valid_0_40; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6337 = ~quene ? _GEN_4281 : valid_0_41; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6338 = ~quene ? _GEN_4282 : valid_0_42; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6339 = ~quene ? _GEN_4283 : valid_0_43; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6340 = ~quene ? _GEN_4284 : valid_0_44; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6341 = ~quene ? _GEN_4285 : valid_0_45; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6342 = ~quene ? _GEN_4286 : valid_0_46; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6343 = ~quene ? _GEN_4287 : valid_0_47; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6344 = ~quene ? _GEN_4288 : valid_0_48; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6345 = ~quene ? _GEN_4289 : valid_0_49; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6346 = ~quene ? _GEN_4290 : valid_0_50; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6347 = ~quene ? _GEN_4291 : valid_0_51; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6348 = ~quene ? _GEN_4292 : valid_0_52; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6349 = ~quene ? _GEN_4293 : valid_0_53; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6350 = ~quene ? _GEN_4294 : valid_0_54; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6351 = ~quene ? _GEN_4295 : valid_0_55; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6352 = ~quene ? _GEN_4296 : valid_0_56; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6353 = ~quene ? _GEN_4297 : valid_0_57; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6354 = ~quene ? _GEN_4298 : valid_0_58; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6355 = ~quene ? _GEN_4299 : valid_0_59; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6356 = ~quene ? _GEN_4300 : valid_0_60; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6357 = ~quene ? _GEN_4301 : valid_0_61; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6358 = ~quene ? _GEN_4302 : valid_0_62; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6359 = ~quene ? _GEN_4303 : valid_0_63; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6360 = ~quene ? _GEN_4304 : valid_0_64; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6361 = ~quene ? _GEN_4305 : valid_0_65; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6362 = ~quene ? _GEN_4306 : valid_0_66; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6363 = ~quene ? _GEN_4307 : valid_0_67; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6364 = ~quene ? _GEN_4308 : valid_0_68; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6365 = ~quene ? _GEN_4309 : valid_0_69; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6366 = ~quene ? _GEN_4310 : valid_0_70; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6367 = ~quene ? _GEN_4311 : valid_0_71; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6368 = ~quene ? _GEN_4312 : valid_0_72; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6369 = ~quene ? _GEN_4313 : valid_0_73; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6370 = ~quene ? _GEN_4314 : valid_0_74; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6371 = ~quene ? _GEN_4315 : valid_0_75; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6372 = ~quene ? _GEN_4316 : valid_0_76; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6373 = ~quene ? _GEN_4317 : valid_0_77; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6374 = ~quene ? _GEN_4318 : valid_0_78; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6375 = ~quene ? _GEN_4319 : valid_0_79; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6376 = ~quene ? _GEN_4320 : valid_0_80; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6377 = ~quene ? _GEN_4321 : valid_0_81; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6378 = ~quene ? _GEN_4322 : valid_0_82; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6379 = ~quene ? _GEN_4323 : valid_0_83; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6380 = ~quene ? _GEN_4324 : valid_0_84; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6381 = ~quene ? _GEN_4325 : valid_0_85; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6382 = ~quene ? _GEN_4326 : valid_0_86; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6383 = ~quene ? _GEN_4327 : valid_0_87; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6384 = ~quene ? _GEN_4328 : valid_0_88; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6385 = ~quene ? _GEN_4329 : valid_0_89; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6386 = ~quene ? _GEN_4330 : valid_0_90; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6387 = ~quene ? _GEN_4331 : valid_0_91; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6388 = ~quene ? _GEN_4332 : valid_0_92; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6389 = ~quene ? _GEN_4333 : valid_0_93; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6390 = ~quene ? _GEN_4334 : valid_0_94; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6391 = ~quene ? _GEN_4335 : valid_0_95; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6392 = ~quene ? _GEN_4336 : valid_0_96; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6393 = ~quene ? _GEN_4337 : valid_0_97; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6394 = ~quene ? _GEN_4338 : valid_0_98; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6395 = ~quene ? _GEN_4339 : valid_0_99; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6396 = ~quene ? _GEN_4340 : valid_0_100; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6397 = ~quene ? _GEN_4341 : valid_0_101; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6398 = ~quene ? _GEN_4342 : valid_0_102; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6399 = ~quene ? _GEN_4343 : valid_0_103; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6400 = ~quene ? _GEN_4344 : valid_0_104; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6401 = ~quene ? _GEN_4345 : valid_0_105; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6402 = ~quene ? _GEN_4346 : valid_0_106; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6403 = ~quene ? _GEN_4347 : valid_0_107; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6404 = ~quene ? _GEN_4348 : valid_0_108; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6405 = ~quene ? _GEN_4349 : valid_0_109; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6406 = ~quene ? _GEN_4350 : valid_0_110; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6407 = ~quene ? _GEN_4351 : valid_0_111; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6408 = ~quene ? _GEN_4352 : valid_0_112; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6409 = ~quene ? _GEN_4353 : valid_0_113; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6410 = ~quene ? _GEN_4354 : valid_0_114; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6411 = ~quene ? _GEN_4355 : valid_0_115; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6412 = ~quene ? _GEN_4356 : valid_0_116; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6413 = ~quene ? _GEN_4357 : valid_0_117; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6414 = ~quene ? _GEN_4358 : valid_0_118; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6415 = ~quene ? _GEN_4359 : valid_0_119; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6416 = ~quene ? _GEN_4360 : valid_0_120; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6417 = ~quene ? _GEN_4361 : valid_0_121; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6418 = ~quene ? _GEN_4362 : valid_0_122; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6419 = ~quene ? _GEN_4363 : valid_0_123; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6420 = ~quene ? _GEN_4364 : valid_0_124; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6421 = ~quene ? _GEN_4365 : valid_0_125; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6422 = ~quene ? _GEN_4366 : valid_0_126; // @[d_cache.scala 132:34 22:26]
  wire  _GEN_6423 = ~quene ? _GEN_4367 : valid_0_127; // @[d_cache.scala 132:34 22:26]
  wire [2:0] _GEN_6424 = ~quene ? _GEN_4368 : _GEN_5908; // @[d_cache.scala 132:34]
  wire [63:0] _GEN_6426 = ~quene ? ram_1_0 : _GEN_5396; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6427 = ~quene ? ram_1_1 : _GEN_5397; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6428 = ~quene ? ram_1_2 : _GEN_5398; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6429 = ~quene ? ram_1_3 : _GEN_5399; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6430 = ~quene ? ram_1_4 : _GEN_5400; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6431 = ~quene ? ram_1_5 : _GEN_5401; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6432 = ~quene ? ram_1_6 : _GEN_5402; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6433 = ~quene ? ram_1_7 : _GEN_5403; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6434 = ~quene ? ram_1_8 : _GEN_5404; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6435 = ~quene ? ram_1_9 : _GEN_5405; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6436 = ~quene ? ram_1_10 : _GEN_5406; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6437 = ~quene ? ram_1_11 : _GEN_5407; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6438 = ~quene ? ram_1_12 : _GEN_5408; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6439 = ~quene ? ram_1_13 : _GEN_5409; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6440 = ~quene ? ram_1_14 : _GEN_5410; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6441 = ~quene ? ram_1_15 : _GEN_5411; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6442 = ~quene ? ram_1_16 : _GEN_5412; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6443 = ~quene ? ram_1_17 : _GEN_5413; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6444 = ~quene ? ram_1_18 : _GEN_5414; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6445 = ~quene ? ram_1_19 : _GEN_5415; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6446 = ~quene ? ram_1_20 : _GEN_5416; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6447 = ~quene ? ram_1_21 : _GEN_5417; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6448 = ~quene ? ram_1_22 : _GEN_5418; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6449 = ~quene ? ram_1_23 : _GEN_5419; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6450 = ~quene ? ram_1_24 : _GEN_5420; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6451 = ~quene ? ram_1_25 : _GEN_5421; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6452 = ~quene ? ram_1_26 : _GEN_5422; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6453 = ~quene ? ram_1_27 : _GEN_5423; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6454 = ~quene ? ram_1_28 : _GEN_5424; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6455 = ~quene ? ram_1_29 : _GEN_5425; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6456 = ~quene ? ram_1_30 : _GEN_5426; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6457 = ~quene ? ram_1_31 : _GEN_5427; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6458 = ~quene ? ram_1_32 : _GEN_5428; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6459 = ~quene ? ram_1_33 : _GEN_5429; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6460 = ~quene ? ram_1_34 : _GEN_5430; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6461 = ~quene ? ram_1_35 : _GEN_5431; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6462 = ~quene ? ram_1_36 : _GEN_5432; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6463 = ~quene ? ram_1_37 : _GEN_5433; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6464 = ~quene ? ram_1_38 : _GEN_5434; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6465 = ~quene ? ram_1_39 : _GEN_5435; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6466 = ~quene ? ram_1_40 : _GEN_5436; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6467 = ~quene ? ram_1_41 : _GEN_5437; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6468 = ~quene ? ram_1_42 : _GEN_5438; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6469 = ~quene ? ram_1_43 : _GEN_5439; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6470 = ~quene ? ram_1_44 : _GEN_5440; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6471 = ~quene ? ram_1_45 : _GEN_5441; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6472 = ~quene ? ram_1_46 : _GEN_5442; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6473 = ~quene ? ram_1_47 : _GEN_5443; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6474 = ~quene ? ram_1_48 : _GEN_5444; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6475 = ~quene ? ram_1_49 : _GEN_5445; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6476 = ~quene ? ram_1_50 : _GEN_5446; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6477 = ~quene ? ram_1_51 : _GEN_5447; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6478 = ~quene ? ram_1_52 : _GEN_5448; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6479 = ~quene ? ram_1_53 : _GEN_5449; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6480 = ~quene ? ram_1_54 : _GEN_5450; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6481 = ~quene ? ram_1_55 : _GEN_5451; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6482 = ~quene ? ram_1_56 : _GEN_5452; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6483 = ~quene ? ram_1_57 : _GEN_5453; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6484 = ~quene ? ram_1_58 : _GEN_5454; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6485 = ~quene ? ram_1_59 : _GEN_5455; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6486 = ~quene ? ram_1_60 : _GEN_5456; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6487 = ~quene ? ram_1_61 : _GEN_5457; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6488 = ~quene ? ram_1_62 : _GEN_5458; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6489 = ~quene ? ram_1_63 : _GEN_5459; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6490 = ~quene ? ram_1_64 : _GEN_5460; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6491 = ~quene ? ram_1_65 : _GEN_5461; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6492 = ~quene ? ram_1_66 : _GEN_5462; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6493 = ~quene ? ram_1_67 : _GEN_5463; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6494 = ~quene ? ram_1_68 : _GEN_5464; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6495 = ~quene ? ram_1_69 : _GEN_5465; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6496 = ~quene ? ram_1_70 : _GEN_5466; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6497 = ~quene ? ram_1_71 : _GEN_5467; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6498 = ~quene ? ram_1_72 : _GEN_5468; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6499 = ~quene ? ram_1_73 : _GEN_5469; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6500 = ~quene ? ram_1_74 : _GEN_5470; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6501 = ~quene ? ram_1_75 : _GEN_5471; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6502 = ~quene ? ram_1_76 : _GEN_5472; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6503 = ~quene ? ram_1_77 : _GEN_5473; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6504 = ~quene ? ram_1_78 : _GEN_5474; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6505 = ~quene ? ram_1_79 : _GEN_5475; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6506 = ~quene ? ram_1_80 : _GEN_5476; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6507 = ~quene ? ram_1_81 : _GEN_5477; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6508 = ~quene ? ram_1_82 : _GEN_5478; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6509 = ~quene ? ram_1_83 : _GEN_5479; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6510 = ~quene ? ram_1_84 : _GEN_5480; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6511 = ~quene ? ram_1_85 : _GEN_5481; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6512 = ~quene ? ram_1_86 : _GEN_5482; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6513 = ~quene ? ram_1_87 : _GEN_5483; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6514 = ~quene ? ram_1_88 : _GEN_5484; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6515 = ~quene ? ram_1_89 : _GEN_5485; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6516 = ~quene ? ram_1_90 : _GEN_5486; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6517 = ~quene ? ram_1_91 : _GEN_5487; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6518 = ~quene ? ram_1_92 : _GEN_5488; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6519 = ~quene ? ram_1_93 : _GEN_5489; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6520 = ~quene ? ram_1_94 : _GEN_5490; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6521 = ~quene ? ram_1_95 : _GEN_5491; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6522 = ~quene ? ram_1_96 : _GEN_5492; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6523 = ~quene ? ram_1_97 : _GEN_5493; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6524 = ~quene ? ram_1_98 : _GEN_5494; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6525 = ~quene ? ram_1_99 : _GEN_5495; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6526 = ~quene ? ram_1_100 : _GEN_5496; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6527 = ~quene ? ram_1_101 : _GEN_5497; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6528 = ~quene ? ram_1_102 : _GEN_5498; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6529 = ~quene ? ram_1_103 : _GEN_5499; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6530 = ~quene ? ram_1_104 : _GEN_5500; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6531 = ~quene ? ram_1_105 : _GEN_5501; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6532 = ~quene ? ram_1_106 : _GEN_5502; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6533 = ~quene ? ram_1_107 : _GEN_5503; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6534 = ~quene ? ram_1_108 : _GEN_5504; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6535 = ~quene ? ram_1_109 : _GEN_5505; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6536 = ~quene ? ram_1_110 : _GEN_5506; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6537 = ~quene ? ram_1_111 : _GEN_5507; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6538 = ~quene ? ram_1_112 : _GEN_5508; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6539 = ~quene ? ram_1_113 : _GEN_5509; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6540 = ~quene ? ram_1_114 : _GEN_5510; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6541 = ~quene ? ram_1_115 : _GEN_5511; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6542 = ~quene ? ram_1_116 : _GEN_5512; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6543 = ~quene ? ram_1_117 : _GEN_5513; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6544 = ~quene ? ram_1_118 : _GEN_5514; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6545 = ~quene ? ram_1_119 : _GEN_5515; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6546 = ~quene ? ram_1_120 : _GEN_5516; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6547 = ~quene ? ram_1_121 : _GEN_5517; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6548 = ~quene ? ram_1_122 : _GEN_5518; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6549 = ~quene ? ram_1_123 : _GEN_5519; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6550 = ~quene ? ram_1_124 : _GEN_5520; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6551 = ~quene ? ram_1_125 : _GEN_5521; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6552 = ~quene ? ram_1_126 : _GEN_5522; // @[d_cache.scala 132:34 19:24]
  wire [63:0] _GEN_6553 = ~quene ? ram_1_127 : _GEN_5523; // @[d_cache.scala 132:34 19:24]
  wire [31:0] _GEN_6554 = ~quene ? tag_1_0 : _GEN_5524; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6555 = ~quene ? tag_1_1 : _GEN_5525; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6556 = ~quene ? tag_1_2 : _GEN_5526; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6557 = ~quene ? tag_1_3 : _GEN_5527; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6558 = ~quene ? tag_1_4 : _GEN_5528; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6559 = ~quene ? tag_1_5 : _GEN_5529; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6560 = ~quene ? tag_1_6 : _GEN_5530; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6561 = ~quene ? tag_1_7 : _GEN_5531; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6562 = ~quene ? tag_1_8 : _GEN_5532; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6563 = ~quene ? tag_1_9 : _GEN_5533; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6564 = ~quene ? tag_1_10 : _GEN_5534; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6565 = ~quene ? tag_1_11 : _GEN_5535; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6566 = ~quene ? tag_1_12 : _GEN_5536; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6567 = ~quene ? tag_1_13 : _GEN_5537; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6568 = ~quene ? tag_1_14 : _GEN_5538; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6569 = ~quene ? tag_1_15 : _GEN_5539; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6570 = ~quene ? tag_1_16 : _GEN_5540; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6571 = ~quene ? tag_1_17 : _GEN_5541; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6572 = ~quene ? tag_1_18 : _GEN_5542; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6573 = ~quene ? tag_1_19 : _GEN_5543; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6574 = ~quene ? tag_1_20 : _GEN_5544; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6575 = ~quene ? tag_1_21 : _GEN_5545; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6576 = ~quene ? tag_1_22 : _GEN_5546; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6577 = ~quene ? tag_1_23 : _GEN_5547; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6578 = ~quene ? tag_1_24 : _GEN_5548; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6579 = ~quene ? tag_1_25 : _GEN_5549; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6580 = ~quene ? tag_1_26 : _GEN_5550; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6581 = ~quene ? tag_1_27 : _GEN_5551; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6582 = ~quene ? tag_1_28 : _GEN_5552; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6583 = ~quene ? tag_1_29 : _GEN_5553; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6584 = ~quene ? tag_1_30 : _GEN_5554; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6585 = ~quene ? tag_1_31 : _GEN_5555; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6586 = ~quene ? tag_1_32 : _GEN_5556; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6587 = ~quene ? tag_1_33 : _GEN_5557; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6588 = ~quene ? tag_1_34 : _GEN_5558; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6589 = ~quene ? tag_1_35 : _GEN_5559; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6590 = ~quene ? tag_1_36 : _GEN_5560; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6591 = ~quene ? tag_1_37 : _GEN_5561; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6592 = ~quene ? tag_1_38 : _GEN_5562; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6593 = ~quene ? tag_1_39 : _GEN_5563; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6594 = ~quene ? tag_1_40 : _GEN_5564; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6595 = ~quene ? tag_1_41 : _GEN_5565; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6596 = ~quene ? tag_1_42 : _GEN_5566; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6597 = ~quene ? tag_1_43 : _GEN_5567; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6598 = ~quene ? tag_1_44 : _GEN_5568; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6599 = ~quene ? tag_1_45 : _GEN_5569; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6600 = ~quene ? tag_1_46 : _GEN_5570; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6601 = ~quene ? tag_1_47 : _GEN_5571; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6602 = ~quene ? tag_1_48 : _GEN_5572; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6603 = ~quene ? tag_1_49 : _GEN_5573; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6604 = ~quene ? tag_1_50 : _GEN_5574; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6605 = ~quene ? tag_1_51 : _GEN_5575; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6606 = ~quene ? tag_1_52 : _GEN_5576; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6607 = ~quene ? tag_1_53 : _GEN_5577; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6608 = ~quene ? tag_1_54 : _GEN_5578; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6609 = ~quene ? tag_1_55 : _GEN_5579; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6610 = ~quene ? tag_1_56 : _GEN_5580; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6611 = ~quene ? tag_1_57 : _GEN_5581; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6612 = ~quene ? tag_1_58 : _GEN_5582; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6613 = ~quene ? tag_1_59 : _GEN_5583; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6614 = ~quene ? tag_1_60 : _GEN_5584; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6615 = ~quene ? tag_1_61 : _GEN_5585; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6616 = ~quene ? tag_1_62 : _GEN_5586; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6617 = ~quene ? tag_1_63 : _GEN_5587; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6618 = ~quene ? tag_1_64 : _GEN_5588; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6619 = ~quene ? tag_1_65 : _GEN_5589; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6620 = ~quene ? tag_1_66 : _GEN_5590; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6621 = ~quene ? tag_1_67 : _GEN_5591; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6622 = ~quene ? tag_1_68 : _GEN_5592; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6623 = ~quene ? tag_1_69 : _GEN_5593; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6624 = ~quene ? tag_1_70 : _GEN_5594; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6625 = ~quene ? tag_1_71 : _GEN_5595; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6626 = ~quene ? tag_1_72 : _GEN_5596; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6627 = ~quene ? tag_1_73 : _GEN_5597; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6628 = ~quene ? tag_1_74 : _GEN_5598; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6629 = ~quene ? tag_1_75 : _GEN_5599; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6630 = ~quene ? tag_1_76 : _GEN_5600; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6631 = ~quene ? tag_1_77 : _GEN_5601; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6632 = ~quene ? tag_1_78 : _GEN_5602; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6633 = ~quene ? tag_1_79 : _GEN_5603; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6634 = ~quene ? tag_1_80 : _GEN_5604; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6635 = ~quene ? tag_1_81 : _GEN_5605; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6636 = ~quene ? tag_1_82 : _GEN_5606; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6637 = ~quene ? tag_1_83 : _GEN_5607; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6638 = ~quene ? tag_1_84 : _GEN_5608; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6639 = ~quene ? tag_1_85 : _GEN_5609; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6640 = ~quene ? tag_1_86 : _GEN_5610; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6641 = ~quene ? tag_1_87 : _GEN_5611; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6642 = ~quene ? tag_1_88 : _GEN_5612; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6643 = ~quene ? tag_1_89 : _GEN_5613; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6644 = ~quene ? tag_1_90 : _GEN_5614; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6645 = ~quene ? tag_1_91 : _GEN_5615; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6646 = ~quene ? tag_1_92 : _GEN_5616; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6647 = ~quene ? tag_1_93 : _GEN_5617; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6648 = ~quene ? tag_1_94 : _GEN_5618; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6649 = ~quene ? tag_1_95 : _GEN_5619; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6650 = ~quene ? tag_1_96 : _GEN_5620; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6651 = ~quene ? tag_1_97 : _GEN_5621; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6652 = ~quene ? tag_1_98 : _GEN_5622; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6653 = ~quene ? tag_1_99 : _GEN_5623; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6654 = ~quene ? tag_1_100 : _GEN_5624; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6655 = ~quene ? tag_1_101 : _GEN_5625; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6656 = ~quene ? tag_1_102 : _GEN_5626; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6657 = ~quene ? tag_1_103 : _GEN_5627; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6658 = ~quene ? tag_1_104 : _GEN_5628; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6659 = ~quene ? tag_1_105 : _GEN_5629; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6660 = ~quene ? tag_1_106 : _GEN_5630; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6661 = ~quene ? tag_1_107 : _GEN_5631; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6662 = ~quene ? tag_1_108 : _GEN_5632; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6663 = ~quene ? tag_1_109 : _GEN_5633; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6664 = ~quene ? tag_1_110 : _GEN_5634; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6665 = ~quene ? tag_1_111 : _GEN_5635; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6666 = ~quene ? tag_1_112 : _GEN_5636; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6667 = ~quene ? tag_1_113 : _GEN_5637; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6668 = ~quene ? tag_1_114 : _GEN_5638; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6669 = ~quene ? tag_1_115 : _GEN_5639; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6670 = ~quene ? tag_1_116 : _GEN_5640; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6671 = ~quene ? tag_1_117 : _GEN_5641; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6672 = ~quene ? tag_1_118 : _GEN_5642; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6673 = ~quene ? tag_1_119 : _GEN_5643; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6674 = ~quene ? tag_1_120 : _GEN_5644; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6675 = ~quene ? tag_1_121 : _GEN_5645; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6676 = ~quene ? tag_1_122 : _GEN_5646; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6677 = ~quene ? tag_1_123 : _GEN_5647; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6678 = ~quene ? tag_1_124 : _GEN_5648; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6679 = ~quene ? tag_1_125 : _GEN_5649; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6680 = ~quene ? tag_1_126 : _GEN_5650; // @[d_cache.scala 132:34 21:24]
  wire [31:0] _GEN_6681 = ~quene ? tag_1_127 : _GEN_5651; // @[d_cache.scala 132:34 21:24]
  wire  _GEN_6682 = ~quene ? dirty_1_0 : _GEN_5652; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6683 = ~quene ? dirty_1_1 : _GEN_5653; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6684 = ~quene ? dirty_1_2 : _GEN_5654; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6685 = ~quene ? dirty_1_3 : _GEN_5655; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6686 = ~quene ? dirty_1_4 : _GEN_5656; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6687 = ~quene ? dirty_1_5 : _GEN_5657; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6688 = ~quene ? dirty_1_6 : _GEN_5658; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6689 = ~quene ? dirty_1_7 : _GEN_5659; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6690 = ~quene ? dirty_1_8 : _GEN_5660; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6691 = ~quene ? dirty_1_9 : _GEN_5661; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6692 = ~quene ? dirty_1_10 : _GEN_5662; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6693 = ~quene ? dirty_1_11 : _GEN_5663; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6694 = ~quene ? dirty_1_12 : _GEN_5664; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6695 = ~quene ? dirty_1_13 : _GEN_5665; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6696 = ~quene ? dirty_1_14 : _GEN_5666; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6697 = ~quene ? dirty_1_15 : _GEN_5667; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6698 = ~quene ? dirty_1_16 : _GEN_5668; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6699 = ~quene ? dirty_1_17 : _GEN_5669; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6700 = ~quene ? dirty_1_18 : _GEN_5670; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6701 = ~quene ? dirty_1_19 : _GEN_5671; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6702 = ~quene ? dirty_1_20 : _GEN_5672; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6703 = ~quene ? dirty_1_21 : _GEN_5673; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6704 = ~quene ? dirty_1_22 : _GEN_5674; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6705 = ~quene ? dirty_1_23 : _GEN_5675; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6706 = ~quene ? dirty_1_24 : _GEN_5676; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6707 = ~quene ? dirty_1_25 : _GEN_5677; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6708 = ~quene ? dirty_1_26 : _GEN_5678; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6709 = ~quene ? dirty_1_27 : _GEN_5679; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6710 = ~quene ? dirty_1_28 : _GEN_5680; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6711 = ~quene ? dirty_1_29 : _GEN_5681; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6712 = ~quene ? dirty_1_30 : _GEN_5682; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6713 = ~quene ? dirty_1_31 : _GEN_5683; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6714 = ~quene ? dirty_1_32 : _GEN_5684; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6715 = ~quene ? dirty_1_33 : _GEN_5685; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6716 = ~quene ? dirty_1_34 : _GEN_5686; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6717 = ~quene ? dirty_1_35 : _GEN_5687; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6718 = ~quene ? dirty_1_36 : _GEN_5688; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6719 = ~quene ? dirty_1_37 : _GEN_5689; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6720 = ~quene ? dirty_1_38 : _GEN_5690; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6721 = ~quene ? dirty_1_39 : _GEN_5691; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6722 = ~quene ? dirty_1_40 : _GEN_5692; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6723 = ~quene ? dirty_1_41 : _GEN_5693; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6724 = ~quene ? dirty_1_42 : _GEN_5694; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6725 = ~quene ? dirty_1_43 : _GEN_5695; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6726 = ~quene ? dirty_1_44 : _GEN_5696; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6727 = ~quene ? dirty_1_45 : _GEN_5697; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6728 = ~quene ? dirty_1_46 : _GEN_5698; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6729 = ~quene ? dirty_1_47 : _GEN_5699; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6730 = ~quene ? dirty_1_48 : _GEN_5700; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6731 = ~quene ? dirty_1_49 : _GEN_5701; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6732 = ~quene ? dirty_1_50 : _GEN_5702; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6733 = ~quene ? dirty_1_51 : _GEN_5703; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6734 = ~quene ? dirty_1_52 : _GEN_5704; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6735 = ~quene ? dirty_1_53 : _GEN_5705; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6736 = ~quene ? dirty_1_54 : _GEN_5706; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6737 = ~quene ? dirty_1_55 : _GEN_5707; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6738 = ~quene ? dirty_1_56 : _GEN_5708; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6739 = ~quene ? dirty_1_57 : _GEN_5709; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6740 = ~quene ? dirty_1_58 : _GEN_5710; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6741 = ~quene ? dirty_1_59 : _GEN_5711; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6742 = ~quene ? dirty_1_60 : _GEN_5712; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6743 = ~quene ? dirty_1_61 : _GEN_5713; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6744 = ~quene ? dirty_1_62 : _GEN_5714; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6745 = ~quene ? dirty_1_63 : _GEN_5715; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6746 = ~quene ? dirty_1_64 : _GEN_5716; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6747 = ~quene ? dirty_1_65 : _GEN_5717; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6748 = ~quene ? dirty_1_66 : _GEN_5718; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6749 = ~quene ? dirty_1_67 : _GEN_5719; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6750 = ~quene ? dirty_1_68 : _GEN_5720; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6751 = ~quene ? dirty_1_69 : _GEN_5721; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6752 = ~quene ? dirty_1_70 : _GEN_5722; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6753 = ~quene ? dirty_1_71 : _GEN_5723; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6754 = ~quene ? dirty_1_72 : _GEN_5724; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6755 = ~quene ? dirty_1_73 : _GEN_5725; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6756 = ~quene ? dirty_1_74 : _GEN_5726; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6757 = ~quene ? dirty_1_75 : _GEN_5727; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6758 = ~quene ? dirty_1_76 : _GEN_5728; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6759 = ~quene ? dirty_1_77 : _GEN_5729; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6760 = ~quene ? dirty_1_78 : _GEN_5730; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6761 = ~quene ? dirty_1_79 : _GEN_5731; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6762 = ~quene ? dirty_1_80 : _GEN_5732; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6763 = ~quene ? dirty_1_81 : _GEN_5733; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6764 = ~quene ? dirty_1_82 : _GEN_5734; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6765 = ~quene ? dirty_1_83 : _GEN_5735; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6766 = ~quene ? dirty_1_84 : _GEN_5736; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6767 = ~quene ? dirty_1_85 : _GEN_5737; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6768 = ~quene ? dirty_1_86 : _GEN_5738; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6769 = ~quene ? dirty_1_87 : _GEN_5739; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6770 = ~quene ? dirty_1_88 : _GEN_5740; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6771 = ~quene ? dirty_1_89 : _GEN_5741; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6772 = ~quene ? dirty_1_90 : _GEN_5742; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6773 = ~quene ? dirty_1_91 : _GEN_5743; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6774 = ~quene ? dirty_1_92 : _GEN_5744; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6775 = ~quene ? dirty_1_93 : _GEN_5745; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6776 = ~quene ? dirty_1_94 : _GEN_5746; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6777 = ~quene ? dirty_1_95 : _GEN_5747; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6778 = ~quene ? dirty_1_96 : _GEN_5748; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6779 = ~quene ? dirty_1_97 : _GEN_5749; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6780 = ~quene ? dirty_1_98 : _GEN_5750; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6781 = ~quene ? dirty_1_99 : _GEN_5751; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6782 = ~quene ? dirty_1_100 : _GEN_5752; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6783 = ~quene ? dirty_1_101 : _GEN_5753; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6784 = ~quene ? dirty_1_102 : _GEN_5754; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6785 = ~quene ? dirty_1_103 : _GEN_5755; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6786 = ~quene ? dirty_1_104 : _GEN_5756; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6787 = ~quene ? dirty_1_105 : _GEN_5757; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6788 = ~quene ? dirty_1_106 : _GEN_5758; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6789 = ~quene ? dirty_1_107 : _GEN_5759; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6790 = ~quene ? dirty_1_108 : _GEN_5760; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6791 = ~quene ? dirty_1_109 : _GEN_5761; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6792 = ~quene ? dirty_1_110 : _GEN_5762; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6793 = ~quene ? dirty_1_111 : _GEN_5763; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6794 = ~quene ? dirty_1_112 : _GEN_5764; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6795 = ~quene ? dirty_1_113 : _GEN_5765; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6796 = ~quene ? dirty_1_114 : _GEN_5766; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6797 = ~quene ? dirty_1_115 : _GEN_5767; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6798 = ~quene ? dirty_1_116 : _GEN_5768; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6799 = ~quene ? dirty_1_117 : _GEN_5769; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6800 = ~quene ? dirty_1_118 : _GEN_5770; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6801 = ~quene ? dirty_1_119 : _GEN_5771; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6802 = ~quene ? dirty_1_120 : _GEN_5772; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6803 = ~quene ? dirty_1_121 : _GEN_5773; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6804 = ~quene ? dirty_1_122 : _GEN_5774; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6805 = ~quene ? dirty_1_123 : _GEN_5775; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6806 = ~quene ? dirty_1_124 : _GEN_5776; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6807 = ~quene ? dirty_1_125 : _GEN_5777; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6808 = ~quene ? dirty_1_126 : _GEN_5778; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6809 = ~quene ? dirty_1_127 : _GEN_5779; // @[d_cache.scala 132:34 25:26]
  wire  _GEN_6810 = ~quene ? valid_1_0 : _GEN_5780; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6811 = ~quene ? valid_1_1 : _GEN_5781; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6812 = ~quene ? valid_1_2 : _GEN_5782; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6813 = ~quene ? valid_1_3 : _GEN_5783; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6814 = ~quene ? valid_1_4 : _GEN_5784; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6815 = ~quene ? valid_1_5 : _GEN_5785; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6816 = ~quene ? valid_1_6 : _GEN_5786; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6817 = ~quene ? valid_1_7 : _GEN_5787; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6818 = ~quene ? valid_1_8 : _GEN_5788; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6819 = ~quene ? valid_1_9 : _GEN_5789; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6820 = ~quene ? valid_1_10 : _GEN_5790; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6821 = ~quene ? valid_1_11 : _GEN_5791; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6822 = ~quene ? valid_1_12 : _GEN_5792; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6823 = ~quene ? valid_1_13 : _GEN_5793; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6824 = ~quene ? valid_1_14 : _GEN_5794; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6825 = ~quene ? valid_1_15 : _GEN_5795; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6826 = ~quene ? valid_1_16 : _GEN_5796; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6827 = ~quene ? valid_1_17 : _GEN_5797; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6828 = ~quene ? valid_1_18 : _GEN_5798; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6829 = ~quene ? valid_1_19 : _GEN_5799; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6830 = ~quene ? valid_1_20 : _GEN_5800; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6831 = ~quene ? valid_1_21 : _GEN_5801; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6832 = ~quene ? valid_1_22 : _GEN_5802; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6833 = ~quene ? valid_1_23 : _GEN_5803; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6834 = ~quene ? valid_1_24 : _GEN_5804; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6835 = ~quene ? valid_1_25 : _GEN_5805; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6836 = ~quene ? valid_1_26 : _GEN_5806; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6837 = ~quene ? valid_1_27 : _GEN_5807; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6838 = ~quene ? valid_1_28 : _GEN_5808; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6839 = ~quene ? valid_1_29 : _GEN_5809; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6840 = ~quene ? valid_1_30 : _GEN_5810; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6841 = ~quene ? valid_1_31 : _GEN_5811; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6842 = ~quene ? valid_1_32 : _GEN_5812; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6843 = ~quene ? valid_1_33 : _GEN_5813; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6844 = ~quene ? valid_1_34 : _GEN_5814; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6845 = ~quene ? valid_1_35 : _GEN_5815; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6846 = ~quene ? valid_1_36 : _GEN_5816; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6847 = ~quene ? valid_1_37 : _GEN_5817; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6848 = ~quene ? valid_1_38 : _GEN_5818; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6849 = ~quene ? valid_1_39 : _GEN_5819; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6850 = ~quene ? valid_1_40 : _GEN_5820; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6851 = ~quene ? valid_1_41 : _GEN_5821; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6852 = ~quene ? valid_1_42 : _GEN_5822; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6853 = ~quene ? valid_1_43 : _GEN_5823; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6854 = ~quene ? valid_1_44 : _GEN_5824; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6855 = ~quene ? valid_1_45 : _GEN_5825; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6856 = ~quene ? valid_1_46 : _GEN_5826; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6857 = ~quene ? valid_1_47 : _GEN_5827; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6858 = ~quene ? valid_1_48 : _GEN_5828; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6859 = ~quene ? valid_1_49 : _GEN_5829; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6860 = ~quene ? valid_1_50 : _GEN_5830; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6861 = ~quene ? valid_1_51 : _GEN_5831; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6862 = ~quene ? valid_1_52 : _GEN_5832; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6863 = ~quene ? valid_1_53 : _GEN_5833; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6864 = ~quene ? valid_1_54 : _GEN_5834; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6865 = ~quene ? valid_1_55 : _GEN_5835; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6866 = ~quene ? valid_1_56 : _GEN_5836; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6867 = ~quene ? valid_1_57 : _GEN_5837; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6868 = ~quene ? valid_1_58 : _GEN_5838; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6869 = ~quene ? valid_1_59 : _GEN_5839; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6870 = ~quene ? valid_1_60 : _GEN_5840; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6871 = ~quene ? valid_1_61 : _GEN_5841; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6872 = ~quene ? valid_1_62 : _GEN_5842; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6873 = ~quene ? valid_1_63 : _GEN_5843; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6874 = ~quene ? valid_1_64 : _GEN_5844; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6875 = ~quene ? valid_1_65 : _GEN_5845; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6876 = ~quene ? valid_1_66 : _GEN_5846; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6877 = ~quene ? valid_1_67 : _GEN_5847; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6878 = ~quene ? valid_1_68 : _GEN_5848; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6879 = ~quene ? valid_1_69 : _GEN_5849; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6880 = ~quene ? valid_1_70 : _GEN_5850; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6881 = ~quene ? valid_1_71 : _GEN_5851; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6882 = ~quene ? valid_1_72 : _GEN_5852; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6883 = ~quene ? valid_1_73 : _GEN_5853; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6884 = ~quene ? valid_1_74 : _GEN_5854; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6885 = ~quene ? valid_1_75 : _GEN_5855; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6886 = ~quene ? valid_1_76 : _GEN_5856; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6887 = ~quene ? valid_1_77 : _GEN_5857; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6888 = ~quene ? valid_1_78 : _GEN_5858; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6889 = ~quene ? valid_1_79 : _GEN_5859; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6890 = ~quene ? valid_1_80 : _GEN_5860; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6891 = ~quene ? valid_1_81 : _GEN_5861; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6892 = ~quene ? valid_1_82 : _GEN_5862; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6893 = ~quene ? valid_1_83 : _GEN_5863; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6894 = ~quene ? valid_1_84 : _GEN_5864; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6895 = ~quene ? valid_1_85 : _GEN_5865; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6896 = ~quene ? valid_1_86 : _GEN_5866; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6897 = ~quene ? valid_1_87 : _GEN_5867; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6898 = ~quene ? valid_1_88 : _GEN_5868; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6899 = ~quene ? valid_1_89 : _GEN_5869; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6900 = ~quene ? valid_1_90 : _GEN_5870; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6901 = ~quene ? valid_1_91 : _GEN_5871; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6902 = ~quene ? valid_1_92 : _GEN_5872; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6903 = ~quene ? valid_1_93 : _GEN_5873; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6904 = ~quene ? valid_1_94 : _GEN_5874; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6905 = ~quene ? valid_1_95 : _GEN_5875; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6906 = ~quene ? valid_1_96 : _GEN_5876; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6907 = ~quene ? valid_1_97 : _GEN_5877; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6908 = ~quene ? valid_1_98 : _GEN_5878; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6909 = ~quene ? valid_1_99 : _GEN_5879; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6910 = ~quene ? valid_1_100 : _GEN_5880; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6911 = ~quene ? valid_1_101 : _GEN_5881; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6912 = ~quene ? valid_1_102 : _GEN_5882; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6913 = ~quene ? valid_1_103 : _GEN_5883; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6914 = ~quene ? valid_1_104 : _GEN_5884; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6915 = ~quene ? valid_1_105 : _GEN_5885; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6916 = ~quene ? valid_1_106 : _GEN_5886; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6917 = ~quene ? valid_1_107 : _GEN_5887; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6918 = ~quene ? valid_1_108 : _GEN_5888; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6919 = ~quene ? valid_1_109 : _GEN_5889; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6920 = ~quene ? valid_1_110 : _GEN_5890; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6921 = ~quene ? valid_1_111 : _GEN_5891; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6922 = ~quene ? valid_1_112 : _GEN_5892; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6923 = ~quene ? valid_1_113 : _GEN_5893; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6924 = ~quene ? valid_1_114 : _GEN_5894; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6925 = ~quene ? valid_1_115 : _GEN_5895; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6926 = ~quene ? valid_1_116 : _GEN_5896; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6927 = ~quene ? valid_1_117 : _GEN_5897; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6928 = ~quene ? valid_1_118 : _GEN_5898; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6929 = ~quene ? valid_1_119 : _GEN_5899; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6930 = ~quene ? valid_1_120 : _GEN_5900; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6931 = ~quene ? valid_1_121 : _GEN_5901; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6932 = ~quene ? valid_1_122 : _GEN_5902; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6933 = ~quene ? valid_1_123 : _GEN_5903; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6934 = ~quene ? valid_1_124 : _GEN_5904; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6935 = ~quene ? valid_1_125 : _GEN_5905; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6936 = ~quene ? valid_1_126 : _GEN_5906; // @[d_cache.scala 132:34 23:26]
  wire  _GEN_6937 = ~quene ? valid_1_127 : _GEN_5907; // @[d_cache.scala 132:34 23:26]
  wire [2:0] _GEN_6938 = unuse_way == 2'h2 ? 3'h7 : _GEN_6424; // @[d_cache.scala 125:40 126:23]
  wire [63:0] _GEN_6939 = unuse_way == 2'h2 ? _GEN_2446 : _GEN_6426; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6940 = unuse_way == 2'h2 ? _GEN_2447 : _GEN_6427; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6941 = unuse_way == 2'h2 ? _GEN_2448 : _GEN_6428; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6942 = unuse_way == 2'h2 ? _GEN_2449 : _GEN_6429; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6943 = unuse_way == 2'h2 ? _GEN_2450 : _GEN_6430; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6944 = unuse_way == 2'h2 ? _GEN_2451 : _GEN_6431; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6945 = unuse_way == 2'h2 ? _GEN_2452 : _GEN_6432; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6946 = unuse_way == 2'h2 ? _GEN_2453 : _GEN_6433; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6947 = unuse_way == 2'h2 ? _GEN_2454 : _GEN_6434; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6948 = unuse_way == 2'h2 ? _GEN_2455 : _GEN_6435; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6949 = unuse_way == 2'h2 ? _GEN_2456 : _GEN_6436; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6950 = unuse_way == 2'h2 ? _GEN_2457 : _GEN_6437; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6951 = unuse_way == 2'h2 ? _GEN_2458 : _GEN_6438; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6952 = unuse_way == 2'h2 ? _GEN_2459 : _GEN_6439; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6953 = unuse_way == 2'h2 ? _GEN_2460 : _GEN_6440; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6954 = unuse_way == 2'h2 ? _GEN_2461 : _GEN_6441; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6955 = unuse_way == 2'h2 ? _GEN_2462 : _GEN_6442; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6956 = unuse_way == 2'h2 ? _GEN_2463 : _GEN_6443; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6957 = unuse_way == 2'h2 ? _GEN_2464 : _GEN_6444; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6958 = unuse_way == 2'h2 ? _GEN_2465 : _GEN_6445; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6959 = unuse_way == 2'h2 ? _GEN_2466 : _GEN_6446; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6960 = unuse_way == 2'h2 ? _GEN_2467 : _GEN_6447; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6961 = unuse_way == 2'h2 ? _GEN_2468 : _GEN_6448; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6962 = unuse_way == 2'h2 ? _GEN_2469 : _GEN_6449; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6963 = unuse_way == 2'h2 ? _GEN_2470 : _GEN_6450; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6964 = unuse_way == 2'h2 ? _GEN_2471 : _GEN_6451; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6965 = unuse_way == 2'h2 ? _GEN_2472 : _GEN_6452; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6966 = unuse_way == 2'h2 ? _GEN_2473 : _GEN_6453; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6967 = unuse_way == 2'h2 ? _GEN_2474 : _GEN_6454; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6968 = unuse_way == 2'h2 ? _GEN_2475 : _GEN_6455; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6969 = unuse_way == 2'h2 ? _GEN_2476 : _GEN_6456; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6970 = unuse_way == 2'h2 ? _GEN_2477 : _GEN_6457; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6971 = unuse_way == 2'h2 ? _GEN_2478 : _GEN_6458; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6972 = unuse_way == 2'h2 ? _GEN_2479 : _GEN_6459; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6973 = unuse_way == 2'h2 ? _GEN_2480 : _GEN_6460; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6974 = unuse_way == 2'h2 ? _GEN_2481 : _GEN_6461; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6975 = unuse_way == 2'h2 ? _GEN_2482 : _GEN_6462; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6976 = unuse_way == 2'h2 ? _GEN_2483 : _GEN_6463; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6977 = unuse_way == 2'h2 ? _GEN_2484 : _GEN_6464; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6978 = unuse_way == 2'h2 ? _GEN_2485 : _GEN_6465; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6979 = unuse_way == 2'h2 ? _GEN_2486 : _GEN_6466; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6980 = unuse_way == 2'h2 ? _GEN_2487 : _GEN_6467; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6981 = unuse_way == 2'h2 ? _GEN_2488 : _GEN_6468; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6982 = unuse_way == 2'h2 ? _GEN_2489 : _GEN_6469; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6983 = unuse_way == 2'h2 ? _GEN_2490 : _GEN_6470; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6984 = unuse_way == 2'h2 ? _GEN_2491 : _GEN_6471; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6985 = unuse_way == 2'h2 ? _GEN_2492 : _GEN_6472; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6986 = unuse_way == 2'h2 ? _GEN_2493 : _GEN_6473; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6987 = unuse_way == 2'h2 ? _GEN_2494 : _GEN_6474; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6988 = unuse_way == 2'h2 ? _GEN_2495 : _GEN_6475; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6989 = unuse_way == 2'h2 ? _GEN_2496 : _GEN_6476; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6990 = unuse_way == 2'h2 ? _GEN_2497 : _GEN_6477; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6991 = unuse_way == 2'h2 ? _GEN_2498 : _GEN_6478; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6992 = unuse_way == 2'h2 ? _GEN_2499 : _GEN_6479; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6993 = unuse_way == 2'h2 ? _GEN_2500 : _GEN_6480; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6994 = unuse_way == 2'h2 ? _GEN_2501 : _GEN_6481; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6995 = unuse_way == 2'h2 ? _GEN_2502 : _GEN_6482; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6996 = unuse_way == 2'h2 ? _GEN_2503 : _GEN_6483; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6997 = unuse_way == 2'h2 ? _GEN_2504 : _GEN_6484; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6998 = unuse_way == 2'h2 ? _GEN_2505 : _GEN_6485; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_6999 = unuse_way == 2'h2 ? _GEN_2506 : _GEN_6486; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7000 = unuse_way == 2'h2 ? _GEN_2507 : _GEN_6487; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7001 = unuse_way == 2'h2 ? _GEN_2508 : _GEN_6488; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7002 = unuse_way == 2'h2 ? _GEN_2509 : _GEN_6489; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7003 = unuse_way == 2'h2 ? _GEN_2510 : _GEN_6490; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7004 = unuse_way == 2'h2 ? _GEN_2511 : _GEN_6491; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7005 = unuse_way == 2'h2 ? _GEN_2512 : _GEN_6492; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7006 = unuse_way == 2'h2 ? _GEN_2513 : _GEN_6493; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7007 = unuse_way == 2'h2 ? _GEN_2514 : _GEN_6494; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7008 = unuse_way == 2'h2 ? _GEN_2515 : _GEN_6495; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7009 = unuse_way == 2'h2 ? _GEN_2516 : _GEN_6496; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7010 = unuse_way == 2'h2 ? _GEN_2517 : _GEN_6497; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7011 = unuse_way == 2'h2 ? _GEN_2518 : _GEN_6498; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7012 = unuse_way == 2'h2 ? _GEN_2519 : _GEN_6499; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7013 = unuse_way == 2'h2 ? _GEN_2520 : _GEN_6500; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7014 = unuse_way == 2'h2 ? _GEN_2521 : _GEN_6501; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7015 = unuse_way == 2'h2 ? _GEN_2522 : _GEN_6502; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7016 = unuse_way == 2'h2 ? _GEN_2523 : _GEN_6503; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7017 = unuse_way == 2'h2 ? _GEN_2524 : _GEN_6504; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7018 = unuse_way == 2'h2 ? _GEN_2525 : _GEN_6505; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7019 = unuse_way == 2'h2 ? _GEN_2526 : _GEN_6506; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7020 = unuse_way == 2'h2 ? _GEN_2527 : _GEN_6507; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7021 = unuse_way == 2'h2 ? _GEN_2528 : _GEN_6508; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7022 = unuse_way == 2'h2 ? _GEN_2529 : _GEN_6509; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7023 = unuse_way == 2'h2 ? _GEN_2530 : _GEN_6510; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7024 = unuse_way == 2'h2 ? _GEN_2531 : _GEN_6511; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7025 = unuse_way == 2'h2 ? _GEN_2532 : _GEN_6512; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7026 = unuse_way == 2'h2 ? _GEN_2533 : _GEN_6513; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7027 = unuse_way == 2'h2 ? _GEN_2534 : _GEN_6514; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7028 = unuse_way == 2'h2 ? _GEN_2535 : _GEN_6515; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7029 = unuse_way == 2'h2 ? _GEN_2536 : _GEN_6516; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7030 = unuse_way == 2'h2 ? _GEN_2537 : _GEN_6517; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7031 = unuse_way == 2'h2 ? _GEN_2538 : _GEN_6518; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7032 = unuse_way == 2'h2 ? _GEN_2539 : _GEN_6519; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7033 = unuse_way == 2'h2 ? _GEN_2540 : _GEN_6520; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7034 = unuse_way == 2'h2 ? _GEN_2541 : _GEN_6521; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7035 = unuse_way == 2'h2 ? _GEN_2542 : _GEN_6522; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7036 = unuse_way == 2'h2 ? _GEN_2543 : _GEN_6523; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7037 = unuse_way == 2'h2 ? _GEN_2544 : _GEN_6524; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7038 = unuse_way == 2'h2 ? _GEN_2545 : _GEN_6525; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7039 = unuse_way == 2'h2 ? _GEN_2546 : _GEN_6526; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7040 = unuse_way == 2'h2 ? _GEN_2547 : _GEN_6527; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7041 = unuse_way == 2'h2 ? _GEN_2548 : _GEN_6528; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7042 = unuse_way == 2'h2 ? _GEN_2549 : _GEN_6529; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7043 = unuse_way == 2'h2 ? _GEN_2550 : _GEN_6530; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7044 = unuse_way == 2'h2 ? _GEN_2551 : _GEN_6531; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7045 = unuse_way == 2'h2 ? _GEN_2552 : _GEN_6532; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7046 = unuse_way == 2'h2 ? _GEN_2553 : _GEN_6533; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7047 = unuse_way == 2'h2 ? _GEN_2554 : _GEN_6534; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7048 = unuse_way == 2'h2 ? _GEN_2555 : _GEN_6535; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7049 = unuse_way == 2'h2 ? _GEN_2556 : _GEN_6536; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7050 = unuse_way == 2'h2 ? _GEN_2557 : _GEN_6537; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7051 = unuse_way == 2'h2 ? _GEN_2558 : _GEN_6538; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7052 = unuse_way == 2'h2 ? _GEN_2559 : _GEN_6539; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7053 = unuse_way == 2'h2 ? _GEN_2560 : _GEN_6540; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7054 = unuse_way == 2'h2 ? _GEN_2561 : _GEN_6541; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7055 = unuse_way == 2'h2 ? _GEN_2562 : _GEN_6542; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7056 = unuse_way == 2'h2 ? _GEN_2563 : _GEN_6543; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7057 = unuse_way == 2'h2 ? _GEN_2564 : _GEN_6544; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7058 = unuse_way == 2'h2 ? _GEN_2565 : _GEN_6545; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7059 = unuse_way == 2'h2 ? _GEN_2566 : _GEN_6546; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7060 = unuse_way == 2'h2 ? _GEN_2567 : _GEN_6547; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7061 = unuse_way == 2'h2 ? _GEN_2568 : _GEN_6548; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7062 = unuse_way == 2'h2 ? _GEN_2569 : _GEN_6549; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7063 = unuse_way == 2'h2 ? _GEN_2570 : _GEN_6550; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7064 = unuse_way == 2'h2 ? _GEN_2571 : _GEN_6551; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7065 = unuse_way == 2'h2 ? _GEN_2572 : _GEN_6552; // @[d_cache.scala 125:40]
  wire [63:0] _GEN_7066 = unuse_way == 2'h2 ? _GEN_2573 : _GEN_6553; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7067 = unuse_way == 2'h2 ? _GEN_2574 : _GEN_6554; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7068 = unuse_way == 2'h2 ? _GEN_2575 : _GEN_6555; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7069 = unuse_way == 2'h2 ? _GEN_2576 : _GEN_6556; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7070 = unuse_way == 2'h2 ? _GEN_2577 : _GEN_6557; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7071 = unuse_way == 2'h2 ? _GEN_2578 : _GEN_6558; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7072 = unuse_way == 2'h2 ? _GEN_2579 : _GEN_6559; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7073 = unuse_way == 2'h2 ? _GEN_2580 : _GEN_6560; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7074 = unuse_way == 2'h2 ? _GEN_2581 : _GEN_6561; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7075 = unuse_way == 2'h2 ? _GEN_2582 : _GEN_6562; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7076 = unuse_way == 2'h2 ? _GEN_2583 : _GEN_6563; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7077 = unuse_way == 2'h2 ? _GEN_2584 : _GEN_6564; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7078 = unuse_way == 2'h2 ? _GEN_2585 : _GEN_6565; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7079 = unuse_way == 2'h2 ? _GEN_2586 : _GEN_6566; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7080 = unuse_way == 2'h2 ? _GEN_2587 : _GEN_6567; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7081 = unuse_way == 2'h2 ? _GEN_2588 : _GEN_6568; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7082 = unuse_way == 2'h2 ? _GEN_2589 : _GEN_6569; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7083 = unuse_way == 2'h2 ? _GEN_2590 : _GEN_6570; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7084 = unuse_way == 2'h2 ? _GEN_2591 : _GEN_6571; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7085 = unuse_way == 2'h2 ? _GEN_2592 : _GEN_6572; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7086 = unuse_way == 2'h2 ? _GEN_2593 : _GEN_6573; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7087 = unuse_way == 2'h2 ? _GEN_2594 : _GEN_6574; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7088 = unuse_way == 2'h2 ? _GEN_2595 : _GEN_6575; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7089 = unuse_way == 2'h2 ? _GEN_2596 : _GEN_6576; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7090 = unuse_way == 2'h2 ? _GEN_2597 : _GEN_6577; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7091 = unuse_way == 2'h2 ? _GEN_2598 : _GEN_6578; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7092 = unuse_way == 2'h2 ? _GEN_2599 : _GEN_6579; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7093 = unuse_way == 2'h2 ? _GEN_2600 : _GEN_6580; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7094 = unuse_way == 2'h2 ? _GEN_2601 : _GEN_6581; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7095 = unuse_way == 2'h2 ? _GEN_2602 : _GEN_6582; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7096 = unuse_way == 2'h2 ? _GEN_2603 : _GEN_6583; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7097 = unuse_way == 2'h2 ? _GEN_2604 : _GEN_6584; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7098 = unuse_way == 2'h2 ? _GEN_2605 : _GEN_6585; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7099 = unuse_way == 2'h2 ? _GEN_2606 : _GEN_6586; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7100 = unuse_way == 2'h2 ? _GEN_2607 : _GEN_6587; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7101 = unuse_way == 2'h2 ? _GEN_2608 : _GEN_6588; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7102 = unuse_way == 2'h2 ? _GEN_2609 : _GEN_6589; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7103 = unuse_way == 2'h2 ? _GEN_2610 : _GEN_6590; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7104 = unuse_way == 2'h2 ? _GEN_2611 : _GEN_6591; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7105 = unuse_way == 2'h2 ? _GEN_2612 : _GEN_6592; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7106 = unuse_way == 2'h2 ? _GEN_2613 : _GEN_6593; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7107 = unuse_way == 2'h2 ? _GEN_2614 : _GEN_6594; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7108 = unuse_way == 2'h2 ? _GEN_2615 : _GEN_6595; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7109 = unuse_way == 2'h2 ? _GEN_2616 : _GEN_6596; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7110 = unuse_way == 2'h2 ? _GEN_2617 : _GEN_6597; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7111 = unuse_way == 2'h2 ? _GEN_2618 : _GEN_6598; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7112 = unuse_way == 2'h2 ? _GEN_2619 : _GEN_6599; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7113 = unuse_way == 2'h2 ? _GEN_2620 : _GEN_6600; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7114 = unuse_way == 2'h2 ? _GEN_2621 : _GEN_6601; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7115 = unuse_way == 2'h2 ? _GEN_2622 : _GEN_6602; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7116 = unuse_way == 2'h2 ? _GEN_2623 : _GEN_6603; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7117 = unuse_way == 2'h2 ? _GEN_2624 : _GEN_6604; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7118 = unuse_way == 2'h2 ? _GEN_2625 : _GEN_6605; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7119 = unuse_way == 2'h2 ? _GEN_2626 : _GEN_6606; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7120 = unuse_way == 2'h2 ? _GEN_2627 : _GEN_6607; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7121 = unuse_way == 2'h2 ? _GEN_2628 : _GEN_6608; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7122 = unuse_way == 2'h2 ? _GEN_2629 : _GEN_6609; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7123 = unuse_way == 2'h2 ? _GEN_2630 : _GEN_6610; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7124 = unuse_way == 2'h2 ? _GEN_2631 : _GEN_6611; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7125 = unuse_way == 2'h2 ? _GEN_2632 : _GEN_6612; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7126 = unuse_way == 2'h2 ? _GEN_2633 : _GEN_6613; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7127 = unuse_way == 2'h2 ? _GEN_2634 : _GEN_6614; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7128 = unuse_way == 2'h2 ? _GEN_2635 : _GEN_6615; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7129 = unuse_way == 2'h2 ? _GEN_2636 : _GEN_6616; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7130 = unuse_way == 2'h2 ? _GEN_2637 : _GEN_6617; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7131 = unuse_way == 2'h2 ? _GEN_2638 : _GEN_6618; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7132 = unuse_way == 2'h2 ? _GEN_2639 : _GEN_6619; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7133 = unuse_way == 2'h2 ? _GEN_2640 : _GEN_6620; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7134 = unuse_way == 2'h2 ? _GEN_2641 : _GEN_6621; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7135 = unuse_way == 2'h2 ? _GEN_2642 : _GEN_6622; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7136 = unuse_way == 2'h2 ? _GEN_2643 : _GEN_6623; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7137 = unuse_way == 2'h2 ? _GEN_2644 : _GEN_6624; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7138 = unuse_way == 2'h2 ? _GEN_2645 : _GEN_6625; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7139 = unuse_way == 2'h2 ? _GEN_2646 : _GEN_6626; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7140 = unuse_way == 2'h2 ? _GEN_2647 : _GEN_6627; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7141 = unuse_way == 2'h2 ? _GEN_2648 : _GEN_6628; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7142 = unuse_way == 2'h2 ? _GEN_2649 : _GEN_6629; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7143 = unuse_way == 2'h2 ? _GEN_2650 : _GEN_6630; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7144 = unuse_way == 2'h2 ? _GEN_2651 : _GEN_6631; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7145 = unuse_way == 2'h2 ? _GEN_2652 : _GEN_6632; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7146 = unuse_way == 2'h2 ? _GEN_2653 : _GEN_6633; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7147 = unuse_way == 2'h2 ? _GEN_2654 : _GEN_6634; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7148 = unuse_way == 2'h2 ? _GEN_2655 : _GEN_6635; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7149 = unuse_way == 2'h2 ? _GEN_2656 : _GEN_6636; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7150 = unuse_way == 2'h2 ? _GEN_2657 : _GEN_6637; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7151 = unuse_way == 2'h2 ? _GEN_2658 : _GEN_6638; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7152 = unuse_way == 2'h2 ? _GEN_2659 : _GEN_6639; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7153 = unuse_way == 2'h2 ? _GEN_2660 : _GEN_6640; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7154 = unuse_way == 2'h2 ? _GEN_2661 : _GEN_6641; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7155 = unuse_way == 2'h2 ? _GEN_2662 : _GEN_6642; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7156 = unuse_way == 2'h2 ? _GEN_2663 : _GEN_6643; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7157 = unuse_way == 2'h2 ? _GEN_2664 : _GEN_6644; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7158 = unuse_way == 2'h2 ? _GEN_2665 : _GEN_6645; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7159 = unuse_way == 2'h2 ? _GEN_2666 : _GEN_6646; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7160 = unuse_way == 2'h2 ? _GEN_2667 : _GEN_6647; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7161 = unuse_way == 2'h2 ? _GEN_2668 : _GEN_6648; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7162 = unuse_way == 2'h2 ? _GEN_2669 : _GEN_6649; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7163 = unuse_way == 2'h2 ? _GEN_2670 : _GEN_6650; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7164 = unuse_way == 2'h2 ? _GEN_2671 : _GEN_6651; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7165 = unuse_way == 2'h2 ? _GEN_2672 : _GEN_6652; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7166 = unuse_way == 2'h2 ? _GEN_2673 : _GEN_6653; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7167 = unuse_way == 2'h2 ? _GEN_2674 : _GEN_6654; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7168 = unuse_way == 2'h2 ? _GEN_2675 : _GEN_6655; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7169 = unuse_way == 2'h2 ? _GEN_2676 : _GEN_6656; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7170 = unuse_way == 2'h2 ? _GEN_2677 : _GEN_6657; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7171 = unuse_way == 2'h2 ? _GEN_2678 : _GEN_6658; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7172 = unuse_way == 2'h2 ? _GEN_2679 : _GEN_6659; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7173 = unuse_way == 2'h2 ? _GEN_2680 : _GEN_6660; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7174 = unuse_way == 2'h2 ? _GEN_2681 : _GEN_6661; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7175 = unuse_way == 2'h2 ? _GEN_2682 : _GEN_6662; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7176 = unuse_way == 2'h2 ? _GEN_2683 : _GEN_6663; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7177 = unuse_way == 2'h2 ? _GEN_2684 : _GEN_6664; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7178 = unuse_way == 2'h2 ? _GEN_2685 : _GEN_6665; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7179 = unuse_way == 2'h2 ? _GEN_2686 : _GEN_6666; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7180 = unuse_way == 2'h2 ? _GEN_2687 : _GEN_6667; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7181 = unuse_way == 2'h2 ? _GEN_2688 : _GEN_6668; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7182 = unuse_way == 2'h2 ? _GEN_2689 : _GEN_6669; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7183 = unuse_way == 2'h2 ? _GEN_2690 : _GEN_6670; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7184 = unuse_way == 2'h2 ? _GEN_2691 : _GEN_6671; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7185 = unuse_way == 2'h2 ? _GEN_2692 : _GEN_6672; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7186 = unuse_way == 2'h2 ? _GEN_2693 : _GEN_6673; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7187 = unuse_way == 2'h2 ? _GEN_2694 : _GEN_6674; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7188 = unuse_way == 2'h2 ? _GEN_2695 : _GEN_6675; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7189 = unuse_way == 2'h2 ? _GEN_2696 : _GEN_6676; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7190 = unuse_way == 2'h2 ? _GEN_2697 : _GEN_6677; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7191 = unuse_way == 2'h2 ? _GEN_2698 : _GEN_6678; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7192 = unuse_way == 2'h2 ? _GEN_2699 : _GEN_6679; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7193 = unuse_way == 2'h2 ? _GEN_2700 : _GEN_6680; // @[d_cache.scala 125:40]
  wire [31:0] _GEN_7194 = unuse_way == 2'h2 ? _GEN_2701 : _GEN_6681; // @[d_cache.scala 125:40]
  wire  _GEN_7195 = unuse_way == 2'h2 ? _GEN_2702 : _GEN_6810; // @[d_cache.scala 125:40]
  wire  _GEN_7196 = unuse_way == 2'h2 ? _GEN_2703 : _GEN_6811; // @[d_cache.scala 125:40]
  wire  _GEN_7197 = unuse_way == 2'h2 ? _GEN_2704 : _GEN_6812; // @[d_cache.scala 125:40]
  wire  _GEN_7198 = unuse_way == 2'h2 ? _GEN_2705 : _GEN_6813; // @[d_cache.scala 125:40]
  wire  _GEN_7199 = unuse_way == 2'h2 ? _GEN_2706 : _GEN_6814; // @[d_cache.scala 125:40]
  wire  _GEN_7200 = unuse_way == 2'h2 ? _GEN_2707 : _GEN_6815; // @[d_cache.scala 125:40]
  wire  _GEN_7201 = unuse_way == 2'h2 ? _GEN_2708 : _GEN_6816; // @[d_cache.scala 125:40]
  wire  _GEN_7202 = unuse_way == 2'h2 ? _GEN_2709 : _GEN_6817; // @[d_cache.scala 125:40]
  wire  _GEN_7203 = unuse_way == 2'h2 ? _GEN_2710 : _GEN_6818; // @[d_cache.scala 125:40]
  wire  _GEN_7204 = unuse_way == 2'h2 ? _GEN_2711 : _GEN_6819; // @[d_cache.scala 125:40]
  wire  _GEN_7205 = unuse_way == 2'h2 ? _GEN_2712 : _GEN_6820; // @[d_cache.scala 125:40]
  wire  _GEN_7206 = unuse_way == 2'h2 ? _GEN_2713 : _GEN_6821; // @[d_cache.scala 125:40]
  wire  _GEN_7207 = unuse_way == 2'h2 ? _GEN_2714 : _GEN_6822; // @[d_cache.scala 125:40]
  wire  _GEN_7208 = unuse_way == 2'h2 ? _GEN_2715 : _GEN_6823; // @[d_cache.scala 125:40]
  wire  _GEN_7209 = unuse_way == 2'h2 ? _GEN_2716 : _GEN_6824; // @[d_cache.scala 125:40]
  wire  _GEN_7210 = unuse_way == 2'h2 ? _GEN_2717 : _GEN_6825; // @[d_cache.scala 125:40]
  wire  _GEN_7211 = unuse_way == 2'h2 ? _GEN_2718 : _GEN_6826; // @[d_cache.scala 125:40]
  wire  _GEN_7212 = unuse_way == 2'h2 ? _GEN_2719 : _GEN_6827; // @[d_cache.scala 125:40]
  wire  _GEN_7213 = unuse_way == 2'h2 ? _GEN_2720 : _GEN_6828; // @[d_cache.scala 125:40]
  wire  _GEN_7214 = unuse_way == 2'h2 ? _GEN_2721 : _GEN_6829; // @[d_cache.scala 125:40]
  wire  _GEN_7215 = unuse_way == 2'h2 ? _GEN_2722 : _GEN_6830; // @[d_cache.scala 125:40]
  wire  _GEN_7216 = unuse_way == 2'h2 ? _GEN_2723 : _GEN_6831; // @[d_cache.scala 125:40]
  wire  _GEN_7217 = unuse_way == 2'h2 ? _GEN_2724 : _GEN_6832; // @[d_cache.scala 125:40]
  wire  _GEN_7218 = unuse_way == 2'h2 ? _GEN_2725 : _GEN_6833; // @[d_cache.scala 125:40]
  wire  _GEN_7219 = unuse_way == 2'h2 ? _GEN_2726 : _GEN_6834; // @[d_cache.scala 125:40]
  wire  _GEN_7220 = unuse_way == 2'h2 ? _GEN_2727 : _GEN_6835; // @[d_cache.scala 125:40]
  wire  _GEN_7221 = unuse_way == 2'h2 ? _GEN_2728 : _GEN_6836; // @[d_cache.scala 125:40]
  wire  _GEN_7222 = unuse_way == 2'h2 ? _GEN_2729 : _GEN_6837; // @[d_cache.scala 125:40]
  wire  _GEN_7223 = unuse_way == 2'h2 ? _GEN_2730 : _GEN_6838; // @[d_cache.scala 125:40]
  wire  _GEN_7224 = unuse_way == 2'h2 ? _GEN_2731 : _GEN_6839; // @[d_cache.scala 125:40]
  wire  _GEN_7225 = unuse_way == 2'h2 ? _GEN_2732 : _GEN_6840; // @[d_cache.scala 125:40]
  wire  _GEN_7226 = unuse_way == 2'h2 ? _GEN_2733 : _GEN_6841; // @[d_cache.scala 125:40]
  wire  _GEN_7227 = unuse_way == 2'h2 ? _GEN_2734 : _GEN_6842; // @[d_cache.scala 125:40]
  wire  _GEN_7228 = unuse_way == 2'h2 ? _GEN_2735 : _GEN_6843; // @[d_cache.scala 125:40]
  wire  _GEN_7229 = unuse_way == 2'h2 ? _GEN_2736 : _GEN_6844; // @[d_cache.scala 125:40]
  wire  _GEN_7230 = unuse_way == 2'h2 ? _GEN_2737 : _GEN_6845; // @[d_cache.scala 125:40]
  wire  _GEN_7231 = unuse_way == 2'h2 ? _GEN_2738 : _GEN_6846; // @[d_cache.scala 125:40]
  wire  _GEN_7232 = unuse_way == 2'h2 ? _GEN_2739 : _GEN_6847; // @[d_cache.scala 125:40]
  wire  _GEN_7233 = unuse_way == 2'h2 ? _GEN_2740 : _GEN_6848; // @[d_cache.scala 125:40]
  wire  _GEN_7234 = unuse_way == 2'h2 ? _GEN_2741 : _GEN_6849; // @[d_cache.scala 125:40]
  wire  _GEN_7235 = unuse_way == 2'h2 ? _GEN_2742 : _GEN_6850; // @[d_cache.scala 125:40]
  wire  _GEN_7236 = unuse_way == 2'h2 ? _GEN_2743 : _GEN_6851; // @[d_cache.scala 125:40]
  wire  _GEN_7237 = unuse_way == 2'h2 ? _GEN_2744 : _GEN_6852; // @[d_cache.scala 125:40]
  wire  _GEN_7238 = unuse_way == 2'h2 ? _GEN_2745 : _GEN_6853; // @[d_cache.scala 125:40]
  wire  _GEN_7239 = unuse_way == 2'h2 ? _GEN_2746 : _GEN_6854; // @[d_cache.scala 125:40]
  wire  _GEN_7240 = unuse_way == 2'h2 ? _GEN_2747 : _GEN_6855; // @[d_cache.scala 125:40]
  wire  _GEN_7241 = unuse_way == 2'h2 ? _GEN_2748 : _GEN_6856; // @[d_cache.scala 125:40]
  wire  _GEN_7242 = unuse_way == 2'h2 ? _GEN_2749 : _GEN_6857; // @[d_cache.scala 125:40]
  wire  _GEN_7243 = unuse_way == 2'h2 ? _GEN_2750 : _GEN_6858; // @[d_cache.scala 125:40]
  wire  _GEN_7244 = unuse_way == 2'h2 ? _GEN_2751 : _GEN_6859; // @[d_cache.scala 125:40]
  wire  _GEN_7245 = unuse_way == 2'h2 ? _GEN_2752 : _GEN_6860; // @[d_cache.scala 125:40]
  wire  _GEN_7246 = unuse_way == 2'h2 ? _GEN_2753 : _GEN_6861; // @[d_cache.scala 125:40]
  wire  _GEN_7247 = unuse_way == 2'h2 ? _GEN_2754 : _GEN_6862; // @[d_cache.scala 125:40]
  wire  _GEN_7248 = unuse_way == 2'h2 ? _GEN_2755 : _GEN_6863; // @[d_cache.scala 125:40]
  wire  _GEN_7249 = unuse_way == 2'h2 ? _GEN_2756 : _GEN_6864; // @[d_cache.scala 125:40]
  wire  _GEN_7250 = unuse_way == 2'h2 ? _GEN_2757 : _GEN_6865; // @[d_cache.scala 125:40]
  wire  _GEN_7251 = unuse_way == 2'h2 ? _GEN_2758 : _GEN_6866; // @[d_cache.scala 125:40]
  wire  _GEN_7252 = unuse_way == 2'h2 ? _GEN_2759 : _GEN_6867; // @[d_cache.scala 125:40]
  wire  _GEN_7253 = unuse_way == 2'h2 ? _GEN_2760 : _GEN_6868; // @[d_cache.scala 125:40]
  wire  _GEN_7254 = unuse_way == 2'h2 ? _GEN_2761 : _GEN_6869; // @[d_cache.scala 125:40]
  wire  _GEN_7255 = unuse_way == 2'h2 ? _GEN_2762 : _GEN_6870; // @[d_cache.scala 125:40]
  wire  _GEN_7256 = unuse_way == 2'h2 ? _GEN_2763 : _GEN_6871; // @[d_cache.scala 125:40]
  wire  _GEN_7257 = unuse_way == 2'h2 ? _GEN_2764 : _GEN_6872; // @[d_cache.scala 125:40]
  wire  _GEN_7258 = unuse_way == 2'h2 ? _GEN_2765 : _GEN_6873; // @[d_cache.scala 125:40]
  wire  _GEN_7259 = unuse_way == 2'h2 ? _GEN_2766 : _GEN_6874; // @[d_cache.scala 125:40]
  wire  _GEN_7260 = unuse_way == 2'h2 ? _GEN_2767 : _GEN_6875; // @[d_cache.scala 125:40]
  wire  _GEN_7261 = unuse_way == 2'h2 ? _GEN_2768 : _GEN_6876; // @[d_cache.scala 125:40]
  wire  _GEN_7262 = unuse_way == 2'h2 ? _GEN_2769 : _GEN_6877; // @[d_cache.scala 125:40]
  wire  _GEN_7263 = unuse_way == 2'h2 ? _GEN_2770 : _GEN_6878; // @[d_cache.scala 125:40]
  wire  _GEN_7264 = unuse_way == 2'h2 ? _GEN_2771 : _GEN_6879; // @[d_cache.scala 125:40]
  wire  _GEN_7265 = unuse_way == 2'h2 ? _GEN_2772 : _GEN_6880; // @[d_cache.scala 125:40]
  wire  _GEN_7266 = unuse_way == 2'h2 ? _GEN_2773 : _GEN_6881; // @[d_cache.scala 125:40]
  wire  _GEN_7267 = unuse_way == 2'h2 ? _GEN_2774 : _GEN_6882; // @[d_cache.scala 125:40]
  wire  _GEN_7268 = unuse_way == 2'h2 ? _GEN_2775 : _GEN_6883; // @[d_cache.scala 125:40]
  wire  _GEN_7269 = unuse_way == 2'h2 ? _GEN_2776 : _GEN_6884; // @[d_cache.scala 125:40]
  wire  _GEN_7270 = unuse_way == 2'h2 ? _GEN_2777 : _GEN_6885; // @[d_cache.scala 125:40]
  wire  _GEN_7271 = unuse_way == 2'h2 ? _GEN_2778 : _GEN_6886; // @[d_cache.scala 125:40]
  wire  _GEN_7272 = unuse_way == 2'h2 ? _GEN_2779 : _GEN_6887; // @[d_cache.scala 125:40]
  wire  _GEN_7273 = unuse_way == 2'h2 ? _GEN_2780 : _GEN_6888; // @[d_cache.scala 125:40]
  wire  _GEN_7274 = unuse_way == 2'h2 ? _GEN_2781 : _GEN_6889; // @[d_cache.scala 125:40]
  wire  _GEN_7275 = unuse_way == 2'h2 ? _GEN_2782 : _GEN_6890; // @[d_cache.scala 125:40]
  wire  _GEN_7276 = unuse_way == 2'h2 ? _GEN_2783 : _GEN_6891; // @[d_cache.scala 125:40]
  wire  _GEN_7277 = unuse_way == 2'h2 ? _GEN_2784 : _GEN_6892; // @[d_cache.scala 125:40]
  wire  _GEN_7278 = unuse_way == 2'h2 ? _GEN_2785 : _GEN_6893; // @[d_cache.scala 125:40]
  wire  _GEN_7279 = unuse_way == 2'h2 ? _GEN_2786 : _GEN_6894; // @[d_cache.scala 125:40]
  wire  _GEN_7280 = unuse_way == 2'h2 ? _GEN_2787 : _GEN_6895; // @[d_cache.scala 125:40]
  wire  _GEN_7281 = unuse_way == 2'h2 ? _GEN_2788 : _GEN_6896; // @[d_cache.scala 125:40]
  wire  _GEN_7282 = unuse_way == 2'h2 ? _GEN_2789 : _GEN_6897; // @[d_cache.scala 125:40]
  wire  _GEN_7283 = unuse_way == 2'h2 ? _GEN_2790 : _GEN_6898; // @[d_cache.scala 125:40]
  wire  _GEN_7284 = unuse_way == 2'h2 ? _GEN_2791 : _GEN_6899; // @[d_cache.scala 125:40]
  wire  _GEN_7285 = unuse_way == 2'h2 ? _GEN_2792 : _GEN_6900; // @[d_cache.scala 125:40]
  wire  _GEN_7286 = unuse_way == 2'h2 ? _GEN_2793 : _GEN_6901; // @[d_cache.scala 125:40]
  wire  _GEN_7287 = unuse_way == 2'h2 ? _GEN_2794 : _GEN_6902; // @[d_cache.scala 125:40]
  wire  _GEN_7288 = unuse_way == 2'h2 ? _GEN_2795 : _GEN_6903; // @[d_cache.scala 125:40]
  wire  _GEN_7289 = unuse_way == 2'h2 ? _GEN_2796 : _GEN_6904; // @[d_cache.scala 125:40]
  wire  _GEN_7290 = unuse_way == 2'h2 ? _GEN_2797 : _GEN_6905; // @[d_cache.scala 125:40]
  wire  _GEN_7291 = unuse_way == 2'h2 ? _GEN_2798 : _GEN_6906; // @[d_cache.scala 125:40]
  wire  _GEN_7292 = unuse_way == 2'h2 ? _GEN_2799 : _GEN_6907; // @[d_cache.scala 125:40]
  wire  _GEN_7293 = unuse_way == 2'h2 ? _GEN_2800 : _GEN_6908; // @[d_cache.scala 125:40]
  wire  _GEN_7294 = unuse_way == 2'h2 ? _GEN_2801 : _GEN_6909; // @[d_cache.scala 125:40]
  wire  _GEN_7295 = unuse_way == 2'h2 ? _GEN_2802 : _GEN_6910; // @[d_cache.scala 125:40]
  wire  _GEN_7296 = unuse_way == 2'h2 ? _GEN_2803 : _GEN_6911; // @[d_cache.scala 125:40]
  wire  _GEN_7297 = unuse_way == 2'h2 ? _GEN_2804 : _GEN_6912; // @[d_cache.scala 125:40]
  wire  _GEN_7298 = unuse_way == 2'h2 ? _GEN_2805 : _GEN_6913; // @[d_cache.scala 125:40]
  wire  _GEN_7299 = unuse_way == 2'h2 ? _GEN_2806 : _GEN_6914; // @[d_cache.scala 125:40]
  wire  _GEN_7300 = unuse_way == 2'h2 ? _GEN_2807 : _GEN_6915; // @[d_cache.scala 125:40]
  wire  _GEN_7301 = unuse_way == 2'h2 ? _GEN_2808 : _GEN_6916; // @[d_cache.scala 125:40]
  wire  _GEN_7302 = unuse_way == 2'h2 ? _GEN_2809 : _GEN_6917; // @[d_cache.scala 125:40]
  wire  _GEN_7303 = unuse_way == 2'h2 ? _GEN_2810 : _GEN_6918; // @[d_cache.scala 125:40]
  wire  _GEN_7304 = unuse_way == 2'h2 ? _GEN_2811 : _GEN_6919; // @[d_cache.scala 125:40]
  wire  _GEN_7305 = unuse_way == 2'h2 ? _GEN_2812 : _GEN_6920; // @[d_cache.scala 125:40]
  wire  _GEN_7306 = unuse_way == 2'h2 ? _GEN_2813 : _GEN_6921; // @[d_cache.scala 125:40]
  wire  _GEN_7307 = unuse_way == 2'h2 ? _GEN_2814 : _GEN_6922; // @[d_cache.scala 125:40]
  wire  _GEN_7308 = unuse_way == 2'h2 ? _GEN_2815 : _GEN_6923; // @[d_cache.scala 125:40]
  wire  _GEN_7309 = unuse_way == 2'h2 ? _GEN_2816 : _GEN_6924; // @[d_cache.scala 125:40]
  wire  _GEN_7310 = unuse_way == 2'h2 ? _GEN_2817 : _GEN_6925; // @[d_cache.scala 125:40]
  wire  _GEN_7311 = unuse_way == 2'h2 ? _GEN_2818 : _GEN_6926; // @[d_cache.scala 125:40]
  wire  _GEN_7312 = unuse_way == 2'h2 ? _GEN_2819 : _GEN_6927; // @[d_cache.scala 125:40]
  wire  _GEN_7313 = unuse_way == 2'h2 ? _GEN_2820 : _GEN_6928; // @[d_cache.scala 125:40]
  wire  _GEN_7314 = unuse_way == 2'h2 ? _GEN_2821 : _GEN_6929; // @[d_cache.scala 125:40]
  wire  _GEN_7315 = unuse_way == 2'h2 ? _GEN_2822 : _GEN_6930; // @[d_cache.scala 125:40]
  wire  _GEN_7316 = unuse_way == 2'h2 ? _GEN_2823 : _GEN_6931; // @[d_cache.scala 125:40]
  wire  _GEN_7317 = unuse_way == 2'h2 ? _GEN_2824 : _GEN_6932; // @[d_cache.scala 125:40]
  wire  _GEN_7318 = unuse_way == 2'h2 ? _GEN_2825 : _GEN_6933; // @[d_cache.scala 125:40]
  wire  _GEN_7319 = unuse_way == 2'h2 ? _GEN_2826 : _GEN_6934; // @[d_cache.scala 125:40]
  wire  _GEN_7320 = unuse_way == 2'h2 ? _GEN_2827 : _GEN_6935; // @[d_cache.scala 125:40]
  wire  _GEN_7321 = unuse_way == 2'h2 ? _GEN_2828 : _GEN_6936; // @[d_cache.scala 125:40]
  wire  _GEN_7322 = unuse_way == 2'h2 ? _GEN_2829 : _GEN_6937; // @[d_cache.scala 125:40]
  wire  _GEN_7323 = unuse_way == 2'h2 ? 1'h0 : _T_28; // @[d_cache.scala 125:40 130:23]
  wire [63:0] _GEN_7324 = unuse_way == 2'h2 ? write_back_data : _GEN_5910; // @[d_cache.scala 125:40 29:34]
  wire [38:0] _GEN_7325 = unuse_way == 2'h2 ? {{7'd0}, write_back_addr} : _GEN_5911; // @[d_cache.scala 125:40 30:34]
  wire [63:0] _GEN_7326 = unuse_way == 2'h2 ? ram_0_0 : _GEN_5912; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7327 = unuse_way == 2'h2 ? ram_0_1 : _GEN_5913; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7328 = unuse_way == 2'h2 ? ram_0_2 : _GEN_5914; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7329 = unuse_way == 2'h2 ? ram_0_3 : _GEN_5915; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7330 = unuse_way == 2'h2 ? ram_0_4 : _GEN_5916; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7331 = unuse_way == 2'h2 ? ram_0_5 : _GEN_5917; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7332 = unuse_way == 2'h2 ? ram_0_6 : _GEN_5918; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7333 = unuse_way == 2'h2 ? ram_0_7 : _GEN_5919; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7334 = unuse_way == 2'h2 ? ram_0_8 : _GEN_5920; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7335 = unuse_way == 2'h2 ? ram_0_9 : _GEN_5921; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7336 = unuse_way == 2'h2 ? ram_0_10 : _GEN_5922; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7337 = unuse_way == 2'h2 ? ram_0_11 : _GEN_5923; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7338 = unuse_way == 2'h2 ? ram_0_12 : _GEN_5924; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7339 = unuse_way == 2'h2 ? ram_0_13 : _GEN_5925; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7340 = unuse_way == 2'h2 ? ram_0_14 : _GEN_5926; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7341 = unuse_way == 2'h2 ? ram_0_15 : _GEN_5927; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7342 = unuse_way == 2'h2 ? ram_0_16 : _GEN_5928; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7343 = unuse_way == 2'h2 ? ram_0_17 : _GEN_5929; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7344 = unuse_way == 2'h2 ? ram_0_18 : _GEN_5930; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7345 = unuse_way == 2'h2 ? ram_0_19 : _GEN_5931; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7346 = unuse_way == 2'h2 ? ram_0_20 : _GEN_5932; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7347 = unuse_way == 2'h2 ? ram_0_21 : _GEN_5933; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7348 = unuse_way == 2'h2 ? ram_0_22 : _GEN_5934; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7349 = unuse_way == 2'h2 ? ram_0_23 : _GEN_5935; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7350 = unuse_way == 2'h2 ? ram_0_24 : _GEN_5936; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7351 = unuse_way == 2'h2 ? ram_0_25 : _GEN_5937; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7352 = unuse_way == 2'h2 ? ram_0_26 : _GEN_5938; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7353 = unuse_way == 2'h2 ? ram_0_27 : _GEN_5939; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7354 = unuse_way == 2'h2 ? ram_0_28 : _GEN_5940; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7355 = unuse_way == 2'h2 ? ram_0_29 : _GEN_5941; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7356 = unuse_way == 2'h2 ? ram_0_30 : _GEN_5942; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7357 = unuse_way == 2'h2 ? ram_0_31 : _GEN_5943; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7358 = unuse_way == 2'h2 ? ram_0_32 : _GEN_5944; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7359 = unuse_way == 2'h2 ? ram_0_33 : _GEN_5945; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7360 = unuse_way == 2'h2 ? ram_0_34 : _GEN_5946; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7361 = unuse_way == 2'h2 ? ram_0_35 : _GEN_5947; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7362 = unuse_way == 2'h2 ? ram_0_36 : _GEN_5948; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7363 = unuse_way == 2'h2 ? ram_0_37 : _GEN_5949; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7364 = unuse_way == 2'h2 ? ram_0_38 : _GEN_5950; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7365 = unuse_way == 2'h2 ? ram_0_39 : _GEN_5951; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7366 = unuse_way == 2'h2 ? ram_0_40 : _GEN_5952; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7367 = unuse_way == 2'h2 ? ram_0_41 : _GEN_5953; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7368 = unuse_way == 2'h2 ? ram_0_42 : _GEN_5954; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7369 = unuse_way == 2'h2 ? ram_0_43 : _GEN_5955; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7370 = unuse_way == 2'h2 ? ram_0_44 : _GEN_5956; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7371 = unuse_way == 2'h2 ? ram_0_45 : _GEN_5957; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7372 = unuse_way == 2'h2 ? ram_0_46 : _GEN_5958; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7373 = unuse_way == 2'h2 ? ram_0_47 : _GEN_5959; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7374 = unuse_way == 2'h2 ? ram_0_48 : _GEN_5960; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7375 = unuse_way == 2'h2 ? ram_0_49 : _GEN_5961; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7376 = unuse_way == 2'h2 ? ram_0_50 : _GEN_5962; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7377 = unuse_way == 2'h2 ? ram_0_51 : _GEN_5963; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7378 = unuse_way == 2'h2 ? ram_0_52 : _GEN_5964; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7379 = unuse_way == 2'h2 ? ram_0_53 : _GEN_5965; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7380 = unuse_way == 2'h2 ? ram_0_54 : _GEN_5966; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7381 = unuse_way == 2'h2 ? ram_0_55 : _GEN_5967; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7382 = unuse_way == 2'h2 ? ram_0_56 : _GEN_5968; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7383 = unuse_way == 2'h2 ? ram_0_57 : _GEN_5969; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7384 = unuse_way == 2'h2 ? ram_0_58 : _GEN_5970; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7385 = unuse_way == 2'h2 ? ram_0_59 : _GEN_5971; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7386 = unuse_way == 2'h2 ? ram_0_60 : _GEN_5972; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7387 = unuse_way == 2'h2 ? ram_0_61 : _GEN_5973; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7388 = unuse_way == 2'h2 ? ram_0_62 : _GEN_5974; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7389 = unuse_way == 2'h2 ? ram_0_63 : _GEN_5975; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7390 = unuse_way == 2'h2 ? ram_0_64 : _GEN_5976; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7391 = unuse_way == 2'h2 ? ram_0_65 : _GEN_5977; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7392 = unuse_way == 2'h2 ? ram_0_66 : _GEN_5978; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7393 = unuse_way == 2'h2 ? ram_0_67 : _GEN_5979; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7394 = unuse_way == 2'h2 ? ram_0_68 : _GEN_5980; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7395 = unuse_way == 2'h2 ? ram_0_69 : _GEN_5981; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7396 = unuse_way == 2'h2 ? ram_0_70 : _GEN_5982; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7397 = unuse_way == 2'h2 ? ram_0_71 : _GEN_5983; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7398 = unuse_way == 2'h2 ? ram_0_72 : _GEN_5984; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7399 = unuse_way == 2'h2 ? ram_0_73 : _GEN_5985; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7400 = unuse_way == 2'h2 ? ram_0_74 : _GEN_5986; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7401 = unuse_way == 2'h2 ? ram_0_75 : _GEN_5987; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7402 = unuse_way == 2'h2 ? ram_0_76 : _GEN_5988; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7403 = unuse_way == 2'h2 ? ram_0_77 : _GEN_5989; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7404 = unuse_way == 2'h2 ? ram_0_78 : _GEN_5990; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7405 = unuse_way == 2'h2 ? ram_0_79 : _GEN_5991; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7406 = unuse_way == 2'h2 ? ram_0_80 : _GEN_5992; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7407 = unuse_way == 2'h2 ? ram_0_81 : _GEN_5993; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7408 = unuse_way == 2'h2 ? ram_0_82 : _GEN_5994; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7409 = unuse_way == 2'h2 ? ram_0_83 : _GEN_5995; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7410 = unuse_way == 2'h2 ? ram_0_84 : _GEN_5996; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7411 = unuse_way == 2'h2 ? ram_0_85 : _GEN_5997; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7412 = unuse_way == 2'h2 ? ram_0_86 : _GEN_5998; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7413 = unuse_way == 2'h2 ? ram_0_87 : _GEN_5999; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7414 = unuse_way == 2'h2 ? ram_0_88 : _GEN_6000; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7415 = unuse_way == 2'h2 ? ram_0_89 : _GEN_6001; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7416 = unuse_way == 2'h2 ? ram_0_90 : _GEN_6002; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7417 = unuse_way == 2'h2 ? ram_0_91 : _GEN_6003; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7418 = unuse_way == 2'h2 ? ram_0_92 : _GEN_6004; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7419 = unuse_way == 2'h2 ? ram_0_93 : _GEN_6005; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7420 = unuse_way == 2'h2 ? ram_0_94 : _GEN_6006; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7421 = unuse_way == 2'h2 ? ram_0_95 : _GEN_6007; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7422 = unuse_way == 2'h2 ? ram_0_96 : _GEN_6008; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7423 = unuse_way == 2'h2 ? ram_0_97 : _GEN_6009; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7424 = unuse_way == 2'h2 ? ram_0_98 : _GEN_6010; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7425 = unuse_way == 2'h2 ? ram_0_99 : _GEN_6011; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7426 = unuse_way == 2'h2 ? ram_0_100 : _GEN_6012; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7427 = unuse_way == 2'h2 ? ram_0_101 : _GEN_6013; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7428 = unuse_way == 2'h2 ? ram_0_102 : _GEN_6014; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7429 = unuse_way == 2'h2 ? ram_0_103 : _GEN_6015; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7430 = unuse_way == 2'h2 ? ram_0_104 : _GEN_6016; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7431 = unuse_way == 2'h2 ? ram_0_105 : _GEN_6017; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7432 = unuse_way == 2'h2 ? ram_0_106 : _GEN_6018; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7433 = unuse_way == 2'h2 ? ram_0_107 : _GEN_6019; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7434 = unuse_way == 2'h2 ? ram_0_108 : _GEN_6020; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7435 = unuse_way == 2'h2 ? ram_0_109 : _GEN_6021; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7436 = unuse_way == 2'h2 ? ram_0_110 : _GEN_6022; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7437 = unuse_way == 2'h2 ? ram_0_111 : _GEN_6023; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7438 = unuse_way == 2'h2 ? ram_0_112 : _GEN_6024; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7439 = unuse_way == 2'h2 ? ram_0_113 : _GEN_6025; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7440 = unuse_way == 2'h2 ? ram_0_114 : _GEN_6026; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7441 = unuse_way == 2'h2 ? ram_0_115 : _GEN_6027; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7442 = unuse_way == 2'h2 ? ram_0_116 : _GEN_6028; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7443 = unuse_way == 2'h2 ? ram_0_117 : _GEN_6029; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7444 = unuse_way == 2'h2 ? ram_0_118 : _GEN_6030; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7445 = unuse_way == 2'h2 ? ram_0_119 : _GEN_6031; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7446 = unuse_way == 2'h2 ? ram_0_120 : _GEN_6032; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7447 = unuse_way == 2'h2 ? ram_0_121 : _GEN_6033; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7448 = unuse_way == 2'h2 ? ram_0_122 : _GEN_6034; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7449 = unuse_way == 2'h2 ? ram_0_123 : _GEN_6035; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7450 = unuse_way == 2'h2 ? ram_0_124 : _GEN_6036; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7451 = unuse_way == 2'h2 ? ram_0_125 : _GEN_6037; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7452 = unuse_way == 2'h2 ? ram_0_126 : _GEN_6038; // @[d_cache.scala 125:40 18:24]
  wire [63:0] _GEN_7453 = unuse_way == 2'h2 ? ram_0_127 : _GEN_6039; // @[d_cache.scala 125:40 18:24]
  wire [31:0] _GEN_7454 = unuse_way == 2'h2 ? tag_0_0 : _GEN_6040; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7455 = unuse_way == 2'h2 ? tag_0_1 : _GEN_6041; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7456 = unuse_way == 2'h2 ? tag_0_2 : _GEN_6042; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7457 = unuse_way == 2'h2 ? tag_0_3 : _GEN_6043; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7458 = unuse_way == 2'h2 ? tag_0_4 : _GEN_6044; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7459 = unuse_way == 2'h2 ? tag_0_5 : _GEN_6045; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7460 = unuse_way == 2'h2 ? tag_0_6 : _GEN_6046; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7461 = unuse_way == 2'h2 ? tag_0_7 : _GEN_6047; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7462 = unuse_way == 2'h2 ? tag_0_8 : _GEN_6048; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7463 = unuse_way == 2'h2 ? tag_0_9 : _GEN_6049; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7464 = unuse_way == 2'h2 ? tag_0_10 : _GEN_6050; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7465 = unuse_way == 2'h2 ? tag_0_11 : _GEN_6051; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7466 = unuse_way == 2'h2 ? tag_0_12 : _GEN_6052; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7467 = unuse_way == 2'h2 ? tag_0_13 : _GEN_6053; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7468 = unuse_way == 2'h2 ? tag_0_14 : _GEN_6054; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7469 = unuse_way == 2'h2 ? tag_0_15 : _GEN_6055; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7470 = unuse_way == 2'h2 ? tag_0_16 : _GEN_6056; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7471 = unuse_way == 2'h2 ? tag_0_17 : _GEN_6057; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7472 = unuse_way == 2'h2 ? tag_0_18 : _GEN_6058; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7473 = unuse_way == 2'h2 ? tag_0_19 : _GEN_6059; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7474 = unuse_way == 2'h2 ? tag_0_20 : _GEN_6060; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7475 = unuse_way == 2'h2 ? tag_0_21 : _GEN_6061; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7476 = unuse_way == 2'h2 ? tag_0_22 : _GEN_6062; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7477 = unuse_way == 2'h2 ? tag_0_23 : _GEN_6063; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7478 = unuse_way == 2'h2 ? tag_0_24 : _GEN_6064; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7479 = unuse_way == 2'h2 ? tag_0_25 : _GEN_6065; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7480 = unuse_way == 2'h2 ? tag_0_26 : _GEN_6066; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7481 = unuse_way == 2'h2 ? tag_0_27 : _GEN_6067; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7482 = unuse_way == 2'h2 ? tag_0_28 : _GEN_6068; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7483 = unuse_way == 2'h2 ? tag_0_29 : _GEN_6069; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7484 = unuse_way == 2'h2 ? tag_0_30 : _GEN_6070; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7485 = unuse_way == 2'h2 ? tag_0_31 : _GEN_6071; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7486 = unuse_way == 2'h2 ? tag_0_32 : _GEN_6072; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7487 = unuse_way == 2'h2 ? tag_0_33 : _GEN_6073; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7488 = unuse_way == 2'h2 ? tag_0_34 : _GEN_6074; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7489 = unuse_way == 2'h2 ? tag_0_35 : _GEN_6075; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7490 = unuse_way == 2'h2 ? tag_0_36 : _GEN_6076; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7491 = unuse_way == 2'h2 ? tag_0_37 : _GEN_6077; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7492 = unuse_way == 2'h2 ? tag_0_38 : _GEN_6078; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7493 = unuse_way == 2'h2 ? tag_0_39 : _GEN_6079; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7494 = unuse_way == 2'h2 ? tag_0_40 : _GEN_6080; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7495 = unuse_way == 2'h2 ? tag_0_41 : _GEN_6081; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7496 = unuse_way == 2'h2 ? tag_0_42 : _GEN_6082; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7497 = unuse_way == 2'h2 ? tag_0_43 : _GEN_6083; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7498 = unuse_way == 2'h2 ? tag_0_44 : _GEN_6084; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7499 = unuse_way == 2'h2 ? tag_0_45 : _GEN_6085; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7500 = unuse_way == 2'h2 ? tag_0_46 : _GEN_6086; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7501 = unuse_way == 2'h2 ? tag_0_47 : _GEN_6087; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7502 = unuse_way == 2'h2 ? tag_0_48 : _GEN_6088; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7503 = unuse_way == 2'h2 ? tag_0_49 : _GEN_6089; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7504 = unuse_way == 2'h2 ? tag_0_50 : _GEN_6090; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7505 = unuse_way == 2'h2 ? tag_0_51 : _GEN_6091; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7506 = unuse_way == 2'h2 ? tag_0_52 : _GEN_6092; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7507 = unuse_way == 2'h2 ? tag_0_53 : _GEN_6093; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7508 = unuse_way == 2'h2 ? tag_0_54 : _GEN_6094; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7509 = unuse_way == 2'h2 ? tag_0_55 : _GEN_6095; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7510 = unuse_way == 2'h2 ? tag_0_56 : _GEN_6096; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7511 = unuse_way == 2'h2 ? tag_0_57 : _GEN_6097; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7512 = unuse_way == 2'h2 ? tag_0_58 : _GEN_6098; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7513 = unuse_way == 2'h2 ? tag_0_59 : _GEN_6099; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7514 = unuse_way == 2'h2 ? tag_0_60 : _GEN_6100; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7515 = unuse_way == 2'h2 ? tag_0_61 : _GEN_6101; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7516 = unuse_way == 2'h2 ? tag_0_62 : _GEN_6102; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7517 = unuse_way == 2'h2 ? tag_0_63 : _GEN_6103; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7518 = unuse_way == 2'h2 ? tag_0_64 : _GEN_6104; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7519 = unuse_way == 2'h2 ? tag_0_65 : _GEN_6105; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7520 = unuse_way == 2'h2 ? tag_0_66 : _GEN_6106; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7521 = unuse_way == 2'h2 ? tag_0_67 : _GEN_6107; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7522 = unuse_way == 2'h2 ? tag_0_68 : _GEN_6108; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7523 = unuse_way == 2'h2 ? tag_0_69 : _GEN_6109; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7524 = unuse_way == 2'h2 ? tag_0_70 : _GEN_6110; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7525 = unuse_way == 2'h2 ? tag_0_71 : _GEN_6111; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7526 = unuse_way == 2'h2 ? tag_0_72 : _GEN_6112; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7527 = unuse_way == 2'h2 ? tag_0_73 : _GEN_6113; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7528 = unuse_way == 2'h2 ? tag_0_74 : _GEN_6114; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7529 = unuse_way == 2'h2 ? tag_0_75 : _GEN_6115; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7530 = unuse_way == 2'h2 ? tag_0_76 : _GEN_6116; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7531 = unuse_way == 2'h2 ? tag_0_77 : _GEN_6117; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7532 = unuse_way == 2'h2 ? tag_0_78 : _GEN_6118; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7533 = unuse_way == 2'h2 ? tag_0_79 : _GEN_6119; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7534 = unuse_way == 2'h2 ? tag_0_80 : _GEN_6120; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7535 = unuse_way == 2'h2 ? tag_0_81 : _GEN_6121; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7536 = unuse_way == 2'h2 ? tag_0_82 : _GEN_6122; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7537 = unuse_way == 2'h2 ? tag_0_83 : _GEN_6123; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7538 = unuse_way == 2'h2 ? tag_0_84 : _GEN_6124; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7539 = unuse_way == 2'h2 ? tag_0_85 : _GEN_6125; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7540 = unuse_way == 2'h2 ? tag_0_86 : _GEN_6126; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7541 = unuse_way == 2'h2 ? tag_0_87 : _GEN_6127; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7542 = unuse_way == 2'h2 ? tag_0_88 : _GEN_6128; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7543 = unuse_way == 2'h2 ? tag_0_89 : _GEN_6129; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7544 = unuse_way == 2'h2 ? tag_0_90 : _GEN_6130; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7545 = unuse_way == 2'h2 ? tag_0_91 : _GEN_6131; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7546 = unuse_way == 2'h2 ? tag_0_92 : _GEN_6132; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7547 = unuse_way == 2'h2 ? tag_0_93 : _GEN_6133; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7548 = unuse_way == 2'h2 ? tag_0_94 : _GEN_6134; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7549 = unuse_way == 2'h2 ? tag_0_95 : _GEN_6135; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7550 = unuse_way == 2'h2 ? tag_0_96 : _GEN_6136; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7551 = unuse_way == 2'h2 ? tag_0_97 : _GEN_6137; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7552 = unuse_way == 2'h2 ? tag_0_98 : _GEN_6138; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7553 = unuse_way == 2'h2 ? tag_0_99 : _GEN_6139; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7554 = unuse_way == 2'h2 ? tag_0_100 : _GEN_6140; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7555 = unuse_way == 2'h2 ? tag_0_101 : _GEN_6141; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7556 = unuse_way == 2'h2 ? tag_0_102 : _GEN_6142; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7557 = unuse_way == 2'h2 ? tag_0_103 : _GEN_6143; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7558 = unuse_way == 2'h2 ? tag_0_104 : _GEN_6144; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7559 = unuse_way == 2'h2 ? tag_0_105 : _GEN_6145; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7560 = unuse_way == 2'h2 ? tag_0_106 : _GEN_6146; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7561 = unuse_way == 2'h2 ? tag_0_107 : _GEN_6147; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7562 = unuse_way == 2'h2 ? tag_0_108 : _GEN_6148; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7563 = unuse_way == 2'h2 ? tag_0_109 : _GEN_6149; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7564 = unuse_way == 2'h2 ? tag_0_110 : _GEN_6150; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7565 = unuse_way == 2'h2 ? tag_0_111 : _GEN_6151; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7566 = unuse_way == 2'h2 ? tag_0_112 : _GEN_6152; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7567 = unuse_way == 2'h2 ? tag_0_113 : _GEN_6153; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7568 = unuse_way == 2'h2 ? tag_0_114 : _GEN_6154; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7569 = unuse_way == 2'h2 ? tag_0_115 : _GEN_6155; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7570 = unuse_way == 2'h2 ? tag_0_116 : _GEN_6156; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7571 = unuse_way == 2'h2 ? tag_0_117 : _GEN_6157; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7572 = unuse_way == 2'h2 ? tag_0_118 : _GEN_6158; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7573 = unuse_way == 2'h2 ? tag_0_119 : _GEN_6159; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7574 = unuse_way == 2'h2 ? tag_0_120 : _GEN_6160; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7575 = unuse_way == 2'h2 ? tag_0_121 : _GEN_6161; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7576 = unuse_way == 2'h2 ? tag_0_122 : _GEN_6162; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7577 = unuse_way == 2'h2 ? tag_0_123 : _GEN_6163; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7578 = unuse_way == 2'h2 ? tag_0_124 : _GEN_6164; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7579 = unuse_way == 2'h2 ? tag_0_125 : _GEN_6165; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7580 = unuse_way == 2'h2 ? tag_0_126 : _GEN_6166; // @[d_cache.scala 125:40 20:24]
  wire [31:0] _GEN_7581 = unuse_way == 2'h2 ? tag_0_127 : _GEN_6167; // @[d_cache.scala 125:40 20:24]
  wire  _GEN_7582 = unuse_way == 2'h2 ? dirty_0_0 : _GEN_6168; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7583 = unuse_way == 2'h2 ? dirty_0_1 : _GEN_6169; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7584 = unuse_way == 2'h2 ? dirty_0_2 : _GEN_6170; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7585 = unuse_way == 2'h2 ? dirty_0_3 : _GEN_6171; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7586 = unuse_way == 2'h2 ? dirty_0_4 : _GEN_6172; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7587 = unuse_way == 2'h2 ? dirty_0_5 : _GEN_6173; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7588 = unuse_way == 2'h2 ? dirty_0_6 : _GEN_6174; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7589 = unuse_way == 2'h2 ? dirty_0_7 : _GEN_6175; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7590 = unuse_way == 2'h2 ? dirty_0_8 : _GEN_6176; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7591 = unuse_way == 2'h2 ? dirty_0_9 : _GEN_6177; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7592 = unuse_way == 2'h2 ? dirty_0_10 : _GEN_6178; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7593 = unuse_way == 2'h2 ? dirty_0_11 : _GEN_6179; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7594 = unuse_way == 2'h2 ? dirty_0_12 : _GEN_6180; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7595 = unuse_way == 2'h2 ? dirty_0_13 : _GEN_6181; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7596 = unuse_way == 2'h2 ? dirty_0_14 : _GEN_6182; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7597 = unuse_way == 2'h2 ? dirty_0_15 : _GEN_6183; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7598 = unuse_way == 2'h2 ? dirty_0_16 : _GEN_6184; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7599 = unuse_way == 2'h2 ? dirty_0_17 : _GEN_6185; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7600 = unuse_way == 2'h2 ? dirty_0_18 : _GEN_6186; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7601 = unuse_way == 2'h2 ? dirty_0_19 : _GEN_6187; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7602 = unuse_way == 2'h2 ? dirty_0_20 : _GEN_6188; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7603 = unuse_way == 2'h2 ? dirty_0_21 : _GEN_6189; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7604 = unuse_way == 2'h2 ? dirty_0_22 : _GEN_6190; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7605 = unuse_way == 2'h2 ? dirty_0_23 : _GEN_6191; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7606 = unuse_way == 2'h2 ? dirty_0_24 : _GEN_6192; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7607 = unuse_way == 2'h2 ? dirty_0_25 : _GEN_6193; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7608 = unuse_way == 2'h2 ? dirty_0_26 : _GEN_6194; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7609 = unuse_way == 2'h2 ? dirty_0_27 : _GEN_6195; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7610 = unuse_way == 2'h2 ? dirty_0_28 : _GEN_6196; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7611 = unuse_way == 2'h2 ? dirty_0_29 : _GEN_6197; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7612 = unuse_way == 2'h2 ? dirty_0_30 : _GEN_6198; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7613 = unuse_way == 2'h2 ? dirty_0_31 : _GEN_6199; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7614 = unuse_way == 2'h2 ? dirty_0_32 : _GEN_6200; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7615 = unuse_way == 2'h2 ? dirty_0_33 : _GEN_6201; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7616 = unuse_way == 2'h2 ? dirty_0_34 : _GEN_6202; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7617 = unuse_way == 2'h2 ? dirty_0_35 : _GEN_6203; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7618 = unuse_way == 2'h2 ? dirty_0_36 : _GEN_6204; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7619 = unuse_way == 2'h2 ? dirty_0_37 : _GEN_6205; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7620 = unuse_way == 2'h2 ? dirty_0_38 : _GEN_6206; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7621 = unuse_way == 2'h2 ? dirty_0_39 : _GEN_6207; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7622 = unuse_way == 2'h2 ? dirty_0_40 : _GEN_6208; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7623 = unuse_way == 2'h2 ? dirty_0_41 : _GEN_6209; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7624 = unuse_way == 2'h2 ? dirty_0_42 : _GEN_6210; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7625 = unuse_way == 2'h2 ? dirty_0_43 : _GEN_6211; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7626 = unuse_way == 2'h2 ? dirty_0_44 : _GEN_6212; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7627 = unuse_way == 2'h2 ? dirty_0_45 : _GEN_6213; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7628 = unuse_way == 2'h2 ? dirty_0_46 : _GEN_6214; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7629 = unuse_way == 2'h2 ? dirty_0_47 : _GEN_6215; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7630 = unuse_way == 2'h2 ? dirty_0_48 : _GEN_6216; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7631 = unuse_way == 2'h2 ? dirty_0_49 : _GEN_6217; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7632 = unuse_way == 2'h2 ? dirty_0_50 : _GEN_6218; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7633 = unuse_way == 2'h2 ? dirty_0_51 : _GEN_6219; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7634 = unuse_way == 2'h2 ? dirty_0_52 : _GEN_6220; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7635 = unuse_way == 2'h2 ? dirty_0_53 : _GEN_6221; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7636 = unuse_way == 2'h2 ? dirty_0_54 : _GEN_6222; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7637 = unuse_way == 2'h2 ? dirty_0_55 : _GEN_6223; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7638 = unuse_way == 2'h2 ? dirty_0_56 : _GEN_6224; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7639 = unuse_way == 2'h2 ? dirty_0_57 : _GEN_6225; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7640 = unuse_way == 2'h2 ? dirty_0_58 : _GEN_6226; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7641 = unuse_way == 2'h2 ? dirty_0_59 : _GEN_6227; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7642 = unuse_way == 2'h2 ? dirty_0_60 : _GEN_6228; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7643 = unuse_way == 2'h2 ? dirty_0_61 : _GEN_6229; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7644 = unuse_way == 2'h2 ? dirty_0_62 : _GEN_6230; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7645 = unuse_way == 2'h2 ? dirty_0_63 : _GEN_6231; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7646 = unuse_way == 2'h2 ? dirty_0_64 : _GEN_6232; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7647 = unuse_way == 2'h2 ? dirty_0_65 : _GEN_6233; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7648 = unuse_way == 2'h2 ? dirty_0_66 : _GEN_6234; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7649 = unuse_way == 2'h2 ? dirty_0_67 : _GEN_6235; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7650 = unuse_way == 2'h2 ? dirty_0_68 : _GEN_6236; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7651 = unuse_way == 2'h2 ? dirty_0_69 : _GEN_6237; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7652 = unuse_way == 2'h2 ? dirty_0_70 : _GEN_6238; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7653 = unuse_way == 2'h2 ? dirty_0_71 : _GEN_6239; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7654 = unuse_way == 2'h2 ? dirty_0_72 : _GEN_6240; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7655 = unuse_way == 2'h2 ? dirty_0_73 : _GEN_6241; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7656 = unuse_way == 2'h2 ? dirty_0_74 : _GEN_6242; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7657 = unuse_way == 2'h2 ? dirty_0_75 : _GEN_6243; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7658 = unuse_way == 2'h2 ? dirty_0_76 : _GEN_6244; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7659 = unuse_way == 2'h2 ? dirty_0_77 : _GEN_6245; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7660 = unuse_way == 2'h2 ? dirty_0_78 : _GEN_6246; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7661 = unuse_way == 2'h2 ? dirty_0_79 : _GEN_6247; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7662 = unuse_way == 2'h2 ? dirty_0_80 : _GEN_6248; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7663 = unuse_way == 2'h2 ? dirty_0_81 : _GEN_6249; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7664 = unuse_way == 2'h2 ? dirty_0_82 : _GEN_6250; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7665 = unuse_way == 2'h2 ? dirty_0_83 : _GEN_6251; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7666 = unuse_way == 2'h2 ? dirty_0_84 : _GEN_6252; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7667 = unuse_way == 2'h2 ? dirty_0_85 : _GEN_6253; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7668 = unuse_way == 2'h2 ? dirty_0_86 : _GEN_6254; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7669 = unuse_way == 2'h2 ? dirty_0_87 : _GEN_6255; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7670 = unuse_way == 2'h2 ? dirty_0_88 : _GEN_6256; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7671 = unuse_way == 2'h2 ? dirty_0_89 : _GEN_6257; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7672 = unuse_way == 2'h2 ? dirty_0_90 : _GEN_6258; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7673 = unuse_way == 2'h2 ? dirty_0_91 : _GEN_6259; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7674 = unuse_way == 2'h2 ? dirty_0_92 : _GEN_6260; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7675 = unuse_way == 2'h2 ? dirty_0_93 : _GEN_6261; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7676 = unuse_way == 2'h2 ? dirty_0_94 : _GEN_6262; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7677 = unuse_way == 2'h2 ? dirty_0_95 : _GEN_6263; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7678 = unuse_way == 2'h2 ? dirty_0_96 : _GEN_6264; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7679 = unuse_way == 2'h2 ? dirty_0_97 : _GEN_6265; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7680 = unuse_way == 2'h2 ? dirty_0_98 : _GEN_6266; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7681 = unuse_way == 2'h2 ? dirty_0_99 : _GEN_6267; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7682 = unuse_way == 2'h2 ? dirty_0_100 : _GEN_6268; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7683 = unuse_way == 2'h2 ? dirty_0_101 : _GEN_6269; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7684 = unuse_way == 2'h2 ? dirty_0_102 : _GEN_6270; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7685 = unuse_way == 2'h2 ? dirty_0_103 : _GEN_6271; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7686 = unuse_way == 2'h2 ? dirty_0_104 : _GEN_6272; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7687 = unuse_way == 2'h2 ? dirty_0_105 : _GEN_6273; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7688 = unuse_way == 2'h2 ? dirty_0_106 : _GEN_6274; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7689 = unuse_way == 2'h2 ? dirty_0_107 : _GEN_6275; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7690 = unuse_way == 2'h2 ? dirty_0_108 : _GEN_6276; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7691 = unuse_way == 2'h2 ? dirty_0_109 : _GEN_6277; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7692 = unuse_way == 2'h2 ? dirty_0_110 : _GEN_6278; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7693 = unuse_way == 2'h2 ? dirty_0_111 : _GEN_6279; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7694 = unuse_way == 2'h2 ? dirty_0_112 : _GEN_6280; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7695 = unuse_way == 2'h2 ? dirty_0_113 : _GEN_6281; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7696 = unuse_way == 2'h2 ? dirty_0_114 : _GEN_6282; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7697 = unuse_way == 2'h2 ? dirty_0_115 : _GEN_6283; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7698 = unuse_way == 2'h2 ? dirty_0_116 : _GEN_6284; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7699 = unuse_way == 2'h2 ? dirty_0_117 : _GEN_6285; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7700 = unuse_way == 2'h2 ? dirty_0_118 : _GEN_6286; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7701 = unuse_way == 2'h2 ? dirty_0_119 : _GEN_6287; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7702 = unuse_way == 2'h2 ? dirty_0_120 : _GEN_6288; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7703 = unuse_way == 2'h2 ? dirty_0_121 : _GEN_6289; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7704 = unuse_way == 2'h2 ? dirty_0_122 : _GEN_6290; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7705 = unuse_way == 2'h2 ? dirty_0_123 : _GEN_6291; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7706 = unuse_way == 2'h2 ? dirty_0_124 : _GEN_6292; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7707 = unuse_way == 2'h2 ? dirty_0_125 : _GEN_6293; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7708 = unuse_way == 2'h2 ? dirty_0_126 : _GEN_6294; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7709 = unuse_way == 2'h2 ? dirty_0_127 : _GEN_6295; // @[d_cache.scala 125:40 24:26]
  wire  _GEN_7710 = unuse_way == 2'h2 ? valid_0_0 : _GEN_6296; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7711 = unuse_way == 2'h2 ? valid_0_1 : _GEN_6297; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7712 = unuse_way == 2'h2 ? valid_0_2 : _GEN_6298; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7713 = unuse_way == 2'h2 ? valid_0_3 : _GEN_6299; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7714 = unuse_way == 2'h2 ? valid_0_4 : _GEN_6300; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7715 = unuse_way == 2'h2 ? valid_0_5 : _GEN_6301; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7716 = unuse_way == 2'h2 ? valid_0_6 : _GEN_6302; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7717 = unuse_way == 2'h2 ? valid_0_7 : _GEN_6303; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7718 = unuse_way == 2'h2 ? valid_0_8 : _GEN_6304; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7719 = unuse_way == 2'h2 ? valid_0_9 : _GEN_6305; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7720 = unuse_way == 2'h2 ? valid_0_10 : _GEN_6306; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7721 = unuse_way == 2'h2 ? valid_0_11 : _GEN_6307; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7722 = unuse_way == 2'h2 ? valid_0_12 : _GEN_6308; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7723 = unuse_way == 2'h2 ? valid_0_13 : _GEN_6309; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7724 = unuse_way == 2'h2 ? valid_0_14 : _GEN_6310; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7725 = unuse_way == 2'h2 ? valid_0_15 : _GEN_6311; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7726 = unuse_way == 2'h2 ? valid_0_16 : _GEN_6312; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7727 = unuse_way == 2'h2 ? valid_0_17 : _GEN_6313; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7728 = unuse_way == 2'h2 ? valid_0_18 : _GEN_6314; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7729 = unuse_way == 2'h2 ? valid_0_19 : _GEN_6315; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7730 = unuse_way == 2'h2 ? valid_0_20 : _GEN_6316; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7731 = unuse_way == 2'h2 ? valid_0_21 : _GEN_6317; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7732 = unuse_way == 2'h2 ? valid_0_22 : _GEN_6318; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7733 = unuse_way == 2'h2 ? valid_0_23 : _GEN_6319; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7734 = unuse_way == 2'h2 ? valid_0_24 : _GEN_6320; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7735 = unuse_way == 2'h2 ? valid_0_25 : _GEN_6321; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7736 = unuse_way == 2'h2 ? valid_0_26 : _GEN_6322; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7737 = unuse_way == 2'h2 ? valid_0_27 : _GEN_6323; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7738 = unuse_way == 2'h2 ? valid_0_28 : _GEN_6324; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7739 = unuse_way == 2'h2 ? valid_0_29 : _GEN_6325; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7740 = unuse_way == 2'h2 ? valid_0_30 : _GEN_6326; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7741 = unuse_way == 2'h2 ? valid_0_31 : _GEN_6327; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7742 = unuse_way == 2'h2 ? valid_0_32 : _GEN_6328; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7743 = unuse_way == 2'h2 ? valid_0_33 : _GEN_6329; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7744 = unuse_way == 2'h2 ? valid_0_34 : _GEN_6330; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7745 = unuse_way == 2'h2 ? valid_0_35 : _GEN_6331; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7746 = unuse_way == 2'h2 ? valid_0_36 : _GEN_6332; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7747 = unuse_way == 2'h2 ? valid_0_37 : _GEN_6333; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7748 = unuse_way == 2'h2 ? valid_0_38 : _GEN_6334; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7749 = unuse_way == 2'h2 ? valid_0_39 : _GEN_6335; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7750 = unuse_way == 2'h2 ? valid_0_40 : _GEN_6336; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7751 = unuse_way == 2'h2 ? valid_0_41 : _GEN_6337; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7752 = unuse_way == 2'h2 ? valid_0_42 : _GEN_6338; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7753 = unuse_way == 2'h2 ? valid_0_43 : _GEN_6339; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7754 = unuse_way == 2'h2 ? valid_0_44 : _GEN_6340; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7755 = unuse_way == 2'h2 ? valid_0_45 : _GEN_6341; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7756 = unuse_way == 2'h2 ? valid_0_46 : _GEN_6342; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7757 = unuse_way == 2'h2 ? valid_0_47 : _GEN_6343; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7758 = unuse_way == 2'h2 ? valid_0_48 : _GEN_6344; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7759 = unuse_way == 2'h2 ? valid_0_49 : _GEN_6345; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7760 = unuse_way == 2'h2 ? valid_0_50 : _GEN_6346; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7761 = unuse_way == 2'h2 ? valid_0_51 : _GEN_6347; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7762 = unuse_way == 2'h2 ? valid_0_52 : _GEN_6348; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7763 = unuse_way == 2'h2 ? valid_0_53 : _GEN_6349; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7764 = unuse_way == 2'h2 ? valid_0_54 : _GEN_6350; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7765 = unuse_way == 2'h2 ? valid_0_55 : _GEN_6351; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7766 = unuse_way == 2'h2 ? valid_0_56 : _GEN_6352; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7767 = unuse_way == 2'h2 ? valid_0_57 : _GEN_6353; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7768 = unuse_way == 2'h2 ? valid_0_58 : _GEN_6354; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7769 = unuse_way == 2'h2 ? valid_0_59 : _GEN_6355; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7770 = unuse_way == 2'h2 ? valid_0_60 : _GEN_6356; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7771 = unuse_way == 2'h2 ? valid_0_61 : _GEN_6357; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7772 = unuse_way == 2'h2 ? valid_0_62 : _GEN_6358; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7773 = unuse_way == 2'h2 ? valid_0_63 : _GEN_6359; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7774 = unuse_way == 2'h2 ? valid_0_64 : _GEN_6360; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7775 = unuse_way == 2'h2 ? valid_0_65 : _GEN_6361; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7776 = unuse_way == 2'h2 ? valid_0_66 : _GEN_6362; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7777 = unuse_way == 2'h2 ? valid_0_67 : _GEN_6363; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7778 = unuse_way == 2'h2 ? valid_0_68 : _GEN_6364; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7779 = unuse_way == 2'h2 ? valid_0_69 : _GEN_6365; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7780 = unuse_way == 2'h2 ? valid_0_70 : _GEN_6366; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7781 = unuse_way == 2'h2 ? valid_0_71 : _GEN_6367; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7782 = unuse_way == 2'h2 ? valid_0_72 : _GEN_6368; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7783 = unuse_way == 2'h2 ? valid_0_73 : _GEN_6369; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7784 = unuse_way == 2'h2 ? valid_0_74 : _GEN_6370; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7785 = unuse_way == 2'h2 ? valid_0_75 : _GEN_6371; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7786 = unuse_way == 2'h2 ? valid_0_76 : _GEN_6372; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7787 = unuse_way == 2'h2 ? valid_0_77 : _GEN_6373; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7788 = unuse_way == 2'h2 ? valid_0_78 : _GEN_6374; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7789 = unuse_way == 2'h2 ? valid_0_79 : _GEN_6375; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7790 = unuse_way == 2'h2 ? valid_0_80 : _GEN_6376; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7791 = unuse_way == 2'h2 ? valid_0_81 : _GEN_6377; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7792 = unuse_way == 2'h2 ? valid_0_82 : _GEN_6378; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7793 = unuse_way == 2'h2 ? valid_0_83 : _GEN_6379; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7794 = unuse_way == 2'h2 ? valid_0_84 : _GEN_6380; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7795 = unuse_way == 2'h2 ? valid_0_85 : _GEN_6381; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7796 = unuse_way == 2'h2 ? valid_0_86 : _GEN_6382; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7797 = unuse_way == 2'h2 ? valid_0_87 : _GEN_6383; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7798 = unuse_way == 2'h2 ? valid_0_88 : _GEN_6384; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7799 = unuse_way == 2'h2 ? valid_0_89 : _GEN_6385; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7800 = unuse_way == 2'h2 ? valid_0_90 : _GEN_6386; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7801 = unuse_way == 2'h2 ? valid_0_91 : _GEN_6387; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7802 = unuse_way == 2'h2 ? valid_0_92 : _GEN_6388; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7803 = unuse_way == 2'h2 ? valid_0_93 : _GEN_6389; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7804 = unuse_way == 2'h2 ? valid_0_94 : _GEN_6390; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7805 = unuse_way == 2'h2 ? valid_0_95 : _GEN_6391; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7806 = unuse_way == 2'h2 ? valid_0_96 : _GEN_6392; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7807 = unuse_way == 2'h2 ? valid_0_97 : _GEN_6393; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7808 = unuse_way == 2'h2 ? valid_0_98 : _GEN_6394; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7809 = unuse_way == 2'h2 ? valid_0_99 : _GEN_6395; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7810 = unuse_way == 2'h2 ? valid_0_100 : _GEN_6396; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7811 = unuse_way == 2'h2 ? valid_0_101 : _GEN_6397; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7812 = unuse_way == 2'h2 ? valid_0_102 : _GEN_6398; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7813 = unuse_way == 2'h2 ? valid_0_103 : _GEN_6399; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7814 = unuse_way == 2'h2 ? valid_0_104 : _GEN_6400; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7815 = unuse_way == 2'h2 ? valid_0_105 : _GEN_6401; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7816 = unuse_way == 2'h2 ? valid_0_106 : _GEN_6402; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7817 = unuse_way == 2'h2 ? valid_0_107 : _GEN_6403; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7818 = unuse_way == 2'h2 ? valid_0_108 : _GEN_6404; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7819 = unuse_way == 2'h2 ? valid_0_109 : _GEN_6405; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7820 = unuse_way == 2'h2 ? valid_0_110 : _GEN_6406; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7821 = unuse_way == 2'h2 ? valid_0_111 : _GEN_6407; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7822 = unuse_way == 2'h2 ? valid_0_112 : _GEN_6408; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7823 = unuse_way == 2'h2 ? valid_0_113 : _GEN_6409; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7824 = unuse_way == 2'h2 ? valid_0_114 : _GEN_6410; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7825 = unuse_way == 2'h2 ? valid_0_115 : _GEN_6411; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7826 = unuse_way == 2'h2 ? valid_0_116 : _GEN_6412; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7827 = unuse_way == 2'h2 ? valid_0_117 : _GEN_6413; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7828 = unuse_way == 2'h2 ? valid_0_118 : _GEN_6414; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7829 = unuse_way == 2'h2 ? valid_0_119 : _GEN_6415; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7830 = unuse_way == 2'h2 ? valid_0_120 : _GEN_6416; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7831 = unuse_way == 2'h2 ? valid_0_121 : _GEN_6417; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7832 = unuse_way == 2'h2 ? valid_0_122 : _GEN_6418; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7833 = unuse_way == 2'h2 ? valid_0_123 : _GEN_6419; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7834 = unuse_way == 2'h2 ? valid_0_124 : _GEN_6420; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7835 = unuse_way == 2'h2 ? valid_0_125 : _GEN_6421; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7836 = unuse_way == 2'h2 ? valid_0_126 : _GEN_6422; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7837 = unuse_way == 2'h2 ? valid_0_127 : _GEN_6423; // @[d_cache.scala 125:40 22:26]
  wire  _GEN_7838 = unuse_way == 2'h2 ? dirty_1_0 : _GEN_6682; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7839 = unuse_way == 2'h2 ? dirty_1_1 : _GEN_6683; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7840 = unuse_way == 2'h2 ? dirty_1_2 : _GEN_6684; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7841 = unuse_way == 2'h2 ? dirty_1_3 : _GEN_6685; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7842 = unuse_way == 2'h2 ? dirty_1_4 : _GEN_6686; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7843 = unuse_way == 2'h2 ? dirty_1_5 : _GEN_6687; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7844 = unuse_way == 2'h2 ? dirty_1_6 : _GEN_6688; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7845 = unuse_way == 2'h2 ? dirty_1_7 : _GEN_6689; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7846 = unuse_way == 2'h2 ? dirty_1_8 : _GEN_6690; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7847 = unuse_way == 2'h2 ? dirty_1_9 : _GEN_6691; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7848 = unuse_way == 2'h2 ? dirty_1_10 : _GEN_6692; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7849 = unuse_way == 2'h2 ? dirty_1_11 : _GEN_6693; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7850 = unuse_way == 2'h2 ? dirty_1_12 : _GEN_6694; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7851 = unuse_way == 2'h2 ? dirty_1_13 : _GEN_6695; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7852 = unuse_way == 2'h2 ? dirty_1_14 : _GEN_6696; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7853 = unuse_way == 2'h2 ? dirty_1_15 : _GEN_6697; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7854 = unuse_way == 2'h2 ? dirty_1_16 : _GEN_6698; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7855 = unuse_way == 2'h2 ? dirty_1_17 : _GEN_6699; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7856 = unuse_way == 2'h2 ? dirty_1_18 : _GEN_6700; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7857 = unuse_way == 2'h2 ? dirty_1_19 : _GEN_6701; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7858 = unuse_way == 2'h2 ? dirty_1_20 : _GEN_6702; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7859 = unuse_way == 2'h2 ? dirty_1_21 : _GEN_6703; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7860 = unuse_way == 2'h2 ? dirty_1_22 : _GEN_6704; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7861 = unuse_way == 2'h2 ? dirty_1_23 : _GEN_6705; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7862 = unuse_way == 2'h2 ? dirty_1_24 : _GEN_6706; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7863 = unuse_way == 2'h2 ? dirty_1_25 : _GEN_6707; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7864 = unuse_way == 2'h2 ? dirty_1_26 : _GEN_6708; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7865 = unuse_way == 2'h2 ? dirty_1_27 : _GEN_6709; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7866 = unuse_way == 2'h2 ? dirty_1_28 : _GEN_6710; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7867 = unuse_way == 2'h2 ? dirty_1_29 : _GEN_6711; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7868 = unuse_way == 2'h2 ? dirty_1_30 : _GEN_6712; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7869 = unuse_way == 2'h2 ? dirty_1_31 : _GEN_6713; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7870 = unuse_way == 2'h2 ? dirty_1_32 : _GEN_6714; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7871 = unuse_way == 2'h2 ? dirty_1_33 : _GEN_6715; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7872 = unuse_way == 2'h2 ? dirty_1_34 : _GEN_6716; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7873 = unuse_way == 2'h2 ? dirty_1_35 : _GEN_6717; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7874 = unuse_way == 2'h2 ? dirty_1_36 : _GEN_6718; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7875 = unuse_way == 2'h2 ? dirty_1_37 : _GEN_6719; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7876 = unuse_way == 2'h2 ? dirty_1_38 : _GEN_6720; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7877 = unuse_way == 2'h2 ? dirty_1_39 : _GEN_6721; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7878 = unuse_way == 2'h2 ? dirty_1_40 : _GEN_6722; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7879 = unuse_way == 2'h2 ? dirty_1_41 : _GEN_6723; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7880 = unuse_way == 2'h2 ? dirty_1_42 : _GEN_6724; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7881 = unuse_way == 2'h2 ? dirty_1_43 : _GEN_6725; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7882 = unuse_way == 2'h2 ? dirty_1_44 : _GEN_6726; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7883 = unuse_way == 2'h2 ? dirty_1_45 : _GEN_6727; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7884 = unuse_way == 2'h2 ? dirty_1_46 : _GEN_6728; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7885 = unuse_way == 2'h2 ? dirty_1_47 : _GEN_6729; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7886 = unuse_way == 2'h2 ? dirty_1_48 : _GEN_6730; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7887 = unuse_way == 2'h2 ? dirty_1_49 : _GEN_6731; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7888 = unuse_way == 2'h2 ? dirty_1_50 : _GEN_6732; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7889 = unuse_way == 2'h2 ? dirty_1_51 : _GEN_6733; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7890 = unuse_way == 2'h2 ? dirty_1_52 : _GEN_6734; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7891 = unuse_way == 2'h2 ? dirty_1_53 : _GEN_6735; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7892 = unuse_way == 2'h2 ? dirty_1_54 : _GEN_6736; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7893 = unuse_way == 2'h2 ? dirty_1_55 : _GEN_6737; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7894 = unuse_way == 2'h2 ? dirty_1_56 : _GEN_6738; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7895 = unuse_way == 2'h2 ? dirty_1_57 : _GEN_6739; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7896 = unuse_way == 2'h2 ? dirty_1_58 : _GEN_6740; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7897 = unuse_way == 2'h2 ? dirty_1_59 : _GEN_6741; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7898 = unuse_way == 2'h2 ? dirty_1_60 : _GEN_6742; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7899 = unuse_way == 2'h2 ? dirty_1_61 : _GEN_6743; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7900 = unuse_way == 2'h2 ? dirty_1_62 : _GEN_6744; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7901 = unuse_way == 2'h2 ? dirty_1_63 : _GEN_6745; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7902 = unuse_way == 2'h2 ? dirty_1_64 : _GEN_6746; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7903 = unuse_way == 2'h2 ? dirty_1_65 : _GEN_6747; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7904 = unuse_way == 2'h2 ? dirty_1_66 : _GEN_6748; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7905 = unuse_way == 2'h2 ? dirty_1_67 : _GEN_6749; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7906 = unuse_way == 2'h2 ? dirty_1_68 : _GEN_6750; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7907 = unuse_way == 2'h2 ? dirty_1_69 : _GEN_6751; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7908 = unuse_way == 2'h2 ? dirty_1_70 : _GEN_6752; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7909 = unuse_way == 2'h2 ? dirty_1_71 : _GEN_6753; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7910 = unuse_way == 2'h2 ? dirty_1_72 : _GEN_6754; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7911 = unuse_way == 2'h2 ? dirty_1_73 : _GEN_6755; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7912 = unuse_way == 2'h2 ? dirty_1_74 : _GEN_6756; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7913 = unuse_way == 2'h2 ? dirty_1_75 : _GEN_6757; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7914 = unuse_way == 2'h2 ? dirty_1_76 : _GEN_6758; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7915 = unuse_way == 2'h2 ? dirty_1_77 : _GEN_6759; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7916 = unuse_way == 2'h2 ? dirty_1_78 : _GEN_6760; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7917 = unuse_way == 2'h2 ? dirty_1_79 : _GEN_6761; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7918 = unuse_way == 2'h2 ? dirty_1_80 : _GEN_6762; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7919 = unuse_way == 2'h2 ? dirty_1_81 : _GEN_6763; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7920 = unuse_way == 2'h2 ? dirty_1_82 : _GEN_6764; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7921 = unuse_way == 2'h2 ? dirty_1_83 : _GEN_6765; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7922 = unuse_way == 2'h2 ? dirty_1_84 : _GEN_6766; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7923 = unuse_way == 2'h2 ? dirty_1_85 : _GEN_6767; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7924 = unuse_way == 2'h2 ? dirty_1_86 : _GEN_6768; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7925 = unuse_way == 2'h2 ? dirty_1_87 : _GEN_6769; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7926 = unuse_way == 2'h2 ? dirty_1_88 : _GEN_6770; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7927 = unuse_way == 2'h2 ? dirty_1_89 : _GEN_6771; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7928 = unuse_way == 2'h2 ? dirty_1_90 : _GEN_6772; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7929 = unuse_way == 2'h2 ? dirty_1_91 : _GEN_6773; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7930 = unuse_way == 2'h2 ? dirty_1_92 : _GEN_6774; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7931 = unuse_way == 2'h2 ? dirty_1_93 : _GEN_6775; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7932 = unuse_way == 2'h2 ? dirty_1_94 : _GEN_6776; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7933 = unuse_way == 2'h2 ? dirty_1_95 : _GEN_6777; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7934 = unuse_way == 2'h2 ? dirty_1_96 : _GEN_6778; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7935 = unuse_way == 2'h2 ? dirty_1_97 : _GEN_6779; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7936 = unuse_way == 2'h2 ? dirty_1_98 : _GEN_6780; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7937 = unuse_way == 2'h2 ? dirty_1_99 : _GEN_6781; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7938 = unuse_way == 2'h2 ? dirty_1_100 : _GEN_6782; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7939 = unuse_way == 2'h2 ? dirty_1_101 : _GEN_6783; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7940 = unuse_way == 2'h2 ? dirty_1_102 : _GEN_6784; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7941 = unuse_way == 2'h2 ? dirty_1_103 : _GEN_6785; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7942 = unuse_way == 2'h2 ? dirty_1_104 : _GEN_6786; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7943 = unuse_way == 2'h2 ? dirty_1_105 : _GEN_6787; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7944 = unuse_way == 2'h2 ? dirty_1_106 : _GEN_6788; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7945 = unuse_way == 2'h2 ? dirty_1_107 : _GEN_6789; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7946 = unuse_way == 2'h2 ? dirty_1_108 : _GEN_6790; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7947 = unuse_way == 2'h2 ? dirty_1_109 : _GEN_6791; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7948 = unuse_way == 2'h2 ? dirty_1_110 : _GEN_6792; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7949 = unuse_way == 2'h2 ? dirty_1_111 : _GEN_6793; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7950 = unuse_way == 2'h2 ? dirty_1_112 : _GEN_6794; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7951 = unuse_way == 2'h2 ? dirty_1_113 : _GEN_6795; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7952 = unuse_way == 2'h2 ? dirty_1_114 : _GEN_6796; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7953 = unuse_way == 2'h2 ? dirty_1_115 : _GEN_6797; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7954 = unuse_way == 2'h2 ? dirty_1_116 : _GEN_6798; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7955 = unuse_way == 2'h2 ? dirty_1_117 : _GEN_6799; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7956 = unuse_way == 2'h2 ? dirty_1_118 : _GEN_6800; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7957 = unuse_way == 2'h2 ? dirty_1_119 : _GEN_6801; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7958 = unuse_way == 2'h2 ? dirty_1_120 : _GEN_6802; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7959 = unuse_way == 2'h2 ? dirty_1_121 : _GEN_6803; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7960 = unuse_way == 2'h2 ? dirty_1_122 : _GEN_6804; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7961 = unuse_way == 2'h2 ? dirty_1_123 : _GEN_6805; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7962 = unuse_way == 2'h2 ? dirty_1_124 : _GEN_6806; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7963 = unuse_way == 2'h2 ? dirty_1_125 : _GEN_6807; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7964 = unuse_way == 2'h2 ? dirty_1_126 : _GEN_6808; // @[d_cache.scala 125:40 25:26]
  wire  _GEN_7965 = unuse_way == 2'h2 ? dirty_1_127 : _GEN_6809; // @[d_cache.scala 125:40 25:26]
  wire [2:0] _GEN_7966 = unuse_way == 2'h1 ? 3'h7 : _GEN_6938; // @[d_cache.scala 119:34 120:23]
  wire [63:0] _GEN_7967 = unuse_way == 2'h1 ? _GEN_2062 : _GEN_7326; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7968 = unuse_way == 2'h1 ? _GEN_2063 : _GEN_7327; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7969 = unuse_way == 2'h1 ? _GEN_2064 : _GEN_7328; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7970 = unuse_way == 2'h1 ? _GEN_2065 : _GEN_7329; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7971 = unuse_way == 2'h1 ? _GEN_2066 : _GEN_7330; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7972 = unuse_way == 2'h1 ? _GEN_2067 : _GEN_7331; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7973 = unuse_way == 2'h1 ? _GEN_2068 : _GEN_7332; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7974 = unuse_way == 2'h1 ? _GEN_2069 : _GEN_7333; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7975 = unuse_way == 2'h1 ? _GEN_2070 : _GEN_7334; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7976 = unuse_way == 2'h1 ? _GEN_2071 : _GEN_7335; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7977 = unuse_way == 2'h1 ? _GEN_2072 : _GEN_7336; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7978 = unuse_way == 2'h1 ? _GEN_2073 : _GEN_7337; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7979 = unuse_way == 2'h1 ? _GEN_2074 : _GEN_7338; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7980 = unuse_way == 2'h1 ? _GEN_2075 : _GEN_7339; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7981 = unuse_way == 2'h1 ? _GEN_2076 : _GEN_7340; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7982 = unuse_way == 2'h1 ? _GEN_2077 : _GEN_7341; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7983 = unuse_way == 2'h1 ? _GEN_2078 : _GEN_7342; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7984 = unuse_way == 2'h1 ? _GEN_2079 : _GEN_7343; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7985 = unuse_way == 2'h1 ? _GEN_2080 : _GEN_7344; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7986 = unuse_way == 2'h1 ? _GEN_2081 : _GEN_7345; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7987 = unuse_way == 2'h1 ? _GEN_2082 : _GEN_7346; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7988 = unuse_way == 2'h1 ? _GEN_2083 : _GEN_7347; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7989 = unuse_way == 2'h1 ? _GEN_2084 : _GEN_7348; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7990 = unuse_way == 2'h1 ? _GEN_2085 : _GEN_7349; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7991 = unuse_way == 2'h1 ? _GEN_2086 : _GEN_7350; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7992 = unuse_way == 2'h1 ? _GEN_2087 : _GEN_7351; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7993 = unuse_way == 2'h1 ? _GEN_2088 : _GEN_7352; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7994 = unuse_way == 2'h1 ? _GEN_2089 : _GEN_7353; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7995 = unuse_way == 2'h1 ? _GEN_2090 : _GEN_7354; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7996 = unuse_way == 2'h1 ? _GEN_2091 : _GEN_7355; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7997 = unuse_way == 2'h1 ? _GEN_2092 : _GEN_7356; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7998 = unuse_way == 2'h1 ? _GEN_2093 : _GEN_7357; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_7999 = unuse_way == 2'h1 ? _GEN_2094 : _GEN_7358; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8000 = unuse_way == 2'h1 ? _GEN_2095 : _GEN_7359; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8001 = unuse_way == 2'h1 ? _GEN_2096 : _GEN_7360; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8002 = unuse_way == 2'h1 ? _GEN_2097 : _GEN_7361; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8003 = unuse_way == 2'h1 ? _GEN_2098 : _GEN_7362; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8004 = unuse_way == 2'h1 ? _GEN_2099 : _GEN_7363; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8005 = unuse_way == 2'h1 ? _GEN_2100 : _GEN_7364; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8006 = unuse_way == 2'h1 ? _GEN_2101 : _GEN_7365; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8007 = unuse_way == 2'h1 ? _GEN_2102 : _GEN_7366; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8008 = unuse_way == 2'h1 ? _GEN_2103 : _GEN_7367; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8009 = unuse_way == 2'h1 ? _GEN_2104 : _GEN_7368; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8010 = unuse_way == 2'h1 ? _GEN_2105 : _GEN_7369; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8011 = unuse_way == 2'h1 ? _GEN_2106 : _GEN_7370; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8012 = unuse_way == 2'h1 ? _GEN_2107 : _GEN_7371; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8013 = unuse_way == 2'h1 ? _GEN_2108 : _GEN_7372; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8014 = unuse_way == 2'h1 ? _GEN_2109 : _GEN_7373; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8015 = unuse_way == 2'h1 ? _GEN_2110 : _GEN_7374; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8016 = unuse_way == 2'h1 ? _GEN_2111 : _GEN_7375; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8017 = unuse_way == 2'h1 ? _GEN_2112 : _GEN_7376; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8018 = unuse_way == 2'h1 ? _GEN_2113 : _GEN_7377; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8019 = unuse_way == 2'h1 ? _GEN_2114 : _GEN_7378; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8020 = unuse_way == 2'h1 ? _GEN_2115 : _GEN_7379; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8021 = unuse_way == 2'h1 ? _GEN_2116 : _GEN_7380; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8022 = unuse_way == 2'h1 ? _GEN_2117 : _GEN_7381; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8023 = unuse_way == 2'h1 ? _GEN_2118 : _GEN_7382; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8024 = unuse_way == 2'h1 ? _GEN_2119 : _GEN_7383; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8025 = unuse_way == 2'h1 ? _GEN_2120 : _GEN_7384; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8026 = unuse_way == 2'h1 ? _GEN_2121 : _GEN_7385; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8027 = unuse_way == 2'h1 ? _GEN_2122 : _GEN_7386; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8028 = unuse_way == 2'h1 ? _GEN_2123 : _GEN_7387; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8029 = unuse_way == 2'h1 ? _GEN_2124 : _GEN_7388; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8030 = unuse_way == 2'h1 ? _GEN_2125 : _GEN_7389; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8031 = unuse_way == 2'h1 ? _GEN_2126 : _GEN_7390; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8032 = unuse_way == 2'h1 ? _GEN_2127 : _GEN_7391; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8033 = unuse_way == 2'h1 ? _GEN_2128 : _GEN_7392; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8034 = unuse_way == 2'h1 ? _GEN_2129 : _GEN_7393; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8035 = unuse_way == 2'h1 ? _GEN_2130 : _GEN_7394; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8036 = unuse_way == 2'h1 ? _GEN_2131 : _GEN_7395; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8037 = unuse_way == 2'h1 ? _GEN_2132 : _GEN_7396; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8038 = unuse_way == 2'h1 ? _GEN_2133 : _GEN_7397; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8039 = unuse_way == 2'h1 ? _GEN_2134 : _GEN_7398; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8040 = unuse_way == 2'h1 ? _GEN_2135 : _GEN_7399; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8041 = unuse_way == 2'h1 ? _GEN_2136 : _GEN_7400; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8042 = unuse_way == 2'h1 ? _GEN_2137 : _GEN_7401; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8043 = unuse_way == 2'h1 ? _GEN_2138 : _GEN_7402; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8044 = unuse_way == 2'h1 ? _GEN_2139 : _GEN_7403; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8045 = unuse_way == 2'h1 ? _GEN_2140 : _GEN_7404; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8046 = unuse_way == 2'h1 ? _GEN_2141 : _GEN_7405; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8047 = unuse_way == 2'h1 ? _GEN_2142 : _GEN_7406; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8048 = unuse_way == 2'h1 ? _GEN_2143 : _GEN_7407; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8049 = unuse_way == 2'h1 ? _GEN_2144 : _GEN_7408; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8050 = unuse_way == 2'h1 ? _GEN_2145 : _GEN_7409; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8051 = unuse_way == 2'h1 ? _GEN_2146 : _GEN_7410; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8052 = unuse_way == 2'h1 ? _GEN_2147 : _GEN_7411; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8053 = unuse_way == 2'h1 ? _GEN_2148 : _GEN_7412; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8054 = unuse_way == 2'h1 ? _GEN_2149 : _GEN_7413; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8055 = unuse_way == 2'h1 ? _GEN_2150 : _GEN_7414; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8056 = unuse_way == 2'h1 ? _GEN_2151 : _GEN_7415; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8057 = unuse_way == 2'h1 ? _GEN_2152 : _GEN_7416; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8058 = unuse_way == 2'h1 ? _GEN_2153 : _GEN_7417; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8059 = unuse_way == 2'h1 ? _GEN_2154 : _GEN_7418; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8060 = unuse_way == 2'h1 ? _GEN_2155 : _GEN_7419; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8061 = unuse_way == 2'h1 ? _GEN_2156 : _GEN_7420; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8062 = unuse_way == 2'h1 ? _GEN_2157 : _GEN_7421; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8063 = unuse_way == 2'h1 ? _GEN_2158 : _GEN_7422; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8064 = unuse_way == 2'h1 ? _GEN_2159 : _GEN_7423; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8065 = unuse_way == 2'h1 ? _GEN_2160 : _GEN_7424; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8066 = unuse_way == 2'h1 ? _GEN_2161 : _GEN_7425; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8067 = unuse_way == 2'h1 ? _GEN_2162 : _GEN_7426; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8068 = unuse_way == 2'h1 ? _GEN_2163 : _GEN_7427; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8069 = unuse_way == 2'h1 ? _GEN_2164 : _GEN_7428; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8070 = unuse_way == 2'h1 ? _GEN_2165 : _GEN_7429; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8071 = unuse_way == 2'h1 ? _GEN_2166 : _GEN_7430; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8072 = unuse_way == 2'h1 ? _GEN_2167 : _GEN_7431; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8073 = unuse_way == 2'h1 ? _GEN_2168 : _GEN_7432; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8074 = unuse_way == 2'h1 ? _GEN_2169 : _GEN_7433; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8075 = unuse_way == 2'h1 ? _GEN_2170 : _GEN_7434; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8076 = unuse_way == 2'h1 ? _GEN_2171 : _GEN_7435; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8077 = unuse_way == 2'h1 ? _GEN_2172 : _GEN_7436; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8078 = unuse_way == 2'h1 ? _GEN_2173 : _GEN_7437; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8079 = unuse_way == 2'h1 ? _GEN_2174 : _GEN_7438; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8080 = unuse_way == 2'h1 ? _GEN_2175 : _GEN_7439; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8081 = unuse_way == 2'h1 ? _GEN_2176 : _GEN_7440; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8082 = unuse_way == 2'h1 ? _GEN_2177 : _GEN_7441; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8083 = unuse_way == 2'h1 ? _GEN_2178 : _GEN_7442; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8084 = unuse_way == 2'h1 ? _GEN_2179 : _GEN_7443; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8085 = unuse_way == 2'h1 ? _GEN_2180 : _GEN_7444; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8086 = unuse_way == 2'h1 ? _GEN_2181 : _GEN_7445; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8087 = unuse_way == 2'h1 ? _GEN_2182 : _GEN_7446; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8088 = unuse_way == 2'h1 ? _GEN_2183 : _GEN_7447; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8089 = unuse_way == 2'h1 ? _GEN_2184 : _GEN_7448; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8090 = unuse_way == 2'h1 ? _GEN_2185 : _GEN_7449; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8091 = unuse_way == 2'h1 ? _GEN_2186 : _GEN_7450; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8092 = unuse_way == 2'h1 ? _GEN_2187 : _GEN_7451; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8093 = unuse_way == 2'h1 ? _GEN_2188 : _GEN_7452; // @[d_cache.scala 119:34]
  wire [63:0] _GEN_8094 = unuse_way == 2'h1 ? _GEN_2189 : _GEN_7453; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8095 = unuse_way == 2'h1 ? _GEN_2190 : _GEN_7454; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8096 = unuse_way == 2'h1 ? _GEN_2191 : _GEN_7455; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8097 = unuse_way == 2'h1 ? _GEN_2192 : _GEN_7456; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8098 = unuse_way == 2'h1 ? _GEN_2193 : _GEN_7457; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8099 = unuse_way == 2'h1 ? _GEN_2194 : _GEN_7458; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8100 = unuse_way == 2'h1 ? _GEN_2195 : _GEN_7459; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8101 = unuse_way == 2'h1 ? _GEN_2196 : _GEN_7460; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8102 = unuse_way == 2'h1 ? _GEN_2197 : _GEN_7461; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8103 = unuse_way == 2'h1 ? _GEN_2198 : _GEN_7462; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8104 = unuse_way == 2'h1 ? _GEN_2199 : _GEN_7463; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8105 = unuse_way == 2'h1 ? _GEN_2200 : _GEN_7464; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8106 = unuse_way == 2'h1 ? _GEN_2201 : _GEN_7465; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8107 = unuse_way == 2'h1 ? _GEN_2202 : _GEN_7466; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8108 = unuse_way == 2'h1 ? _GEN_2203 : _GEN_7467; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8109 = unuse_way == 2'h1 ? _GEN_2204 : _GEN_7468; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8110 = unuse_way == 2'h1 ? _GEN_2205 : _GEN_7469; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8111 = unuse_way == 2'h1 ? _GEN_2206 : _GEN_7470; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8112 = unuse_way == 2'h1 ? _GEN_2207 : _GEN_7471; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8113 = unuse_way == 2'h1 ? _GEN_2208 : _GEN_7472; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8114 = unuse_way == 2'h1 ? _GEN_2209 : _GEN_7473; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8115 = unuse_way == 2'h1 ? _GEN_2210 : _GEN_7474; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8116 = unuse_way == 2'h1 ? _GEN_2211 : _GEN_7475; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8117 = unuse_way == 2'h1 ? _GEN_2212 : _GEN_7476; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8118 = unuse_way == 2'h1 ? _GEN_2213 : _GEN_7477; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8119 = unuse_way == 2'h1 ? _GEN_2214 : _GEN_7478; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8120 = unuse_way == 2'h1 ? _GEN_2215 : _GEN_7479; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8121 = unuse_way == 2'h1 ? _GEN_2216 : _GEN_7480; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8122 = unuse_way == 2'h1 ? _GEN_2217 : _GEN_7481; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8123 = unuse_way == 2'h1 ? _GEN_2218 : _GEN_7482; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8124 = unuse_way == 2'h1 ? _GEN_2219 : _GEN_7483; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8125 = unuse_way == 2'h1 ? _GEN_2220 : _GEN_7484; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8126 = unuse_way == 2'h1 ? _GEN_2221 : _GEN_7485; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8127 = unuse_way == 2'h1 ? _GEN_2222 : _GEN_7486; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8128 = unuse_way == 2'h1 ? _GEN_2223 : _GEN_7487; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8129 = unuse_way == 2'h1 ? _GEN_2224 : _GEN_7488; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8130 = unuse_way == 2'h1 ? _GEN_2225 : _GEN_7489; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8131 = unuse_way == 2'h1 ? _GEN_2226 : _GEN_7490; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8132 = unuse_way == 2'h1 ? _GEN_2227 : _GEN_7491; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8133 = unuse_way == 2'h1 ? _GEN_2228 : _GEN_7492; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8134 = unuse_way == 2'h1 ? _GEN_2229 : _GEN_7493; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8135 = unuse_way == 2'h1 ? _GEN_2230 : _GEN_7494; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8136 = unuse_way == 2'h1 ? _GEN_2231 : _GEN_7495; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8137 = unuse_way == 2'h1 ? _GEN_2232 : _GEN_7496; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8138 = unuse_way == 2'h1 ? _GEN_2233 : _GEN_7497; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8139 = unuse_way == 2'h1 ? _GEN_2234 : _GEN_7498; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8140 = unuse_way == 2'h1 ? _GEN_2235 : _GEN_7499; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8141 = unuse_way == 2'h1 ? _GEN_2236 : _GEN_7500; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8142 = unuse_way == 2'h1 ? _GEN_2237 : _GEN_7501; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8143 = unuse_way == 2'h1 ? _GEN_2238 : _GEN_7502; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8144 = unuse_way == 2'h1 ? _GEN_2239 : _GEN_7503; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8145 = unuse_way == 2'h1 ? _GEN_2240 : _GEN_7504; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8146 = unuse_way == 2'h1 ? _GEN_2241 : _GEN_7505; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8147 = unuse_way == 2'h1 ? _GEN_2242 : _GEN_7506; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8148 = unuse_way == 2'h1 ? _GEN_2243 : _GEN_7507; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8149 = unuse_way == 2'h1 ? _GEN_2244 : _GEN_7508; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8150 = unuse_way == 2'h1 ? _GEN_2245 : _GEN_7509; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8151 = unuse_way == 2'h1 ? _GEN_2246 : _GEN_7510; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8152 = unuse_way == 2'h1 ? _GEN_2247 : _GEN_7511; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8153 = unuse_way == 2'h1 ? _GEN_2248 : _GEN_7512; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8154 = unuse_way == 2'h1 ? _GEN_2249 : _GEN_7513; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8155 = unuse_way == 2'h1 ? _GEN_2250 : _GEN_7514; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8156 = unuse_way == 2'h1 ? _GEN_2251 : _GEN_7515; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8157 = unuse_way == 2'h1 ? _GEN_2252 : _GEN_7516; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8158 = unuse_way == 2'h1 ? _GEN_2253 : _GEN_7517; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8159 = unuse_way == 2'h1 ? _GEN_2254 : _GEN_7518; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8160 = unuse_way == 2'h1 ? _GEN_2255 : _GEN_7519; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8161 = unuse_way == 2'h1 ? _GEN_2256 : _GEN_7520; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8162 = unuse_way == 2'h1 ? _GEN_2257 : _GEN_7521; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8163 = unuse_way == 2'h1 ? _GEN_2258 : _GEN_7522; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8164 = unuse_way == 2'h1 ? _GEN_2259 : _GEN_7523; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8165 = unuse_way == 2'h1 ? _GEN_2260 : _GEN_7524; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8166 = unuse_way == 2'h1 ? _GEN_2261 : _GEN_7525; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8167 = unuse_way == 2'h1 ? _GEN_2262 : _GEN_7526; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8168 = unuse_way == 2'h1 ? _GEN_2263 : _GEN_7527; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8169 = unuse_way == 2'h1 ? _GEN_2264 : _GEN_7528; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8170 = unuse_way == 2'h1 ? _GEN_2265 : _GEN_7529; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8171 = unuse_way == 2'h1 ? _GEN_2266 : _GEN_7530; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8172 = unuse_way == 2'h1 ? _GEN_2267 : _GEN_7531; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8173 = unuse_way == 2'h1 ? _GEN_2268 : _GEN_7532; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8174 = unuse_way == 2'h1 ? _GEN_2269 : _GEN_7533; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8175 = unuse_way == 2'h1 ? _GEN_2270 : _GEN_7534; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8176 = unuse_way == 2'h1 ? _GEN_2271 : _GEN_7535; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8177 = unuse_way == 2'h1 ? _GEN_2272 : _GEN_7536; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8178 = unuse_way == 2'h1 ? _GEN_2273 : _GEN_7537; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8179 = unuse_way == 2'h1 ? _GEN_2274 : _GEN_7538; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8180 = unuse_way == 2'h1 ? _GEN_2275 : _GEN_7539; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8181 = unuse_way == 2'h1 ? _GEN_2276 : _GEN_7540; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8182 = unuse_way == 2'h1 ? _GEN_2277 : _GEN_7541; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8183 = unuse_way == 2'h1 ? _GEN_2278 : _GEN_7542; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8184 = unuse_way == 2'h1 ? _GEN_2279 : _GEN_7543; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8185 = unuse_way == 2'h1 ? _GEN_2280 : _GEN_7544; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8186 = unuse_way == 2'h1 ? _GEN_2281 : _GEN_7545; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8187 = unuse_way == 2'h1 ? _GEN_2282 : _GEN_7546; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8188 = unuse_way == 2'h1 ? _GEN_2283 : _GEN_7547; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8189 = unuse_way == 2'h1 ? _GEN_2284 : _GEN_7548; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8190 = unuse_way == 2'h1 ? _GEN_2285 : _GEN_7549; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8191 = unuse_way == 2'h1 ? _GEN_2286 : _GEN_7550; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8192 = unuse_way == 2'h1 ? _GEN_2287 : _GEN_7551; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8193 = unuse_way == 2'h1 ? _GEN_2288 : _GEN_7552; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8194 = unuse_way == 2'h1 ? _GEN_2289 : _GEN_7553; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8195 = unuse_way == 2'h1 ? _GEN_2290 : _GEN_7554; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8196 = unuse_way == 2'h1 ? _GEN_2291 : _GEN_7555; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8197 = unuse_way == 2'h1 ? _GEN_2292 : _GEN_7556; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8198 = unuse_way == 2'h1 ? _GEN_2293 : _GEN_7557; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8199 = unuse_way == 2'h1 ? _GEN_2294 : _GEN_7558; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8200 = unuse_way == 2'h1 ? _GEN_2295 : _GEN_7559; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8201 = unuse_way == 2'h1 ? _GEN_2296 : _GEN_7560; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8202 = unuse_way == 2'h1 ? _GEN_2297 : _GEN_7561; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8203 = unuse_way == 2'h1 ? _GEN_2298 : _GEN_7562; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8204 = unuse_way == 2'h1 ? _GEN_2299 : _GEN_7563; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8205 = unuse_way == 2'h1 ? _GEN_2300 : _GEN_7564; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8206 = unuse_way == 2'h1 ? _GEN_2301 : _GEN_7565; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8207 = unuse_way == 2'h1 ? _GEN_2302 : _GEN_7566; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8208 = unuse_way == 2'h1 ? _GEN_2303 : _GEN_7567; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8209 = unuse_way == 2'h1 ? _GEN_2304 : _GEN_7568; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8210 = unuse_way == 2'h1 ? _GEN_2305 : _GEN_7569; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8211 = unuse_way == 2'h1 ? _GEN_2306 : _GEN_7570; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8212 = unuse_way == 2'h1 ? _GEN_2307 : _GEN_7571; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8213 = unuse_way == 2'h1 ? _GEN_2308 : _GEN_7572; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8214 = unuse_way == 2'h1 ? _GEN_2309 : _GEN_7573; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8215 = unuse_way == 2'h1 ? _GEN_2310 : _GEN_7574; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8216 = unuse_way == 2'h1 ? _GEN_2311 : _GEN_7575; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8217 = unuse_way == 2'h1 ? _GEN_2312 : _GEN_7576; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8218 = unuse_way == 2'h1 ? _GEN_2313 : _GEN_7577; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8219 = unuse_way == 2'h1 ? _GEN_2314 : _GEN_7578; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8220 = unuse_way == 2'h1 ? _GEN_2315 : _GEN_7579; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8221 = unuse_way == 2'h1 ? _GEN_2316 : _GEN_7580; // @[d_cache.scala 119:34]
  wire [31:0] _GEN_8222 = unuse_way == 2'h1 ? _GEN_2317 : _GEN_7581; // @[d_cache.scala 119:34]
  wire  _GEN_8223 = unuse_way == 2'h1 ? _GEN_2318 : _GEN_7710; // @[d_cache.scala 119:34]
  wire  _GEN_8224 = unuse_way == 2'h1 ? _GEN_2319 : _GEN_7711; // @[d_cache.scala 119:34]
  wire  _GEN_8225 = unuse_way == 2'h1 ? _GEN_2320 : _GEN_7712; // @[d_cache.scala 119:34]
  wire  _GEN_8226 = unuse_way == 2'h1 ? _GEN_2321 : _GEN_7713; // @[d_cache.scala 119:34]
  wire  _GEN_8227 = unuse_way == 2'h1 ? _GEN_2322 : _GEN_7714; // @[d_cache.scala 119:34]
  wire  _GEN_8228 = unuse_way == 2'h1 ? _GEN_2323 : _GEN_7715; // @[d_cache.scala 119:34]
  wire  _GEN_8229 = unuse_way == 2'h1 ? _GEN_2324 : _GEN_7716; // @[d_cache.scala 119:34]
  wire  _GEN_8230 = unuse_way == 2'h1 ? _GEN_2325 : _GEN_7717; // @[d_cache.scala 119:34]
  wire  _GEN_8231 = unuse_way == 2'h1 ? _GEN_2326 : _GEN_7718; // @[d_cache.scala 119:34]
  wire  _GEN_8232 = unuse_way == 2'h1 ? _GEN_2327 : _GEN_7719; // @[d_cache.scala 119:34]
  wire  _GEN_8233 = unuse_way == 2'h1 ? _GEN_2328 : _GEN_7720; // @[d_cache.scala 119:34]
  wire  _GEN_8234 = unuse_way == 2'h1 ? _GEN_2329 : _GEN_7721; // @[d_cache.scala 119:34]
  wire  _GEN_8235 = unuse_way == 2'h1 ? _GEN_2330 : _GEN_7722; // @[d_cache.scala 119:34]
  wire  _GEN_8236 = unuse_way == 2'h1 ? _GEN_2331 : _GEN_7723; // @[d_cache.scala 119:34]
  wire  _GEN_8237 = unuse_way == 2'h1 ? _GEN_2332 : _GEN_7724; // @[d_cache.scala 119:34]
  wire  _GEN_8238 = unuse_way == 2'h1 ? _GEN_2333 : _GEN_7725; // @[d_cache.scala 119:34]
  wire  _GEN_8239 = unuse_way == 2'h1 ? _GEN_2334 : _GEN_7726; // @[d_cache.scala 119:34]
  wire  _GEN_8240 = unuse_way == 2'h1 ? _GEN_2335 : _GEN_7727; // @[d_cache.scala 119:34]
  wire  _GEN_8241 = unuse_way == 2'h1 ? _GEN_2336 : _GEN_7728; // @[d_cache.scala 119:34]
  wire  _GEN_8242 = unuse_way == 2'h1 ? _GEN_2337 : _GEN_7729; // @[d_cache.scala 119:34]
  wire  _GEN_8243 = unuse_way == 2'h1 ? _GEN_2338 : _GEN_7730; // @[d_cache.scala 119:34]
  wire  _GEN_8244 = unuse_way == 2'h1 ? _GEN_2339 : _GEN_7731; // @[d_cache.scala 119:34]
  wire  _GEN_8245 = unuse_way == 2'h1 ? _GEN_2340 : _GEN_7732; // @[d_cache.scala 119:34]
  wire  _GEN_8246 = unuse_way == 2'h1 ? _GEN_2341 : _GEN_7733; // @[d_cache.scala 119:34]
  wire  _GEN_8247 = unuse_way == 2'h1 ? _GEN_2342 : _GEN_7734; // @[d_cache.scala 119:34]
  wire  _GEN_8248 = unuse_way == 2'h1 ? _GEN_2343 : _GEN_7735; // @[d_cache.scala 119:34]
  wire  _GEN_8249 = unuse_way == 2'h1 ? _GEN_2344 : _GEN_7736; // @[d_cache.scala 119:34]
  wire  _GEN_8250 = unuse_way == 2'h1 ? _GEN_2345 : _GEN_7737; // @[d_cache.scala 119:34]
  wire  _GEN_8251 = unuse_way == 2'h1 ? _GEN_2346 : _GEN_7738; // @[d_cache.scala 119:34]
  wire  _GEN_8252 = unuse_way == 2'h1 ? _GEN_2347 : _GEN_7739; // @[d_cache.scala 119:34]
  wire  _GEN_8253 = unuse_way == 2'h1 ? _GEN_2348 : _GEN_7740; // @[d_cache.scala 119:34]
  wire  _GEN_8254 = unuse_way == 2'h1 ? _GEN_2349 : _GEN_7741; // @[d_cache.scala 119:34]
  wire  _GEN_8255 = unuse_way == 2'h1 ? _GEN_2350 : _GEN_7742; // @[d_cache.scala 119:34]
  wire  _GEN_8256 = unuse_way == 2'h1 ? _GEN_2351 : _GEN_7743; // @[d_cache.scala 119:34]
  wire  _GEN_8257 = unuse_way == 2'h1 ? _GEN_2352 : _GEN_7744; // @[d_cache.scala 119:34]
  wire  _GEN_8258 = unuse_way == 2'h1 ? _GEN_2353 : _GEN_7745; // @[d_cache.scala 119:34]
  wire  _GEN_8259 = unuse_way == 2'h1 ? _GEN_2354 : _GEN_7746; // @[d_cache.scala 119:34]
  wire  _GEN_8260 = unuse_way == 2'h1 ? _GEN_2355 : _GEN_7747; // @[d_cache.scala 119:34]
  wire  _GEN_8261 = unuse_way == 2'h1 ? _GEN_2356 : _GEN_7748; // @[d_cache.scala 119:34]
  wire  _GEN_8262 = unuse_way == 2'h1 ? _GEN_2357 : _GEN_7749; // @[d_cache.scala 119:34]
  wire  _GEN_8263 = unuse_way == 2'h1 ? _GEN_2358 : _GEN_7750; // @[d_cache.scala 119:34]
  wire  _GEN_8264 = unuse_way == 2'h1 ? _GEN_2359 : _GEN_7751; // @[d_cache.scala 119:34]
  wire  _GEN_8265 = unuse_way == 2'h1 ? _GEN_2360 : _GEN_7752; // @[d_cache.scala 119:34]
  wire  _GEN_8266 = unuse_way == 2'h1 ? _GEN_2361 : _GEN_7753; // @[d_cache.scala 119:34]
  wire  _GEN_8267 = unuse_way == 2'h1 ? _GEN_2362 : _GEN_7754; // @[d_cache.scala 119:34]
  wire  _GEN_8268 = unuse_way == 2'h1 ? _GEN_2363 : _GEN_7755; // @[d_cache.scala 119:34]
  wire  _GEN_8269 = unuse_way == 2'h1 ? _GEN_2364 : _GEN_7756; // @[d_cache.scala 119:34]
  wire  _GEN_8270 = unuse_way == 2'h1 ? _GEN_2365 : _GEN_7757; // @[d_cache.scala 119:34]
  wire  _GEN_8271 = unuse_way == 2'h1 ? _GEN_2366 : _GEN_7758; // @[d_cache.scala 119:34]
  wire  _GEN_8272 = unuse_way == 2'h1 ? _GEN_2367 : _GEN_7759; // @[d_cache.scala 119:34]
  wire  _GEN_8273 = unuse_way == 2'h1 ? _GEN_2368 : _GEN_7760; // @[d_cache.scala 119:34]
  wire  _GEN_8274 = unuse_way == 2'h1 ? _GEN_2369 : _GEN_7761; // @[d_cache.scala 119:34]
  wire  _GEN_8275 = unuse_way == 2'h1 ? _GEN_2370 : _GEN_7762; // @[d_cache.scala 119:34]
  wire  _GEN_8276 = unuse_way == 2'h1 ? _GEN_2371 : _GEN_7763; // @[d_cache.scala 119:34]
  wire  _GEN_8277 = unuse_way == 2'h1 ? _GEN_2372 : _GEN_7764; // @[d_cache.scala 119:34]
  wire  _GEN_8278 = unuse_way == 2'h1 ? _GEN_2373 : _GEN_7765; // @[d_cache.scala 119:34]
  wire  _GEN_8279 = unuse_way == 2'h1 ? _GEN_2374 : _GEN_7766; // @[d_cache.scala 119:34]
  wire  _GEN_8280 = unuse_way == 2'h1 ? _GEN_2375 : _GEN_7767; // @[d_cache.scala 119:34]
  wire  _GEN_8281 = unuse_way == 2'h1 ? _GEN_2376 : _GEN_7768; // @[d_cache.scala 119:34]
  wire  _GEN_8282 = unuse_way == 2'h1 ? _GEN_2377 : _GEN_7769; // @[d_cache.scala 119:34]
  wire  _GEN_8283 = unuse_way == 2'h1 ? _GEN_2378 : _GEN_7770; // @[d_cache.scala 119:34]
  wire  _GEN_8284 = unuse_way == 2'h1 ? _GEN_2379 : _GEN_7771; // @[d_cache.scala 119:34]
  wire  _GEN_8285 = unuse_way == 2'h1 ? _GEN_2380 : _GEN_7772; // @[d_cache.scala 119:34]
  wire  _GEN_8286 = unuse_way == 2'h1 ? _GEN_2381 : _GEN_7773; // @[d_cache.scala 119:34]
  wire  _GEN_8287 = unuse_way == 2'h1 ? _GEN_2382 : _GEN_7774; // @[d_cache.scala 119:34]
  wire  _GEN_8288 = unuse_way == 2'h1 ? _GEN_2383 : _GEN_7775; // @[d_cache.scala 119:34]
  wire  _GEN_8289 = unuse_way == 2'h1 ? _GEN_2384 : _GEN_7776; // @[d_cache.scala 119:34]
  wire  _GEN_8290 = unuse_way == 2'h1 ? _GEN_2385 : _GEN_7777; // @[d_cache.scala 119:34]
  wire  _GEN_8291 = unuse_way == 2'h1 ? _GEN_2386 : _GEN_7778; // @[d_cache.scala 119:34]
  wire  _GEN_8292 = unuse_way == 2'h1 ? _GEN_2387 : _GEN_7779; // @[d_cache.scala 119:34]
  wire  _GEN_8293 = unuse_way == 2'h1 ? _GEN_2388 : _GEN_7780; // @[d_cache.scala 119:34]
  wire  _GEN_8294 = unuse_way == 2'h1 ? _GEN_2389 : _GEN_7781; // @[d_cache.scala 119:34]
  wire  _GEN_8295 = unuse_way == 2'h1 ? _GEN_2390 : _GEN_7782; // @[d_cache.scala 119:34]
  wire  _GEN_8296 = unuse_way == 2'h1 ? _GEN_2391 : _GEN_7783; // @[d_cache.scala 119:34]
  wire  _GEN_8297 = unuse_way == 2'h1 ? _GEN_2392 : _GEN_7784; // @[d_cache.scala 119:34]
  wire  _GEN_8298 = unuse_way == 2'h1 ? _GEN_2393 : _GEN_7785; // @[d_cache.scala 119:34]
  wire  _GEN_8299 = unuse_way == 2'h1 ? _GEN_2394 : _GEN_7786; // @[d_cache.scala 119:34]
  wire  _GEN_8300 = unuse_way == 2'h1 ? _GEN_2395 : _GEN_7787; // @[d_cache.scala 119:34]
  wire  _GEN_8301 = unuse_way == 2'h1 ? _GEN_2396 : _GEN_7788; // @[d_cache.scala 119:34]
  wire  _GEN_8302 = unuse_way == 2'h1 ? _GEN_2397 : _GEN_7789; // @[d_cache.scala 119:34]
  wire  _GEN_8303 = unuse_way == 2'h1 ? _GEN_2398 : _GEN_7790; // @[d_cache.scala 119:34]
  wire  _GEN_8304 = unuse_way == 2'h1 ? _GEN_2399 : _GEN_7791; // @[d_cache.scala 119:34]
  wire  _GEN_8305 = unuse_way == 2'h1 ? _GEN_2400 : _GEN_7792; // @[d_cache.scala 119:34]
  wire  _GEN_8306 = unuse_way == 2'h1 ? _GEN_2401 : _GEN_7793; // @[d_cache.scala 119:34]
  wire  _GEN_8307 = unuse_way == 2'h1 ? _GEN_2402 : _GEN_7794; // @[d_cache.scala 119:34]
  wire  _GEN_8308 = unuse_way == 2'h1 ? _GEN_2403 : _GEN_7795; // @[d_cache.scala 119:34]
  wire  _GEN_8309 = unuse_way == 2'h1 ? _GEN_2404 : _GEN_7796; // @[d_cache.scala 119:34]
  wire  _GEN_8310 = unuse_way == 2'h1 ? _GEN_2405 : _GEN_7797; // @[d_cache.scala 119:34]
  wire  _GEN_8311 = unuse_way == 2'h1 ? _GEN_2406 : _GEN_7798; // @[d_cache.scala 119:34]
  wire  _GEN_8312 = unuse_way == 2'h1 ? _GEN_2407 : _GEN_7799; // @[d_cache.scala 119:34]
  wire  _GEN_8313 = unuse_way == 2'h1 ? _GEN_2408 : _GEN_7800; // @[d_cache.scala 119:34]
  wire  _GEN_8314 = unuse_way == 2'h1 ? _GEN_2409 : _GEN_7801; // @[d_cache.scala 119:34]
  wire  _GEN_8315 = unuse_way == 2'h1 ? _GEN_2410 : _GEN_7802; // @[d_cache.scala 119:34]
  wire  _GEN_8316 = unuse_way == 2'h1 ? _GEN_2411 : _GEN_7803; // @[d_cache.scala 119:34]
  wire  _GEN_8317 = unuse_way == 2'h1 ? _GEN_2412 : _GEN_7804; // @[d_cache.scala 119:34]
  wire  _GEN_8318 = unuse_way == 2'h1 ? _GEN_2413 : _GEN_7805; // @[d_cache.scala 119:34]
  wire  _GEN_8319 = unuse_way == 2'h1 ? _GEN_2414 : _GEN_7806; // @[d_cache.scala 119:34]
  wire  _GEN_8320 = unuse_way == 2'h1 ? _GEN_2415 : _GEN_7807; // @[d_cache.scala 119:34]
  wire  _GEN_8321 = unuse_way == 2'h1 ? _GEN_2416 : _GEN_7808; // @[d_cache.scala 119:34]
  wire  _GEN_8322 = unuse_way == 2'h1 ? _GEN_2417 : _GEN_7809; // @[d_cache.scala 119:34]
  wire  _GEN_8323 = unuse_way == 2'h1 ? _GEN_2418 : _GEN_7810; // @[d_cache.scala 119:34]
  wire  _GEN_8324 = unuse_way == 2'h1 ? _GEN_2419 : _GEN_7811; // @[d_cache.scala 119:34]
  wire  _GEN_8325 = unuse_way == 2'h1 ? _GEN_2420 : _GEN_7812; // @[d_cache.scala 119:34]
  wire  _GEN_8326 = unuse_way == 2'h1 ? _GEN_2421 : _GEN_7813; // @[d_cache.scala 119:34]
  wire  _GEN_8327 = unuse_way == 2'h1 ? _GEN_2422 : _GEN_7814; // @[d_cache.scala 119:34]
  wire  _GEN_8328 = unuse_way == 2'h1 ? _GEN_2423 : _GEN_7815; // @[d_cache.scala 119:34]
  wire  _GEN_8329 = unuse_way == 2'h1 ? _GEN_2424 : _GEN_7816; // @[d_cache.scala 119:34]
  wire  _GEN_8330 = unuse_way == 2'h1 ? _GEN_2425 : _GEN_7817; // @[d_cache.scala 119:34]
  wire  _GEN_8331 = unuse_way == 2'h1 ? _GEN_2426 : _GEN_7818; // @[d_cache.scala 119:34]
  wire  _GEN_8332 = unuse_way == 2'h1 ? _GEN_2427 : _GEN_7819; // @[d_cache.scala 119:34]
  wire  _GEN_8333 = unuse_way == 2'h1 ? _GEN_2428 : _GEN_7820; // @[d_cache.scala 119:34]
  wire  _GEN_8334 = unuse_way == 2'h1 ? _GEN_2429 : _GEN_7821; // @[d_cache.scala 119:34]
  wire  _GEN_8335 = unuse_way == 2'h1 ? _GEN_2430 : _GEN_7822; // @[d_cache.scala 119:34]
  wire  _GEN_8336 = unuse_way == 2'h1 ? _GEN_2431 : _GEN_7823; // @[d_cache.scala 119:34]
  wire  _GEN_8337 = unuse_way == 2'h1 ? _GEN_2432 : _GEN_7824; // @[d_cache.scala 119:34]
  wire  _GEN_8338 = unuse_way == 2'h1 ? _GEN_2433 : _GEN_7825; // @[d_cache.scala 119:34]
  wire  _GEN_8339 = unuse_way == 2'h1 ? _GEN_2434 : _GEN_7826; // @[d_cache.scala 119:34]
  wire  _GEN_8340 = unuse_way == 2'h1 ? _GEN_2435 : _GEN_7827; // @[d_cache.scala 119:34]
  wire  _GEN_8341 = unuse_way == 2'h1 ? _GEN_2436 : _GEN_7828; // @[d_cache.scala 119:34]
  wire  _GEN_8342 = unuse_way == 2'h1 ? _GEN_2437 : _GEN_7829; // @[d_cache.scala 119:34]
  wire  _GEN_8343 = unuse_way == 2'h1 ? _GEN_2438 : _GEN_7830; // @[d_cache.scala 119:34]
  wire  _GEN_8344 = unuse_way == 2'h1 ? _GEN_2439 : _GEN_7831; // @[d_cache.scala 119:34]
  wire  _GEN_8345 = unuse_way == 2'h1 ? _GEN_2440 : _GEN_7832; // @[d_cache.scala 119:34]
  wire  _GEN_8346 = unuse_way == 2'h1 ? _GEN_2441 : _GEN_7833; // @[d_cache.scala 119:34]
  wire  _GEN_8347 = unuse_way == 2'h1 ? _GEN_2442 : _GEN_7834; // @[d_cache.scala 119:34]
  wire  _GEN_8348 = unuse_way == 2'h1 ? _GEN_2443 : _GEN_7835; // @[d_cache.scala 119:34]
  wire  _GEN_8349 = unuse_way == 2'h1 ? _GEN_2444 : _GEN_7836; // @[d_cache.scala 119:34]
  wire  _GEN_8350 = unuse_way == 2'h1 ? _GEN_2445 : _GEN_7837; // @[d_cache.scala 119:34]
  wire  _GEN_8351 = unuse_way == 2'h1 | _GEN_7323; // @[d_cache.scala 119:34 124:23]
  wire [63:0] _GEN_8352 = unuse_way == 2'h1 ? ram_1_0 : _GEN_6939; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8353 = unuse_way == 2'h1 ? ram_1_1 : _GEN_6940; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8354 = unuse_way == 2'h1 ? ram_1_2 : _GEN_6941; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8355 = unuse_way == 2'h1 ? ram_1_3 : _GEN_6942; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8356 = unuse_way == 2'h1 ? ram_1_4 : _GEN_6943; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8357 = unuse_way == 2'h1 ? ram_1_5 : _GEN_6944; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8358 = unuse_way == 2'h1 ? ram_1_6 : _GEN_6945; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8359 = unuse_way == 2'h1 ? ram_1_7 : _GEN_6946; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8360 = unuse_way == 2'h1 ? ram_1_8 : _GEN_6947; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8361 = unuse_way == 2'h1 ? ram_1_9 : _GEN_6948; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8362 = unuse_way == 2'h1 ? ram_1_10 : _GEN_6949; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8363 = unuse_way == 2'h1 ? ram_1_11 : _GEN_6950; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8364 = unuse_way == 2'h1 ? ram_1_12 : _GEN_6951; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8365 = unuse_way == 2'h1 ? ram_1_13 : _GEN_6952; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8366 = unuse_way == 2'h1 ? ram_1_14 : _GEN_6953; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8367 = unuse_way == 2'h1 ? ram_1_15 : _GEN_6954; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8368 = unuse_way == 2'h1 ? ram_1_16 : _GEN_6955; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8369 = unuse_way == 2'h1 ? ram_1_17 : _GEN_6956; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8370 = unuse_way == 2'h1 ? ram_1_18 : _GEN_6957; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8371 = unuse_way == 2'h1 ? ram_1_19 : _GEN_6958; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8372 = unuse_way == 2'h1 ? ram_1_20 : _GEN_6959; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8373 = unuse_way == 2'h1 ? ram_1_21 : _GEN_6960; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8374 = unuse_way == 2'h1 ? ram_1_22 : _GEN_6961; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8375 = unuse_way == 2'h1 ? ram_1_23 : _GEN_6962; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8376 = unuse_way == 2'h1 ? ram_1_24 : _GEN_6963; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8377 = unuse_way == 2'h1 ? ram_1_25 : _GEN_6964; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8378 = unuse_way == 2'h1 ? ram_1_26 : _GEN_6965; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8379 = unuse_way == 2'h1 ? ram_1_27 : _GEN_6966; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8380 = unuse_way == 2'h1 ? ram_1_28 : _GEN_6967; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8381 = unuse_way == 2'h1 ? ram_1_29 : _GEN_6968; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8382 = unuse_way == 2'h1 ? ram_1_30 : _GEN_6969; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8383 = unuse_way == 2'h1 ? ram_1_31 : _GEN_6970; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8384 = unuse_way == 2'h1 ? ram_1_32 : _GEN_6971; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8385 = unuse_way == 2'h1 ? ram_1_33 : _GEN_6972; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8386 = unuse_way == 2'h1 ? ram_1_34 : _GEN_6973; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8387 = unuse_way == 2'h1 ? ram_1_35 : _GEN_6974; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8388 = unuse_way == 2'h1 ? ram_1_36 : _GEN_6975; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8389 = unuse_way == 2'h1 ? ram_1_37 : _GEN_6976; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8390 = unuse_way == 2'h1 ? ram_1_38 : _GEN_6977; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8391 = unuse_way == 2'h1 ? ram_1_39 : _GEN_6978; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8392 = unuse_way == 2'h1 ? ram_1_40 : _GEN_6979; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8393 = unuse_way == 2'h1 ? ram_1_41 : _GEN_6980; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8394 = unuse_way == 2'h1 ? ram_1_42 : _GEN_6981; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8395 = unuse_way == 2'h1 ? ram_1_43 : _GEN_6982; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8396 = unuse_way == 2'h1 ? ram_1_44 : _GEN_6983; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8397 = unuse_way == 2'h1 ? ram_1_45 : _GEN_6984; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8398 = unuse_way == 2'h1 ? ram_1_46 : _GEN_6985; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8399 = unuse_way == 2'h1 ? ram_1_47 : _GEN_6986; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8400 = unuse_way == 2'h1 ? ram_1_48 : _GEN_6987; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8401 = unuse_way == 2'h1 ? ram_1_49 : _GEN_6988; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8402 = unuse_way == 2'h1 ? ram_1_50 : _GEN_6989; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8403 = unuse_way == 2'h1 ? ram_1_51 : _GEN_6990; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8404 = unuse_way == 2'h1 ? ram_1_52 : _GEN_6991; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8405 = unuse_way == 2'h1 ? ram_1_53 : _GEN_6992; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8406 = unuse_way == 2'h1 ? ram_1_54 : _GEN_6993; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8407 = unuse_way == 2'h1 ? ram_1_55 : _GEN_6994; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8408 = unuse_way == 2'h1 ? ram_1_56 : _GEN_6995; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8409 = unuse_way == 2'h1 ? ram_1_57 : _GEN_6996; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8410 = unuse_way == 2'h1 ? ram_1_58 : _GEN_6997; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8411 = unuse_way == 2'h1 ? ram_1_59 : _GEN_6998; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8412 = unuse_way == 2'h1 ? ram_1_60 : _GEN_6999; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8413 = unuse_way == 2'h1 ? ram_1_61 : _GEN_7000; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8414 = unuse_way == 2'h1 ? ram_1_62 : _GEN_7001; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8415 = unuse_way == 2'h1 ? ram_1_63 : _GEN_7002; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8416 = unuse_way == 2'h1 ? ram_1_64 : _GEN_7003; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8417 = unuse_way == 2'h1 ? ram_1_65 : _GEN_7004; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8418 = unuse_way == 2'h1 ? ram_1_66 : _GEN_7005; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8419 = unuse_way == 2'h1 ? ram_1_67 : _GEN_7006; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8420 = unuse_way == 2'h1 ? ram_1_68 : _GEN_7007; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8421 = unuse_way == 2'h1 ? ram_1_69 : _GEN_7008; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8422 = unuse_way == 2'h1 ? ram_1_70 : _GEN_7009; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8423 = unuse_way == 2'h1 ? ram_1_71 : _GEN_7010; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8424 = unuse_way == 2'h1 ? ram_1_72 : _GEN_7011; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8425 = unuse_way == 2'h1 ? ram_1_73 : _GEN_7012; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8426 = unuse_way == 2'h1 ? ram_1_74 : _GEN_7013; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8427 = unuse_way == 2'h1 ? ram_1_75 : _GEN_7014; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8428 = unuse_way == 2'h1 ? ram_1_76 : _GEN_7015; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8429 = unuse_way == 2'h1 ? ram_1_77 : _GEN_7016; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8430 = unuse_way == 2'h1 ? ram_1_78 : _GEN_7017; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8431 = unuse_way == 2'h1 ? ram_1_79 : _GEN_7018; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8432 = unuse_way == 2'h1 ? ram_1_80 : _GEN_7019; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8433 = unuse_way == 2'h1 ? ram_1_81 : _GEN_7020; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8434 = unuse_way == 2'h1 ? ram_1_82 : _GEN_7021; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8435 = unuse_way == 2'h1 ? ram_1_83 : _GEN_7022; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8436 = unuse_way == 2'h1 ? ram_1_84 : _GEN_7023; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8437 = unuse_way == 2'h1 ? ram_1_85 : _GEN_7024; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8438 = unuse_way == 2'h1 ? ram_1_86 : _GEN_7025; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8439 = unuse_way == 2'h1 ? ram_1_87 : _GEN_7026; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8440 = unuse_way == 2'h1 ? ram_1_88 : _GEN_7027; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8441 = unuse_way == 2'h1 ? ram_1_89 : _GEN_7028; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8442 = unuse_way == 2'h1 ? ram_1_90 : _GEN_7029; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8443 = unuse_way == 2'h1 ? ram_1_91 : _GEN_7030; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8444 = unuse_way == 2'h1 ? ram_1_92 : _GEN_7031; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8445 = unuse_way == 2'h1 ? ram_1_93 : _GEN_7032; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8446 = unuse_way == 2'h1 ? ram_1_94 : _GEN_7033; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8447 = unuse_way == 2'h1 ? ram_1_95 : _GEN_7034; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8448 = unuse_way == 2'h1 ? ram_1_96 : _GEN_7035; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8449 = unuse_way == 2'h1 ? ram_1_97 : _GEN_7036; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8450 = unuse_way == 2'h1 ? ram_1_98 : _GEN_7037; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8451 = unuse_way == 2'h1 ? ram_1_99 : _GEN_7038; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8452 = unuse_way == 2'h1 ? ram_1_100 : _GEN_7039; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8453 = unuse_way == 2'h1 ? ram_1_101 : _GEN_7040; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8454 = unuse_way == 2'h1 ? ram_1_102 : _GEN_7041; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8455 = unuse_way == 2'h1 ? ram_1_103 : _GEN_7042; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8456 = unuse_way == 2'h1 ? ram_1_104 : _GEN_7043; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8457 = unuse_way == 2'h1 ? ram_1_105 : _GEN_7044; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8458 = unuse_way == 2'h1 ? ram_1_106 : _GEN_7045; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8459 = unuse_way == 2'h1 ? ram_1_107 : _GEN_7046; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8460 = unuse_way == 2'h1 ? ram_1_108 : _GEN_7047; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8461 = unuse_way == 2'h1 ? ram_1_109 : _GEN_7048; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8462 = unuse_way == 2'h1 ? ram_1_110 : _GEN_7049; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8463 = unuse_way == 2'h1 ? ram_1_111 : _GEN_7050; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8464 = unuse_way == 2'h1 ? ram_1_112 : _GEN_7051; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8465 = unuse_way == 2'h1 ? ram_1_113 : _GEN_7052; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8466 = unuse_way == 2'h1 ? ram_1_114 : _GEN_7053; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8467 = unuse_way == 2'h1 ? ram_1_115 : _GEN_7054; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8468 = unuse_way == 2'h1 ? ram_1_116 : _GEN_7055; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8469 = unuse_way == 2'h1 ? ram_1_117 : _GEN_7056; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8470 = unuse_way == 2'h1 ? ram_1_118 : _GEN_7057; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8471 = unuse_way == 2'h1 ? ram_1_119 : _GEN_7058; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8472 = unuse_way == 2'h1 ? ram_1_120 : _GEN_7059; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8473 = unuse_way == 2'h1 ? ram_1_121 : _GEN_7060; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8474 = unuse_way == 2'h1 ? ram_1_122 : _GEN_7061; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8475 = unuse_way == 2'h1 ? ram_1_123 : _GEN_7062; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8476 = unuse_way == 2'h1 ? ram_1_124 : _GEN_7063; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8477 = unuse_way == 2'h1 ? ram_1_125 : _GEN_7064; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8478 = unuse_way == 2'h1 ? ram_1_126 : _GEN_7065; // @[d_cache.scala 119:34 19:24]
  wire [63:0] _GEN_8479 = unuse_way == 2'h1 ? ram_1_127 : _GEN_7066; // @[d_cache.scala 119:34 19:24]
  wire [31:0] _GEN_8480 = unuse_way == 2'h1 ? tag_1_0 : _GEN_7067; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8481 = unuse_way == 2'h1 ? tag_1_1 : _GEN_7068; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8482 = unuse_way == 2'h1 ? tag_1_2 : _GEN_7069; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8483 = unuse_way == 2'h1 ? tag_1_3 : _GEN_7070; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8484 = unuse_way == 2'h1 ? tag_1_4 : _GEN_7071; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8485 = unuse_way == 2'h1 ? tag_1_5 : _GEN_7072; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8486 = unuse_way == 2'h1 ? tag_1_6 : _GEN_7073; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8487 = unuse_way == 2'h1 ? tag_1_7 : _GEN_7074; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8488 = unuse_way == 2'h1 ? tag_1_8 : _GEN_7075; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8489 = unuse_way == 2'h1 ? tag_1_9 : _GEN_7076; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8490 = unuse_way == 2'h1 ? tag_1_10 : _GEN_7077; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8491 = unuse_way == 2'h1 ? tag_1_11 : _GEN_7078; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8492 = unuse_way == 2'h1 ? tag_1_12 : _GEN_7079; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8493 = unuse_way == 2'h1 ? tag_1_13 : _GEN_7080; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8494 = unuse_way == 2'h1 ? tag_1_14 : _GEN_7081; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8495 = unuse_way == 2'h1 ? tag_1_15 : _GEN_7082; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8496 = unuse_way == 2'h1 ? tag_1_16 : _GEN_7083; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8497 = unuse_way == 2'h1 ? tag_1_17 : _GEN_7084; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8498 = unuse_way == 2'h1 ? tag_1_18 : _GEN_7085; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8499 = unuse_way == 2'h1 ? tag_1_19 : _GEN_7086; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8500 = unuse_way == 2'h1 ? tag_1_20 : _GEN_7087; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8501 = unuse_way == 2'h1 ? tag_1_21 : _GEN_7088; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8502 = unuse_way == 2'h1 ? tag_1_22 : _GEN_7089; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8503 = unuse_way == 2'h1 ? tag_1_23 : _GEN_7090; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8504 = unuse_way == 2'h1 ? tag_1_24 : _GEN_7091; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8505 = unuse_way == 2'h1 ? tag_1_25 : _GEN_7092; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8506 = unuse_way == 2'h1 ? tag_1_26 : _GEN_7093; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8507 = unuse_way == 2'h1 ? tag_1_27 : _GEN_7094; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8508 = unuse_way == 2'h1 ? tag_1_28 : _GEN_7095; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8509 = unuse_way == 2'h1 ? tag_1_29 : _GEN_7096; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8510 = unuse_way == 2'h1 ? tag_1_30 : _GEN_7097; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8511 = unuse_way == 2'h1 ? tag_1_31 : _GEN_7098; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8512 = unuse_way == 2'h1 ? tag_1_32 : _GEN_7099; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8513 = unuse_way == 2'h1 ? tag_1_33 : _GEN_7100; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8514 = unuse_way == 2'h1 ? tag_1_34 : _GEN_7101; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8515 = unuse_way == 2'h1 ? tag_1_35 : _GEN_7102; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8516 = unuse_way == 2'h1 ? tag_1_36 : _GEN_7103; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8517 = unuse_way == 2'h1 ? tag_1_37 : _GEN_7104; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8518 = unuse_way == 2'h1 ? tag_1_38 : _GEN_7105; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8519 = unuse_way == 2'h1 ? tag_1_39 : _GEN_7106; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8520 = unuse_way == 2'h1 ? tag_1_40 : _GEN_7107; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8521 = unuse_way == 2'h1 ? tag_1_41 : _GEN_7108; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8522 = unuse_way == 2'h1 ? tag_1_42 : _GEN_7109; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8523 = unuse_way == 2'h1 ? tag_1_43 : _GEN_7110; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8524 = unuse_way == 2'h1 ? tag_1_44 : _GEN_7111; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8525 = unuse_way == 2'h1 ? tag_1_45 : _GEN_7112; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8526 = unuse_way == 2'h1 ? tag_1_46 : _GEN_7113; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8527 = unuse_way == 2'h1 ? tag_1_47 : _GEN_7114; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8528 = unuse_way == 2'h1 ? tag_1_48 : _GEN_7115; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8529 = unuse_way == 2'h1 ? tag_1_49 : _GEN_7116; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8530 = unuse_way == 2'h1 ? tag_1_50 : _GEN_7117; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8531 = unuse_way == 2'h1 ? tag_1_51 : _GEN_7118; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8532 = unuse_way == 2'h1 ? tag_1_52 : _GEN_7119; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8533 = unuse_way == 2'h1 ? tag_1_53 : _GEN_7120; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8534 = unuse_way == 2'h1 ? tag_1_54 : _GEN_7121; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8535 = unuse_way == 2'h1 ? tag_1_55 : _GEN_7122; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8536 = unuse_way == 2'h1 ? tag_1_56 : _GEN_7123; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8537 = unuse_way == 2'h1 ? tag_1_57 : _GEN_7124; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8538 = unuse_way == 2'h1 ? tag_1_58 : _GEN_7125; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8539 = unuse_way == 2'h1 ? tag_1_59 : _GEN_7126; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8540 = unuse_way == 2'h1 ? tag_1_60 : _GEN_7127; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8541 = unuse_way == 2'h1 ? tag_1_61 : _GEN_7128; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8542 = unuse_way == 2'h1 ? tag_1_62 : _GEN_7129; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8543 = unuse_way == 2'h1 ? tag_1_63 : _GEN_7130; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8544 = unuse_way == 2'h1 ? tag_1_64 : _GEN_7131; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8545 = unuse_way == 2'h1 ? tag_1_65 : _GEN_7132; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8546 = unuse_way == 2'h1 ? tag_1_66 : _GEN_7133; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8547 = unuse_way == 2'h1 ? tag_1_67 : _GEN_7134; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8548 = unuse_way == 2'h1 ? tag_1_68 : _GEN_7135; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8549 = unuse_way == 2'h1 ? tag_1_69 : _GEN_7136; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8550 = unuse_way == 2'h1 ? tag_1_70 : _GEN_7137; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8551 = unuse_way == 2'h1 ? tag_1_71 : _GEN_7138; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8552 = unuse_way == 2'h1 ? tag_1_72 : _GEN_7139; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8553 = unuse_way == 2'h1 ? tag_1_73 : _GEN_7140; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8554 = unuse_way == 2'h1 ? tag_1_74 : _GEN_7141; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8555 = unuse_way == 2'h1 ? tag_1_75 : _GEN_7142; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8556 = unuse_way == 2'h1 ? tag_1_76 : _GEN_7143; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8557 = unuse_way == 2'h1 ? tag_1_77 : _GEN_7144; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8558 = unuse_way == 2'h1 ? tag_1_78 : _GEN_7145; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8559 = unuse_way == 2'h1 ? tag_1_79 : _GEN_7146; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8560 = unuse_way == 2'h1 ? tag_1_80 : _GEN_7147; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8561 = unuse_way == 2'h1 ? tag_1_81 : _GEN_7148; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8562 = unuse_way == 2'h1 ? tag_1_82 : _GEN_7149; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8563 = unuse_way == 2'h1 ? tag_1_83 : _GEN_7150; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8564 = unuse_way == 2'h1 ? tag_1_84 : _GEN_7151; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8565 = unuse_way == 2'h1 ? tag_1_85 : _GEN_7152; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8566 = unuse_way == 2'h1 ? tag_1_86 : _GEN_7153; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8567 = unuse_way == 2'h1 ? tag_1_87 : _GEN_7154; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8568 = unuse_way == 2'h1 ? tag_1_88 : _GEN_7155; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8569 = unuse_way == 2'h1 ? tag_1_89 : _GEN_7156; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8570 = unuse_way == 2'h1 ? tag_1_90 : _GEN_7157; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8571 = unuse_way == 2'h1 ? tag_1_91 : _GEN_7158; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8572 = unuse_way == 2'h1 ? tag_1_92 : _GEN_7159; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8573 = unuse_way == 2'h1 ? tag_1_93 : _GEN_7160; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8574 = unuse_way == 2'h1 ? tag_1_94 : _GEN_7161; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8575 = unuse_way == 2'h1 ? tag_1_95 : _GEN_7162; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8576 = unuse_way == 2'h1 ? tag_1_96 : _GEN_7163; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8577 = unuse_way == 2'h1 ? tag_1_97 : _GEN_7164; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8578 = unuse_way == 2'h1 ? tag_1_98 : _GEN_7165; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8579 = unuse_way == 2'h1 ? tag_1_99 : _GEN_7166; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8580 = unuse_way == 2'h1 ? tag_1_100 : _GEN_7167; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8581 = unuse_way == 2'h1 ? tag_1_101 : _GEN_7168; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8582 = unuse_way == 2'h1 ? tag_1_102 : _GEN_7169; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8583 = unuse_way == 2'h1 ? tag_1_103 : _GEN_7170; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8584 = unuse_way == 2'h1 ? tag_1_104 : _GEN_7171; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8585 = unuse_way == 2'h1 ? tag_1_105 : _GEN_7172; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8586 = unuse_way == 2'h1 ? tag_1_106 : _GEN_7173; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8587 = unuse_way == 2'h1 ? tag_1_107 : _GEN_7174; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8588 = unuse_way == 2'h1 ? tag_1_108 : _GEN_7175; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8589 = unuse_way == 2'h1 ? tag_1_109 : _GEN_7176; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8590 = unuse_way == 2'h1 ? tag_1_110 : _GEN_7177; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8591 = unuse_way == 2'h1 ? tag_1_111 : _GEN_7178; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8592 = unuse_way == 2'h1 ? tag_1_112 : _GEN_7179; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8593 = unuse_way == 2'h1 ? tag_1_113 : _GEN_7180; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8594 = unuse_way == 2'h1 ? tag_1_114 : _GEN_7181; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8595 = unuse_way == 2'h1 ? tag_1_115 : _GEN_7182; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8596 = unuse_way == 2'h1 ? tag_1_116 : _GEN_7183; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8597 = unuse_way == 2'h1 ? tag_1_117 : _GEN_7184; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8598 = unuse_way == 2'h1 ? tag_1_118 : _GEN_7185; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8599 = unuse_way == 2'h1 ? tag_1_119 : _GEN_7186; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8600 = unuse_way == 2'h1 ? tag_1_120 : _GEN_7187; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8601 = unuse_way == 2'h1 ? tag_1_121 : _GEN_7188; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8602 = unuse_way == 2'h1 ? tag_1_122 : _GEN_7189; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8603 = unuse_way == 2'h1 ? tag_1_123 : _GEN_7190; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8604 = unuse_way == 2'h1 ? tag_1_124 : _GEN_7191; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8605 = unuse_way == 2'h1 ? tag_1_125 : _GEN_7192; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8606 = unuse_way == 2'h1 ? tag_1_126 : _GEN_7193; // @[d_cache.scala 119:34 21:24]
  wire [31:0] _GEN_8607 = unuse_way == 2'h1 ? tag_1_127 : _GEN_7194; // @[d_cache.scala 119:34 21:24]
  wire  _GEN_8608 = unuse_way == 2'h1 ? valid_1_0 : _GEN_7195; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8609 = unuse_way == 2'h1 ? valid_1_1 : _GEN_7196; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8610 = unuse_way == 2'h1 ? valid_1_2 : _GEN_7197; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8611 = unuse_way == 2'h1 ? valid_1_3 : _GEN_7198; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8612 = unuse_way == 2'h1 ? valid_1_4 : _GEN_7199; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8613 = unuse_way == 2'h1 ? valid_1_5 : _GEN_7200; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8614 = unuse_way == 2'h1 ? valid_1_6 : _GEN_7201; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8615 = unuse_way == 2'h1 ? valid_1_7 : _GEN_7202; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8616 = unuse_way == 2'h1 ? valid_1_8 : _GEN_7203; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8617 = unuse_way == 2'h1 ? valid_1_9 : _GEN_7204; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8618 = unuse_way == 2'h1 ? valid_1_10 : _GEN_7205; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8619 = unuse_way == 2'h1 ? valid_1_11 : _GEN_7206; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8620 = unuse_way == 2'h1 ? valid_1_12 : _GEN_7207; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8621 = unuse_way == 2'h1 ? valid_1_13 : _GEN_7208; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8622 = unuse_way == 2'h1 ? valid_1_14 : _GEN_7209; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8623 = unuse_way == 2'h1 ? valid_1_15 : _GEN_7210; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8624 = unuse_way == 2'h1 ? valid_1_16 : _GEN_7211; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8625 = unuse_way == 2'h1 ? valid_1_17 : _GEN_7212; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8626 = unuse_way == 2'h1 ? valid_1_18 : _GEN_7213; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8627 = unuse_way == 2'h1 ? valid_1_19 : _GEN_7214; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8628 = unuse_way == 2'h1 ? valid_1_20 : _GEN_7215; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8629 = unuse_way == 2'h1 ? valid_1_21 : _GEN_7216; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8630 = unuse_way == 2'h1 ? valid_1_22 : _GEN_7217; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8631 = unuse_way == 2'h1 ? valid_1_23 : _GEN_7218; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8632 = unuse_way == 2'h1 ? valid_1_24 : _GEN_7219; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8633 = unuse_way == 2'h1 ? valid_1_25 : _GEN_7220; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8634 = unuse_way == 2'h1 ? valid_1_26 : _GEN_7221; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8635 = unuse_way == 2'h1 ? valid_1_27 : _GEN_7222; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8636 = unuse_way == 2'h1 ? valid_1_28 : _GEN_7223; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8637 = unuse_way == 2'h1 ? valid_1_29 : _GEN_7224; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8638 = unuse_way == 2'h1 ? valid_1_30 : _GEN_7225; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8639 = unuse_way == 2'h1 ? valid_1_31 : _GEN_7226; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8640 = unuse_way == 2'h1 ? valid_1_32 : _GEN_7227; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8641 = unuse_way == 2'h1 ? valid_1_33 : _GEN_7228; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8642 = unuse_way == 2'h1 ? valid_1_34 : _GEN_7229; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8643 = unuse_way == 2'h1 ? valid_1_35 : _GEN_7230; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8644 = unuse_way == 2'h1 ? valid_1_36 : _GEN_7231; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8645 = unuse_way == 2'h1 ? valid_1_37 : _GEN_7232; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8646 = unuse_way == 2'h1 ? valid_1_38 : _GEN_7233; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8647 = unuse_way == 2'h1 ? valid_1_39 : _GEN_7234; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8648 = unuse_way == 2'h1 ? valid_1_40 : _GEN_7235; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8649 = unuse_way == 2'h1 ? valid_1_41 : _GEN_7236; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8650 = unuse_way == 2'h1 ? valid_1_42 : _GEN_7237; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8651 = unuse_way == 2'h1 ? valid_1_43 : _GEN_7238; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8652 = unuse_way == 2'h1 ? valid_1_44 : _GEN_7239; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8653 = unuse_way == 2'h1 ? valid_1_45 : _GEN_7240; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8654 = unuse_way == 2'h1 ? valid_1_46 : _GEN_7241; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8655 = unuse_way == 2'h1 ? valid_1_47 : _GEN_7242; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8656 = unuse_way == 2'h1 ? valid_1_48 : _GEN_7243; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8657 = unuse_way == 2'h1 ? valid_1_49 : _GEN_7244; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8658 = unuse_way == 2'h1 ? valid_1_50 : _GEN_7245; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8659 = unuse_way == 2'h1 ? valid_1_51 : _GEN_7246; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8660 = unuse_way == 2'h1 ? valid_1_52 : _GEN_7247; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8661 = unuse_way == 2'h1 ? valid_1_53 : _GEN_7248; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8662 = unuse_way == 2'h1 ? valid_1_54 : _GEN_7249; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8663 = unuse_way == 2'h1 ? valid_1_55 : _GEN_7250; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8664 = unuse_way == 2'h1 ? valid_1_56 : _GEN_7251; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8665 = unuse_way == 2'h1 ? valid_1_57 : _GEN_7252; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8666 = unuse_way == 2'h1 ? valid_1_58 : _GEN_7253; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8667 = unuse_way == 2'h1 ? valid_1_59 : _GEN_7254; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8668 = unuse_way == 2'h1 ? valid_1_60 : _GEN_7255; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8669 = unuse_way == 2'h1 ? valid_1_61 : _GEN_7256; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8670 = unuse_way == 2'h1 ? valid_1_62 : _GEN_7257; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8671 = unuse_way == 2'h1 ? valid_1_63 : _GEN_7258; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8672 = unuse_way == 2'h1 ? valid_1_64 : _GEN_7259; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8673 = unuse_way == 2'h1 ? valid_1_65 : _GEN_7260; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8674 = unuse_way == 2'h1 ? valid_1_66 : _GEN_7261; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8675 = unuse_way == 2'h1 ? valid_1_67 : _GEN_7262; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8676 = unuse_way == 2'h1 ? valid_1_68 : _GEN_7263; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8677 = unuse_way == 2'h1 ? valid_1_69 : _GEN_7264; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8678 = unuse_way == 2'h1 ? valid_1_70 : _GEN_7265; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8679 = unuse_way == 2'h1 ? valid_1_71 : _GEN_7266; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8680 = unuse_way == 2'h1 ? valid_1_72 : _GEN_7267; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8681 = unuse_way == 2'h1 ? valid_1_73 : _GEN_7268; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8682 = unuse_way == 2'h1 ? valid_1_74 : _GEN_7269; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8683 = unuse_way == 2'h1 ? valid_1_75 : _GEN_7270; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8684 = unuse_way == 2'h1 ? valid_1_76 : _GEN_7271; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8685 = unuse_way == 2'h1 ? valid_1_77 : _GEN_7272; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8686 = unuse_way == 2'h1 ? valid_1_78 : _GEN_7273; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8687 = unuse_way == 2'h1 ? valid_1_79 : _GEN_7274; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8688 = unuse_way == 2'h1 ? valid_1_80 : _GEN_7275; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8689 = unuse_way == 2'h1 ? valid_1_81 : _GEN_7276; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8690 = unuse_way == 2'h1 ? valid_1_82 : _GEN_7277; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8691 = unuse_way == 2'h1 ? valid_1_83 : _GEN_7278; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8692 = unuse_way == 2'h1 ? valid_1_84 : _GEN_7279; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8693 = unuse_way == 2'h1 ? valid_1_85 : _GEN_7280; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8694 = unuse_way == 2'h1 ? valid_1_86 : _GEN_7281; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8695 = unuse_way == 2'h1 ? valid_1_87 : _GEN_7282; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8696 = unuse_way == 2'h1 ? valid_1_88 : _GEN_7283; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8697 = unuse_way == 2'h1 ? valid_1_89 : _GEN_7284; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8698 = unuse_way == 2'h1 ? valid_1_90 : _GEN_7285; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8699 = unuse_way == 2'h1 ? valid_1_91 : _GEN_7286; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8700 = unuse_way == 2'h1 ? valid_1_92 : _GEN_7287; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8701 = unuse_way == 2'h1 ? valid_1_93 : _GEN_7288; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8702 = unuse_way == 2'h1 ? valid_1_94 : _GEN_7289; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8703 = unuse_way == 2'h1 ? valid_1_95 : _GEN_7290; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8704 = unuse_way == 2'h1 ? valid_1_96 : _GEN_7291; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8705 = unuse_way == 2'h1 ? valid_1_97 : _GEN_7292; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8706 = unuse_way == 2'h1 ? valid_1_98 : _GEN_7293; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8707 = unuse_way == 2'h1 ? valid_1_99 : _GEN_7294; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8708 = unuse_way == 2'h1 ? valid_1_100 : _GEN_7295; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8709 = unuse_way == 2'h1 ? valid_1_101 : _GEN_7296; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8710 = unuse_way == 2'h1 ? valid_1_102 : _GEN_7297; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8711 = unuse_way == 2'h1 ? valid_1_103 : _GEN_7298; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8712 = unuse_way == 2'h1 ? valid_1_104 : _GEN_7299; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8713 = unuse_way == 2'h1 ? valid_1_105 : _GEN_7300; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8714 = unuse_way == 2'h1 ? valid_1_106 : _GEN_7301; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8715 = unuse_way == 2'h1 ? valid_1_107 : _GEN_7302; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8716 = unuse_way == 2'h1 ? valid_1_108 : _GEN_7303; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8717 = unuse_way == 2'h1 ? valid_1_109 : _GEN_7304; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8718 = unuse_way == 2'h1 ? valid_1_110 : _GEN_7305; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8719 = unuse_way == 2'h1 ? valid_1_111 : _GEN_7306; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8720 = unuse_way == 2'h1 ? valid_1_112 : _GEN_7307; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8721 = unuse_way == 2'h1 ? valid_1_113 : _GEN_7308; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8722 = unuse_way == 2'h1 ? valid_1_114 : _GEN_7309; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8723 = unuse_way == 2'h1 ? valid_1_115 : _GEN_7310; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8724 = unuse_way == 2'h1 ? valid_1_116 : _GEN_7311; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8725 = unuse_way == 2'h1 ? valid_1_117 : _GEN_7312; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8726 = unuse_way == 2'h1 ? valid_1_118 : _GEN_7313; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8727 = unuse_way == 2'h1 ? valid_1_119 : _GEN_7314; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8728 = unuse_way == 2'h1 ? valid_1_120 : _GEN_7315; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8729 = unuse_way == 2'h1 ? valid_1_121 : _GEN_7316; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8730 = unuse_way == 2'h1 ? valid_1_122 : _GEN_7317; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8731 = unuse_way == 2'h1 ? valid_1_123 : _GEN_7318; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8732 = unuse_way == 2'h1 ? valid_1_124 : _GEN_7319; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8733 = unuse_way == 2'h1 ? valid_1_125 : _GEN_7320; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8734 = unuse_way == 2'h1 ? valid_1_126 : _GEN_7321; // @[d_cache.scala 119:34 23:26]
  wire  _GEN_8735 = unuse_way == 2'h1 ? valid_1_127 : _GEN_7322; // @[d_cache.scala 119:34 23:26]
  wire [63:0] _GEN_8736 = unuse_way == 2'h1 ? write_back_data : _GEN_7324; // @[d_cache.scala 119:34 29:34]
  wire [38:0] _GEN_8737 = unuse_way == 2'h1 ? {{7'd0}, write_back_addr} : _GEN_7325; // @[d_cache.scala 119:34 30:34]
  wire  _GEN_8738 = unuse_way == 2'h1 ? dirty_0_0 : _GEN_7582; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8739 = unuse_way == 2'h1 ? dirty_0_1 : _GEN_7583; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8740 = unuse_way == 2'h1 ? dirty_0_2 : _GEN_7584; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8741 = unuse_way == 2'h1 ? dirty_0_3 : _GEN_7585; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8742 = unuse_way == 2'h1 ? dirty_0_4 : _GEN_7586; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8743 = unuse_way == 2'h1 ? dirty_0_5 : _GEN_7587; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8744 = unuse_way == 2'h1 ? dirty_0_6 : _GEN_7588; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8745 = unuse_way == 2'h1 ? dirty_0_7 : _GEN_7589; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8746 = unuse_way == 2'h1 ? dirty_0_8 : _GEN_7590; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8747 = unuse_way == 2'h1 ? dirty_0_9 : _GEN_7591; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8748 = unuse_way == 2'h1 ? dirty_0_10 : _GEN_7592; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8749 = unuse_way == 2'h1 ? dirty_0_11 : _GEN_7593; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8750 = unuse_way == 2'h1 ? dirty_0_12 : _GEN_7594; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8751 = unuse_way == 2'h1 ? dirty_0_13 : _GEN_7595; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8752 = unuse_way == 2'h1 ? dirty_0_14 : _GEN_7596; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8753 = unuse_way == 2'h1 ? dirty_0_15 : _GEN_7597; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8754 = unuse_way == 2'h1 ? dirty_0_16 : _GEN_7598; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8755 = unuse_way == 2'h1 ? dirty_0_17 : _GEN_7599; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8756 = unuse_way == 2'h1 ? dirty_0_18 : _GEN_7600; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8757 = unuse_way == 2'h1 ? dirty_0_19 : _GEN_7601; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8758 = unuse_way == 2'h1 ? dirty_0_20 : _GEN_7602; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8759 = unuse_way == 2'h1 ? dirty_0_21 : _GEN_7603; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8760 = unuse_way == 2'h1 ? dirty_0_22 : _GEN_7604; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8761 = unuse_way == 2'h1 ? dirty_0_23 : _GEN_7605; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8762 = unuse_way == 2'h1 ? dirty_0_24 : _GEN_7606; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8763 = unuse_way == 2'h1 ? dirty_0_25 : _GEN_7607; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8764 = unuse_way == 2'h1 ? dirty_0_26 : _GEN_7608; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8765 = unuse_way == 2'h1 ? dirty_0_27 : _GEN_7609; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8766 = unuse_way == 2'h1 ? dirty_0_28 : _GEN_7610; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8767 = unuse_way == 2'h1 ? dirty_0_29 : _GEN_7611; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8768 = unuse_way == 2'h1 ? dirty_0_30 : _GEN_7612; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8769 = unuse_way == 2'h1 ? dirty_0_31 : _GEN_7613; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8770 = unuse_way == 2'h1 ? dirty_0_32 : _GEN_7614; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8771 = unuse_way == 2'h1 ? dirty_0_33 : _GEN_7615; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8772 = unuse_way == 2'h1 ? dirty_0_34 : _GEN_7616; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8773 = unuse_way == 2'h1 ? dirty_0_35 : _GEN_7617; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8774 = unuse_way == 2'h1 ? dirty_0_36 : _GEN_7618; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8775 = unuse_way == 2'h1 ? dirty_0_37 : _GEN_7619; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8776 = unuse_way == 2'h1 ? dirty_0_38 : _GEN_7620; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8777 = unuse_way == 2'h1 ? dirty_0_39 : _GEN_7621; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8778 = unuse_way == 2'h1 ? dirty_0_40 : _GEN_7622; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8779 = unuse_way == 2'h1 ? dirty_0_41 : _GEN_7623; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8780 = unuse_way == 2'h1 ? dirty_0_42 : _GEN_7624; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8781 = unuse_way == 2'h1 ? dirty_0_43 : _GEN_7625; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8782 = unuse_way == 2'h1 ? dirty_0_44 : _GEN_7626; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8783 = unuse_way == 2'h1 ? dirty_0_45 : _GEN_7627; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8784 = unuse_way == 2'h1 ? dirty_0_46 : _GEN_7628; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8785 = unuse_way == 2'h1 ? dirty_0_47 : _GEN_7629; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8786 = unuse_way == 2'h1 ? dirty_0_48 : _GEN_7630; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8787 = unuse_way == 2'h1 ? dirty_0_49 : _GEN_7631; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8788 = unuse_way == 2'h1 ? dirty_0_50 : _GEN_7632; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8789 = unuse_way == 2'h1 ? dirty_0_51 : _GEN_7633; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8790 = unuse_way == 2'h1 ? dirty_0_52 : _GEN_7634; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8791 = unuse_way == 2'h1 ? dirty_0_53 : _GEN_7635; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8792 = unuse_way == 2'h1 ? dirty_0_54 : _GEN_7636; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8793 = unuse_way == 2'h1 ? dirty_0_55 : _GEN_7637; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8794 = unuse_way == 2'h1 ? dirty_0_56 : _GEN_7638; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8795 = unuse_way == 2'h1 ? dirty_0_57 : _GEN_7639; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8796 = unuse_way == 2'h1 ? dirty_0_58 : _GEN_7640; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8797 = unuse_way == 2'h1 ? dirty_0_59 : _GEN_7641; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8798 = unuse_way == 2'h1 ? dirty_0_60 : _GEN_7642; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8799 = unuse_way == 2'h1 ? dirty_0_61 : _GEN_7643; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8800 = unuse_way == 2'h1 ? dirty_0_62 : _GEN_7644; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8801 = unuse_way == 2'h1 ? dirty_0_63 : _GEN_7645; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8802 = unuse_way == 2'h1 ? dirty_0_64 : _GEN_7646; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8803 = unuse_way == 2'h1 ? dirty_0_65 : _GEN_7647; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8804 = unuse_way == 2'h1 ? dirty_0_66 : _GEN_7648; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8805 = unuse_way == 2'h1 ? dirty_0_67 : _GEN_7649; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8806 = unuse_way == 2'h1 ? dirty_0_68 : _GEN_7650; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8807 = unuse_way == 2'h1 ? dirty_0_69 : _GEN_7651; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8808 = unuse_way == 2'h1 ? dirty_0_70 : _GEN_7652; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8809 = unuse_way == 2'h1 ? dirty_0_71 : _GEN_7653; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8810 = unuse_way == 2'h1 ? dirty_0_72 : _GEN_7654; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8811 = unuse_way == 2'h1 ? dirty_0_73 : _GEN_7655; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8812 = unuse_way == 2'h1 ? dirty_0_74 : _GEN_7656; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8813 = unuse_way == 2'h1 ? dirty_0_75 : _GEN_7657; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8814 = unuse_way == 2'h1 ? dirty_0_76 : _GEN_7658; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8815 = unuse_way == 2'h1 ? dirty_0_77 : _GEN_7659; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8816 = unuse_way == 2'h1 ? dirty_0_78 : _GEN_7660; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8817 = unuse_way == 2'h1 ? dirty_0_79 : _GEN_7661; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8818 = unuse_way == 2'h1 ? dirty_0_80 : _GEN_7662; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8819 = unuse_way == 2'h1 ? dirty_0_81 : _GEN_7663; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8820 = unuse_way == 2'h1 ? dirty_0_82 : _GEN_7664; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8821 = unuse_way == 2'h1 ? dirty_0_83 : _GEN_7665; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8822 = unuse_way == 2'h1 ? dirty_0_84 : _GEN_7666; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8823 = unuse_way == 2'h1 ? dirty_0_85 : _GEN_7667; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8824 = unuse_way == 2'h1 ? dirty_0_86 : _GEN_7668; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8825 = unuse_way == 2'h1 ? dirty_0_87 : _GEN_7669; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8826 = unuse_way == 2'h1 ? dirty_0_88 : _GEN_7670; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8827 = unuse_way == 2'h1 ? dirty_0_89 : _GEN_7671; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8828 = unuse_way == 2'h1 ? dirty_0_90 : _GEN_7672; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8829 = unuse_way == 2'h1 ? dirty_0_91 : _GEN_7673; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8830 = unuse_way == 2'h1 ? dirty_0_92 : _GEN_7674; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8831 = unuse_way == 2'h1 ? dirty_0_93 : _GEN_7675; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8832 = unuse_way == 2'h1 ? dirty_0_94 : _GEN_7676; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8833 = unuse_way == 2'h1 ? dirty_0_95 : _GEN_7677; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8834 = unuse_way == 2'h1 ? dirty_0_96 : _GEN_7678; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8835 = unuse_way == 2'h1 ? dirty_0_97 : _GEN_7679; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8836 = unuse_way == 2'h1 ? dirty_0_98 : _GEN_7680; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8837 = unuse_way == 2'h1 ? dirty_0_99 : _GEN_7681; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8838 = unuse_way == 2'h1 ? dirty_0_100 : _GEN_7682; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8839 = unuse_way == 2'h1 ? dirty_0_101 : _GEN_7683; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8840 = unuse_way == 2'h1 ? dirty_0_102 : _GEN_7684; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8841 = unuse_way == 2'h1 ? dirty_0_103 : _GEN_7685; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8842 = unuse_way == 2'h1 ? dirty_0_104 : _GEN_7686; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8843 = unuse_way == 2'h1 ? dirty_0_105 : _GEN_7687; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8844 = unuse_way == 2'h1 ? dirty_0_106 : _GEN_7688; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8845 = unuse_way == 2'h1 ? dirty_0_107 : _GEN_7689; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8846 = unuse_way == 2'h1 ? dirty_0_108 : _GEN_7690; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8847 = unuse_way == 2'h1 ? dirty_0_109 : _GEN_7691; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8848 = unuse_way == 2'h1 ? dirty_0_110 : _GEN_7692; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8849 = unuse_way == 2'h1 ? dirty_0_111 : _GEN_7693; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8850 = unuse_way == 2'h1 ? dirty_0_112 : _GEN_7694; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8851 = unuse_way == 2'h1 ? dirty_0_113 : _GEN_7695; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8852 = unuse_way == 2'h1 ? dirty_0_114 : _GEN_7696; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8853 = unuse_way == 2'h1 ? dirty_0_115 : _GEN_7697; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8854 = unuse_way == 2'h1 ? dirty_0_116 : _GEN_7698; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8855 = unuse_way == 2'h1 ? dirty_0_117 : _GEN_7699; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8856 = unuse_way == 2'h1 ? dirty_0_118 : _GEN_7700; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8857 = unuse_way == 2'h1 ? dirty_0_119 : _GEN_7701; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8858 = unuse_way == 2'h1 ? dirty_0_120 : _GEN_7702; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8859 = unuse_way == 2'h1 ? dirty_0_121 : _GEN_7703; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8860 = unuse_way == 2'h1 ? dirty_0_122 : _GEN_7704; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8861 = unuse_way == 2'h1 ? dirty_0_123 : _GEN_7705; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8862 = unuse_way == 2'h1 ? dirty_0_124 : _GEN_7706; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8863 = unuse_way == 2'h1 ? dirty_0_125 : _GEN_7707; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8864 = unuse_way == 2'h1 ? dirty_0_126 : _GEN_7708; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8865 = unuse_way == 2'h1 ? dirty_0_127 : _GEN_7709; // @[d_cache.scala 119:34 24:26]
  wire  _GEN_8866 = unuse_way == 2'h1 ? dirty_1_0 : _GEN_7838; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8867 = unuse_way == 2'h1 ? dirty_1_1 : _GEN_7839; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8868 = unuse_way == 2'h1 ? dirty_1_2 : _GEN_7840; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8869 = unuse_way == 2'h1 ? dirty_1_3 : _GEN_7841; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8870 = unuse_way == 2'h1 ? dirty_1_4 : _GEN_7842; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8871 = unuse_way == 2'h1 ? dirty_1_5 : _GEN_7843; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8872 = unuse_way == 2'h1 ? dirty_1_6 : _GEN_7844; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8873 = unuse_way == 2'h1 ? dirty_1_7 : _GEN_7845; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8874 = unuse_way == 2'h1 ? dirty_1_8 : _GEN_7846; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8875 = unuse_way == 2'h1 ? dirty_1_9 : _GEN_7847; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8876 = unuse_way == 2'h1 ? dirty_1_10 : _GEN_7848; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8877 = unuse_way == 2'h1 ? dirty_1_11 : _GEN_7849; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8878 = unuse_way == 2'h1 ? dirty_1_12 : _GEN_7850; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8879 = unuse_way == 2'h1 ? dirty_1_13 : _GEN_7851; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8880 = unuse_way == 2'h1 ? dirty_1_14 : _GEN_7852; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8881 = unuse_way == 2'h1 ? dirty_1_15 : _GEN_7853; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8882 = unuse_way == 2'h1 ? dirty_1_16 : _GEN_7854; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8883 = unuse_way == 2'h1 ? dirty_1_17 : _GEN_7855; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8884 = unuse_way == 2'h1 ? dirty_1_18 : _GEN_7856; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8885 = unuse_way == 2'h1 ? dirty_1_19 : _GEN_7857; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8886 = unuse_way == 2'h1 ? dirty_1_20 : _GEN_7858; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8887 = unuse_way == 2'h1 ? dirty_1_21 : _GEN_7859; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8888 = unuse_way == 2'h1 ? dirty_1_22 : _GEN_7860; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8889 = unuse_way == 2'h1 ? dirty_1_23 : _GEN_7861; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8890 = unuse_way == 2'h1 ? dirty_1_24 : _GEN_7862; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8891 = unuse_way == 2'h1 ? dirty_1_25 : _GEN_7863; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8892 = unuse_way == 2'h1 ? dirty_1_26 : _GEN_7864; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8893 = unuse_way == 2'h1 ? dirty_1_27 : _GEN_7865; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8894 = unuse_way == 2'h1 ? dirty_1_28 : _GEN_7866; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8895 = unuse_way == 2'h1 ? dirty_1_29 : _GEN_7867; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8896 = unuse_way == 2'h1 ? dirty_1_30 : _GEN_7868; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8897 = unuse_way == 2'h1 ? dirty_1_31 : _GEN_7869; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8898 = unuse_way == 2'h1 ? dirty_1_32 : _GEN_7870; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8899 = unuse_way == 2'h1 ? dirty_1_33 : _GEN_7871; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8900 = unuse_way == 2'h1 ? dirty_1_34 : _GEN_7872; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8901 = unuse_way == 2'h1 ? dirty_1_35 : _GEN_7873; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8902 = unuse_way == 2'h1 ? dirty_1_36 : _GEN_7874; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8903 = unuse_way == 2'h1 ? dirty_1_37 : _GEN_7875; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8904 = unuse_way == 2'h1 ? dirty_1_38 : _GEN_7876; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8905 = unuse_way == 2'h1 ? dirty_1_39 : _GEN_7877; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8906 = unuse_way == 2'h1 ? dirty_1_40 : _GEN_7878; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8907 = unuse_way == 2'h1 ? dirty_1_41 : _GEN_7879; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8908 = unuse_way == 2'h1 ? dirty_1_42 : _GEN_7880; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8909 = unuse_way == 2'h1 ? dirty_1_43 : _GEN_7881; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8910 = unuse_way == 2'h1 ? dirty_1_44 : _GEN_7882; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8911 = unuse_way == 2'h1 ? dirty_1_45 : _GEN_7883; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8912 = unuse_way == 2'h1 ? dirty_1_46 : _GEN_7884; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8913 = unuse_way == 2'h1 ? dirty_1_47 : _GEN_7885; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8914 = unuse_way == 2'h1 ? dirty_1_48 : _GEN_7886; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8915 = unuse_way == 2'h1 ? dirty_1_49 : _GEN_7887; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8916 = unuse_way == 2'h1 ? dirty_1_50 : _GEN_7888; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8917 = unuse_way == 2'h1 ? dirty_1_51 : _GEN_7889; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8918 = unuse_way == 2'h1 ? dirty_1_52 : _GEN_7890; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8919 = unuse_way == 2'h1 ? dirty_1_53 : _GEN_7891; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8920 = unuse_way == 2'h1 ? dirty_1_54 : _GEN_7892; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8921 = unuse_way == 2'h1 ? dirty_1_55 : _GEN_7893; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8922 = unuse_way == 2'h1 ? dirty_1_56 : _GEN_7894; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8923 = unuse_way == 2'h1 ? dirty_1_57 : _GEN_7895; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8924 = unuse_way == 2'h1 ? dirty_1_58 : _GEN_7896; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8925 = unuse_way == 2'h1 ? dirty_1_59 : _GEN_7897; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8926 = unuse_way == 2'h1 ? dirty_1_60 : _GEN_7898; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8927 = unuse_way == 2'h1 ? dirty_1_61 : _GEN_7899; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8928 = unuse_way == 2'h1 ? dirty_1_62 : _GEN_7900; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8929 = unuse_way == 2'h1 ? dirty_1_63 : _GEN_7901; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8930 = unuse_way == 2'h1 ? dirty_1_64 : _GEN_7902; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8931 = unuse_way == 2'h1 ? dirty_1_65 : _GEN_7903; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8932 = unuse_way == 2'h1 ? dirty_1_66 : _GEN_7904; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8933 = unuse_way == 2'h1 ? dirty_1_67 : _GEN_7905; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8934 = unuse_way == 2'h1 ? dirty_1_68 : _GEN_7906; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8935 = unuse_way == 2'h1 ? dirty_1_69 : _GEN_7907; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8936 = unuse_way == 2'h1 ? dirty_1_70 : _GEN_7908; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8937 = unuse_way == 2'h1 ? dirty_1_71 : _GEN_7909; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8938 = unuse_way == 2'h1 ? dirty_1_72 : _GEN_7910; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8939 = unuse_way == 2'h1 ? dirty_1_73 : _GEN_7911; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8940 = unuse_way == 2'h1 ? dirty_1_74 : _GEN_7912; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8941 = unuse_way == 2'h1 ? dirty_1_75 : _GEN_7913; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8942 = unuse_way == 2'h1 ? dirty_1_76 : _GEN_7914; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8943 = unuse_way == 2'h1 ? dirty_1_77 : _GEN_7915; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8944 = unuse_way == 2'h1 ? dirty_1_78 : _GEN_7916; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8945 = unuse_way == 2'h1 ? dirty_1_79 : _GEN_7917; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8946 = unuse_way == 2'h1 ? dirty_1_80 : _GEN_7918; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8947 = unuse_way == 2'h1 ? dirty_1_81 : _GEN_7919; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8948 = unuse_way == 2'h1 ? dirty_1_82 : _GEN_7920; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8949 = unuse_way == 2'h1 ? dirty_1_83 : _GEN_7921; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8950 = unuse_way == 2'h1 ? dirty_1_84 : _GEN_7922; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8951 = unuse_way == 2'h1 ? dirty_1_85 : _GEN_7923; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8952 = unuse_way == 2'h1 ? dirty_1_86 : _GEN_7924; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8953 = unuse_way == 2'h1 ? dirty_1_87 : _GEN_7925; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8954 = unuse_way == 2'h1 ? dirty_1_88 : _GEN_7926; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8955 = unuse_way == 2'h1 ? dirty_1_89 : _GEN_7927; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8956 = unuse_way == 2'h1 ? dirty_1_90 : _GEN_7928; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8957 = unuse_way == 2'h1 ? dirty_1_91 : _GEN_7929; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8958 = unuse_way == 2'h1 ? dirty_1_92 : _GEN_7930; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8959 = unuse_way == 2'h1 ? dirty_1_93 : _GEN_7931; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8960 = unuse_way == 2'h1 ? dirty_1_94 : _GEN_7932; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8961 = unuse_way == 2'h1 ? dirty_1_95 : _GEN_7933; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8962 = unuse_way == 2'h1 ? dirty_1_96 : _GEN_7934; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8963 = unuse_way == 2'h1 ? dirty_1_97 : _GEN_7935; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8964 = unuse_way == 2'h1 ? dirty_1_98 : _GEN_7936; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8965 = unuse_way == 2'h1 ? dirty_1_99 : _GEN_7937; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8966 = unuse_way == 2'h1 ? dirty_1_100 : _GEN_7938; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8967 = unuse_way == 2'h1 ? dirty_1_101 : _GEN_7939; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8968 = unuse_way == 2'h1 ? dirty_1_102 : _GEN_7940; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8969 = unuse_way == 2'h1 ? dirty_1_103 : _GEN_7941; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8970 = unuse_way == 2'h1 ? dirty_1_104 : _GEN_7942; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8971 = unuse_way == 2'h1 ? dirty_1_105 : _GEN_7943; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8972 = unuse_way == 2'h1 ? dirty_1_106 : _GEN_7944; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8973 = unuse_way == 2'h1 ? dirty_1_107 : _GEN_7945; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8974 = unuse_way == 2'h1 ? dirty_1_108 : _GEN_7946; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8975 = unuse_way == 2'h1 ? dirty_1_109 : _GEN_7947; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8976 = unuse_way == 2'h1 ? dirty_1_110 : _GEN_7948; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8977 = unuse_way == 2'h1 ? dirty_1_111 : _GEN_7949; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8978 = unuse_way == 2'h1 ? dirty_1_112 : _GEN_7950; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8979 = unuse_way == 2'h1 ? dirty_1_113 : _GEN_7951; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8980 = unuse_way == 2'h1 ? dirty_1_114 : _GEN_7952; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8981 = unuse_way == 2'h1 ? dirty_1_115 : _GEN_7953; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8982 = unuse_way == 2'h1 ? dirty_1_116 : _GEN_7954; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8983 = unuse_way == 2'h1 ? dirty_1_117 : _GEN_7955; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8984 = unuse_way == 2'h1 ? dirty_1_118 : _GEN_7956; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8985 = unuse_way == 2'h1 ? dirty_1_119 : _GEN_7957; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8986 = unuse_way == 2'h1 ? dirty_1_120 : _GEN_7958; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8987 = unuse_way == 2'h1 ? dirty_1_121 : _GEN_7959; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8988 = unuse_way == 2'h1 ? dirty_1_122 : _GEN_7960; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8989 = unuse_way == 2'h1 ? dirty_1_123 : _GEN_7961; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8990 = unuse_way == 2'h1 ? dirty_1_124 : _GEN_7962; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8991 = unuse_way == 2'h1 ? dirty_1_125 : _GEN_7963; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8992 = unuse_way == 2'h1 ? dirty_1_126 : _GEN_7964; // @[d_cache.scala 119:34 25:26]
  wire  _GEN_8993 = unuse_way == 2'h1 ? dirty_1_127 : _GEN_7965; // @[d_cache.scala 119:34 25:26]
  wire [2:0] _GEN_8994 = io_from_axi_bvalid ? 3'h5 : state; // @[d_cache.scala 171:37 172:23 60:24]
  wire [2:0] _GEN_8995 = 3'h7 == state ? 3'h1 : state; // @[d_cache.scala 64:18 176:19 60:24]
  wire [2:0] _GEN_8996 = 3'h6 == state ? _GEN_8994 : _GEN_8995; // @[d_cache.scala 64:18]
  wire [2:0] _GEN_8997 = 3'h5 == state ? _GEN_7966 : _GEN_8996; // @[d_cache.scala 64:18]
  wire [63:0] _GEN_8998 = 3'h5 == state ? _GEN_7967 : ram_0_0; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_8999 = 3'h5 == state ? _GEN_7968 : ram_0_1; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9000 = 3'h5 == state ? _GEN_7969 : ram_0_2; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9001 = 3'h5 == state ? _GEN_7970 : ram_0_3; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9002 = 3'h5 == state ? _GEN_7971 : ram_0_4; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9003 = 3'h5 == state ? _GEN_7972 : ram_0_5; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9004 = 3'h5 == state ? _GEN_7973 : ram_0_6; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9005 = 3'h5 == state ? _GEN_7974 : ram_0_7; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9006 = 3'h5 == state ? _GEN_7975 : ram_0_8; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9007 = 3'h5 == state ? _GEN_7976 : ram_0_9; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9008 = 3'h5 == state ? _GEN_7977 : ram_0_10; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9009 = 3'h5 == state ? _GEN_7978 : ram_0_11; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9010 = 3'h5 == state ? _GEN_7979 : ram_0_12; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9011 = 3'h5 == state ? _GEN_7980 : ram_0_13; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9012 = 3'h5 == state ? _GEN_7981 : ram_0_14; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9013 = 3'h5 == state ? _GEN_7982 : ram_0_15; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9014 = 3'h5 == state ? _GEN_7983 : ram_0_16; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9015 = 3'h5 == state ? _GEN_7984 : ram_0_17; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9016 = 3'h5 == state ? _GEN_7985 : ram_0_18; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9017 = 3'h5 == state ? _GEN_7986 : ram_0_19; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9018 = 3'h5 == state ? _GEN_7987 : ram_0_20; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9019 = 3'h5 == state ? _GEN_7988 : ram_0_21; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9020 = 3'h5 == state ? _GEN_7989 : ram_0_22; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9021 = 3'h5 == state ? _GEN_7990 : ram_0_23; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9022 = 3'h5 == state ? _GEN_7991 : ram_0_24; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9023 = 3'h5 == state ? _GEN_7992 : ram_0_25; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9024 = 3'h5 == state ? _GEN_7993 : ram_0_26; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9025 = 3'h5 == state ? _GEN_7994 : ram_0_27; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9026 = 3'h5 == state ? _GEN_7995 : ram_0_28; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9027 = 3'h5 == state ? _GEN_7996 : ram_0_29; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9028 = 3'h5 == state ? _GEN_7997 : ram_0_30; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9029 = 3'h5 == state ? _GEN_7998 : ram_0_31; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9030 = 3'h5 == state ? _GEN_7999 : ram_0_32; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9031 = 3'h5 == state ? _GEN_8000 : ram_0_33; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9032 = 3'h5 == state ? _GEN_8001 : ram_0_34; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9033 = 3'h5 == state ? _GEN_8002 : ram_0_35; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9034 = 3'h5 == state ? _GEN_8003 : ram_0_36; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9035 = 3'h5 == state ? _GEN_8004 : ram_0_37; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9036 = 3'h5 == state ? _GEN_8005 : ram_0_38; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9037 = 3'h5 == state ? _GEN_8006 : ram_0_39; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9038 = 3'h5 == state ? _GEN_8007 : ram_0_40; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9039 = 3'h5 == state ? _GEN_8008 : ram_0_41; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9040 = 3'h5 == state ? _GEN_8009 : ram_0_42; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9041 = 3'h5 == state ? _GEN_8010 : ram_0_43; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9042 = 3'h5 == state ? _GEN_8011 : ram_0_44; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9043 = 3'h5 == state ? _GEN_8012 : ram_0_45; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9044 = 3'h5 == state ? _GEN_8013 : ram_0_46; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9045 = 3'h5 == state ? _GEN_8014 : ram_0_47; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9046 = 3'h5 == state ? _GEN_8015 : ram_0_48; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9047 = 3'h5 == state ? _GEN_8016 : ram_0_49; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9048 = 3'h5 == state ? _GEN_8017 : ram_0_50; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9049 = 3'h5 == state ? _GEN_8018 : ram_0_51; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9050 = 3'h5 == state ? _GEN_8019 : ram_0_52; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9051 = 3'h5 == state ? _GEN_8020 : ram_0_53; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9052 = 3'h5 == state ? _GEN_8021 : ram_0_54; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9053 = 3'h5 == state ? _GEN_8022 : ram_0_55; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9054 = 3'h5 == state ? _GEN_8023 : ram_0_56; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9055 = 3'h5 == state ? _GEN_8024 : ram_0_57; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9056 = 3'h5 == state ? _GEN_8025 : ram_0_58; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9057 = 3'h5 == state ? _GEN_8026 : ram_0_59; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9058 = 3'h5 == state ? _GEN_8027 : ram_0_60; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9059 = 3'h5 == state ? _GEN_8028 : ram_0_61; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9060 = 3'h5 == state ? _GEN_8029 : ram_0_62; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9061 = 3'h5 == state ? _GEN_8030 : ram_0_63; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9062 = 3'h5 == state ? _GEN_8031 : ram_0_64; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9063 = 3'h5 == state ? _GEN_8032 : ram_0_65; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9064 = 3'h5 == state ? _GEN_8033 : ram_0_66; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9065 = 3'h5 == state ? _GEN_8034 : ram_0_67; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9066 = 3'h5 == state ? _GEN_8035 : ram_0_68; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9067 = 3'h5 == state ? _GEN_8036 : ram_0_69; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9068 = 3'h5 == state ? _GEN_8037 : ram_0_70; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9069 = 3'h5 == state ? _GEN_8038 : ram_0_71; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9070 = 3'h5 == state ? _GEN_8039 : ram_0_72; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9071 = 3'h5 == state ? _GEN_8040 : ram_0_73; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9072 = 3'h5 == state ? _GEN_8041 : ram_0_74; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9073 = 3'h5 == state ? _GEN_8042 : ram_0_75; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9074 = 3'h5 == state ? _GEN_8043 : ram_0_76; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9075 = 3'h5 == state ? _GEN_8044 : ram_0_77; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9076 = 3'h5 == state ? _GEN_8045 : ram_0_78; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9077 = 3'h5 == state ? _GEN_8046 : ram_0_79; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9078 = 3'h5 == state ? _GEN_8047 : ram_0_80; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9079 = 3'h5 == state ? _GEN_8048 : ram_0_81; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9080 = 3'h5 == state ? _GEN_8049 : ram_0_82; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9081 = 3'h5 == state ? _GEN_8050 : ram_0_83; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9082 = 3'h5 == state ? _GEN_8051 : ram_0_84; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9083 = 3'h5 == state ? _GEN_8052 : ram_0_85; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9084 = 3'h5 == state ? _GEN_8053 : ram_0_86; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9085 = 3'h5 == state ? _GEN_8054 : ram_0_87; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9086 = 3'h5 == state ? _GEN_8055 : ram_0_88; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9087 = 3'h5 == state ? _GEN_8056 : ram_0_89; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9088 = 3'h5 == state ? _GEN_8057 : ram_0_90; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9089 = 3'h5 == state ? _GEN_8058 : ram_0_91; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9090 = 3'h5 == state ? _GEN_8059 : ram_0_92; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9091 = 3'h5 == state ? _GEN_8060 : ram_0_93; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9092 = 3'h5 == state ? _GEN_8061 : ram_0_94; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9093 = 3'h5 == state ? _GEN_8062 : ram_0_95; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9094 = 3'h5 == state ? _GEN_8063 : ram_0_96; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9095 = 3'h5 == state ? _GEN_8064 : ram_0_97; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9096 = 3'h5 == state ? _GEN_8065 : ram_0_98; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9097 = 3'h5 == state ? _GEN_8066 : ram_0_99; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9098 = 3'h5 == state ? _GEN_8067 : ram_0_100; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9099 = 3'h5 == state ? _GEN_8068 : ram_0_101; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9100 = 3'h5 == state ? _GEN_8069 : ram_0_102; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9101 = 3'h5 == state ? _GEN_8070 : ram_0_103; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9102 = 3'h5 == state ? _GEN_8071 : ram_0_104; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9103 = 3'h5 == state ? _GEN_8072 : ram_0_105; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9104 = 3'h5 == state ? _GEN_8073 : ram_0_106; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9105 = 3'h5 == state ? _GEN_8074 : ram_0_107; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9106 = 3'h5 == state ? _GEN_8075 : ram_0_108; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9107 = 3'h5 == state ? _GEN_8076 : ram_0_109; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9108 = 3'h5 == state ? _GEN_8077 : ram_0_110; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9109 = 3'h5 == state ? _GEN_8078 : ram_0_111; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9110 = 3'h5 == state ? _GEN_8079 : ram_0_112; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9111 = 3'h5 == state ? _GEN_8080 : ram_0_113; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9112 = 3'h5 == state ? _GEN_8081 : ram_0_114; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9113 = 3'h5 == state ? _GEN_8082 : ram_0_115; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9114 = 3'h5 == state ? _GEN_8083 : ram_0_116; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9115 = 3'h5 == state ? _GEN_8084 : ram_0_117; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9116 = 3'h5 == state ? _GEN_8085 : ram_0_118; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9117 = 3'h5 == state ? _GEN_8086 : ram_0_119; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9118 = 3'h5 == state ? _GEN_8087 : ram_0_120; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9119 = 3'h5 == state ? _GEN_8088 : ram_0_121; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9120 = 3'h5 == state ? _GEN_8089 : ram_0_122; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9121 = 3'h5 == state ? _GEN_8090 : ram_0_123; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9122 = 3'h5 == state ? _GEN_8091 : ram_0_124; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9123 = 3'h5 == state ? _GEN_8092 : ram_0_125; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9124 = 3'h5 == state ? _GEN_8093 : ram_0_126; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_9125 = 3'h5 == state ? _GEN_8094 : ram_0_127; // @[d_cache.scala 64:18 18:24]
  wire [31:0] _GEN_9126 = 3'h5 == state ? _GEN_8095 : tag_0_0; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9127 = 3'h5 == state ? _GEN_8096 : tag_0_1; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9128 = 3'h5 == state ? _GEN_8097 : tag_0_2; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9129 = 3'h5 == state ? _GEN_8098 : tag_0_3; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9130 = 3'h5 == state ? _GEN_8099 : tag_0_4; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9131 = 3'h5 == state ? _GEN_8100 : tag_0_5; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9132 = 3'h5 == state ? _GEN_8101 : tag_0_6; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9133 = 3'h5 == state ? _GEN_8102 : tag_0_7; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9134 = 3'h5 == state ? _GEN_8103 : tag_0_8; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9135 = 3'h5 == state ? _GEN_8104 : tag_0_9; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9136 = 3'h5 == state ? _GEN_8105 : tag_0_10; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9137 = 3'h5 == state ? _GEN_8106 : tag_0_11; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9138 = 3'h5 == state ? _GEN_8107 : tag_0_12; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9139 = 3'h5 == state ? _GEN_8108 : tag_0_13; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9140 = 3'h5 == state ? _GEN_8109 : tag_0_14; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9141 = 3'h5 == state ? _GEN_8110 : tag_0_15; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9142 = 3'h5 == state ? _GEN_8111 : tag_0_16; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9143 = 3'h5 == state ? _GEN_8112 : tag_0_17; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9144 = 3'h5 == state ? _GEN_8113 : tag_0_18; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9145 = 3'h5 == state ? _GEN_8114 : tag_0_19; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9146 = 3'h5 == state ? _GEN_8115 : tag_0_20; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9147 = 3'h5 == state ? _GEN_8116 : tag_0_21; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9148 = 3'h5 == state ? _GEN_8117 : tag_0_22; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9149 = 3'h5 == state ? _GEN_8118 : tag_0_23; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9150 = 3'h5 == state ? _GEN_8119 : tag_0_24; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9151 = 3'h5 == state ? _GEN_8120 : tag_0_25; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9152 = 3'h5 == state ? _GEN_8121 : tag_0_26; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9153 = 3'h5 == state ? _GEN_8122 : tag_0_27; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9154 = 3'h5 == state ? _GEN_8123 : tag_0_28; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9155 = 3'h5 == state ? _GEN_8124 : tag_0_29; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9156 = 3'h5 == state ? _GEN_8125 : tag_0_30; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9157 = 3'h5 == state ? _GEN_8126 : tag_0_31; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9158 = 3'h5 == state ? _GEN_8127 : tag_0_32; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9159 = 3'h5 == state ? _GEN_8128 : tag_0_33; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9160 = 3'h5 == state ? _GEN_8129 : tag_0_34; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9161 = 3'h5 == state ? _GEN_8130 : tag_0_35; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9162 = 3'h5 == state ? _GEN_8131 : tag_0_36; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9163 = 3'h5 == state ? _GEN_8132 : tag_0_37; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9164 = 3'h5 == state ? _GEN_8133 : tag_0_38; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9165 = 3'h5 == state ? _GEN_8134 : tag_0_39; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9166 = 3'h5 == state ? _GEN_8135 : tag_0_40; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9167 = 3'h5 == state ? _GEN_8136 : tag_0_41; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9168 = 3'h5 == state ? _GEN_8137 : tag_0_42; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9169 = 3'h5 == state ? _GEN_8138 : tag_0_43; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9170 = 3'h5 == state ? _GEN_8139 : tag_0_44; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9171 = 3'h5 == state ? _GEN_8140 : tag_0_45; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9172 = 3'h5 == state ? _GEN_8141 : tag_0_46; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9173 = 3'h5 == state ? _GEN_8142 : tag_0_47; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9174 = 3'h5 == state ? _GEN_8143 : tag_0_48; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9175 = 3'h5 == state ? _GEN_8144 : tag_0_49; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9176 = 3'h5 == state ? _GEN_8145 : tag_0_50; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9177 = 3'h5 == state ? _GEN_8146 : tag_0_51; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9178 = 3'h5 == state ? _GEN_8147 : tag_0_52; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9179 = 3'h5 == state ? _GEN_8148 : tag_0_53; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9180 = 3'h5 == state ? _GEN_8149 : tag_0_54; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9181 = 3'h5 == state ? _GEN_8150 : tag_0_55; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9182 = 3'h5 == state ? _GEN_8151 : tag_0_56; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9183 = 3'h5 == state ? _GEN_8152 : tag_0_57; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9184 = 3'h5 == state ? _GEN_8153 : tag_0_58; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9185 = 3'h5 == state ? _GEN_8154 : tag_0_59; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9186 = 3'h5 == state ? _GEN_8155 : tag_0_60; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9187 = 3'h5 == state ? _GEN_8156 : tag_0_61; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9188 = 3'h5 == state ? _GEN_8157 : tag_0_62; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9189 = 3'h5 == state ? _GEN_8158 : tag_0_63; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9190 = 3'h5 == state ? _GEN_8159 : tag_0_64; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9191 = 3'h5 == state ? _GEN_8160 : tag_0_65; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9192 = 3'h5 == state ? _GEN_8161 : tag_0_66; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9193 = 3'h5 == state ? _GEN_8162 : tag_0_67; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9194 = 3'h5 == state ? _GEN_8163 : tag_0_68; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9195 = 3'h5 == state ? _GEN_8164 : tag_0_69; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9196 = 3'h5 == state ? _GEN_8165 : tag_0_70; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9197 = 3'h5 == state ? _GEN_8166 : tag_0_71; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9198 = 3'h5 == state ? _GEN_8167 : tag_0_72; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9199 = 3'h5 == state ? _GEN_8168 : tag_0_73; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9200 = 3'h5 == state ? _GEN_8169 : tag_0_74; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9201 = 3'h5 == state ? _GEN_8170 : tag_0_75; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9202 = 3'h5 == state ? _GEN_8171 : tag_0_76; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9203 = 3'h5 == state ? _GEN_8172 : tag_0_77; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9204 = 3'h5 == state ? _GEN_8173 : tag_0_78; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9205 = 3'h5 == state ? _GEN_8174 : tag_0_79; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9206 = 3'h5 == state ? _GEN_8175 : tag_0_80; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9207 = 3'h5 == state ? _GEN_8176 : tag_0_81; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9208 = 3'h5 == state ? _GEN_8177 : tag_0_82; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9209 = 3'h5 == state ? _GEN_8178 : tag_0_83; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9210 = 3'h5 == state ? _GEN_8179 : tag_0_84; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9211 = 3'h5 == state ? _GEN_8180 : tag_0_85; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9212 = 3'h5 == state ? _GEN_8181 : tag_0_86; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9213 = 3'h5 == state ? _GEN_8182 : tag_0_87; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9214 = 3'h5 == state ? _GEN_8183 : tag_0_88; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9215 = 3'h5 == state ? _GEN_8184 : tag_0_89; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9216 = 3'h5 == state ? _GEN_8185 : tag_0_90; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9217 = 3'h5 == state ? _GEN_8186 : tag_0_91; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9218 = 3'h5 == state ? _GEN_8187 : tag_0_92; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9219 = 3'h5 == state ? _GEN_8188 : tag_0_93; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9220 = 3'h5 == state ? _GEN_8189 : tag_0_94; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9221 = 3'h5 == state ? _GEN_8190 : tag_0_95; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9222 = 3'h5 == state ? _GEN_8191 : tag_0_96; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9223 = 3'h5 == state ? _GEN_8192 : tag_0_97; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9224 = 3'h5 == state ? _GEN_8193 : tag_0_98; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9225 = 3'h5 == state ? _GEN_8194 : tag_0_99; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9226 = 3'h5 == state ? _GEN_8195 : tag_0_100; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9227 = 3'h5 == state ? _GEN_8196 : tag_0_101; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9228 = 3'h5 == state ? _GEN_8197 : tag_0_102; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9229 = 3'h5 == state ? _GEN_8198 : tag_0_103; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9230 = 3'h5 == state ? _GEN_8199 : tag_0_104; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9231 = 3'h5 == state ? _GEN_8200 : tag_0_105; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9232 = 3'h5 == state ? _GEN_8201 : tag_0_106; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9233 = 3'h5 == state ? _GEN_8202 : tag_0_107; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9234 = 3'h5 == state ? _GEN_8203 : tag_0_108; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9235 = 3'h5 == state ? _GEN_8204 : tag_0_109; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9236 = 3'h5 == state ? _GEN_8205 : tag_0_110; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9237 = 3'h5 == state ? _GEN_8206 : tag_0_111; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9238 = 3'h5 == state ? _GEN_8207 : tag_0_112; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9239 = 3'h5 == state ? _GEN_8208 : tag_0_113; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9240 = 3'h5 == state ? _GEN_8209 : tag_0_114; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9241 = 3'h5 == state ? _GEN_8210 : tag_0_115; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9242 = 3'h5 == state ? _GEN_8211 : tag_0_116; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9243 = 3'h5 == state ? _GEN_8212 : tag_0_117; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9244 = 3'h5 == state ? _GEN_8213 : tag_0_118; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9245 = 3'h5 == state ? _GEN_8214 : tag_0_119; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9246 = 3'h5 == state ? _GEN_8215 : tag_0_120; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9247 = 3'h5 == state ? _GEN_8216 : tag_0_121; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9248 = 3'h5 == state ? _GEN_8217 : tag_0_122; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9249 = 3'h5 == state ? _GEN_8218 : tag_0_123; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9250 = 3'h5 == state ? _GEN_8219 : tag_0_124; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9251 = 3'h5 == state ? _GEN_8220 : tag_0_125; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9252 = 3'h5 == state ? _GEN_8221 : tag_0_126; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_9253 = 3'h5 == state ? _GEN_8222 : tag_0_127; // @[d_cache.scala 64:18 20:24]
  wire  _GEN_9254 = 3'h5 == state ? _GEN_8223 : valid_0_0; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9255 = 3'h5 == state ? _GEN_8224 : valid_0_1; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9256 = 3'h5 == state ? _GEN_8225 : valid_0_2; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9257 = 3'h5 == state ? _GEN_8226 : valid_0_3; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9258 = 3'h5 == state ? _GEN_8227 : valid_0_4; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9259 = 3'h5 == state ? _GEN_8228 : valid_0_5; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9260 = 3'h5 == state ? _GEN_8229 : valid_0_6; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9261 = 3'h5 == state ? _GEN_8230 : valid_0_7; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9262 = 3'h5 == state ? _GEN_8231 : valid_0_8; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9263 = 3'h5 == state ? _GEN_8232 : valid_0_9; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9264 = 3'h5 == state ? _GEN_8233 : valid_0_10; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9265 = 3'h5 == state ? _GEN_8234 : valid_0_11; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9266 = 3'h5 == state ? _GEN_8235 : valid_0_12; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9267 = 3'h5 == state ? _GEN_8236 : valid_0_13; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9268 = 3'h5 == state ? _GEN_8237 : valid_0_14; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9269 = 3'h5 == state ? _GEN_8238 : valid_0_15; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9270 = 3'h5 == state ? _GEN_8239 : valid_0_16; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9271 = 3'h5 == state ? _GEN_8240 : valid_0_17; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9272 = 3'h5 == state ? _GEN_8241 : valid_0_18; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9273 = 3'h5 == state ? _GEN_8242 : valid_0_19; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9274 = 3'h5 == state ? _GEN_8243 : valid_0_20; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9275 = 3'h5 == state ? _GEN_8244 : valid_0_21; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9276 = 3'h5 == state ? _GEN_8245 : valid_0_22; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9277 = 3'h5 == state ? _GEN_8246 : valid_0_23; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9278 = 3'h5 == state ? _GEN_8247 : valid_0_24; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9279 = 3'h5 == state ? _GEN_8248 : valid_0_25; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9280 = 3'h5 == state ? _GEN_8249 : valid_0_26; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9281 = 3'h5 == state ? _GEN_8250 : valid_0_27; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9282 = 3'h5 == state ? _GEN_8251 : valid_0_28; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9283 = 3'h5 == state ? _GEN_8252 : valid_0_29; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9284 = 3'h5 == state ? _GEN_8253 : valid_0_30; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9285 = 3'h5 == state ? _GEN_8254 : valid_0_31; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9286 = 3'h5 == state ? _GEN_8255 : valid_0_32; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9287 = 3'h5 == state ? _GEN_8256 : valid_0_33; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9288 = 3'h5 == state ? _GEN_8257 : valid_0_34; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9289 = 3'h5 == state ? _GEN_8258 : valid_0_35; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9290 = 3'h5 == state ? _GEN_8259 : valid_0_36; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9291 = 3'h5 == state ? _GEN_8260 : valid_0_37; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9292 = 3'h5 == state ? _GEN_8261 : valid_0_38; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9293 = 3'h5 == state ? _GEN_8262 : valid_0_39; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9294 = 3'h5 == state ? _GEN_8263 : valid_0_40; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9295 = 3'h5 == state ? _GEN_8264 : valid_0_41; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9296 = 3'h5 == state ? _GEN_8265 : valid_0_42; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9297 = 3'h5 == state ? _GEN_8266 : valid_0_43; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9298 = 3'h5 == state ? _GEN_8267 : valid_0_44; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9299 = 3'h5 == state ? _GEN_8268 : valid_0_45; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9300 = 3'h5 == state ? _GEN_8269 : valid_0_46; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9301 = 3'h5 == state ? _GEN_8270 : valid_0_47; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9302 = 3'h5 == state ? _GEN_8271 : valid_0_48; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9303 = 3'h5 == state ? _GEN_8272 : valid_0_49; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9304 = 3'h5 == state ? _GEN_8273 : valid_0_50; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9305 = 3'h5 == state ? _GEN_8274 : valid_0_51; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9306 = 3'h5 == state ? _GEN_8275 : valid_0_52; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9307 = 3'h5 == state ? _GEN_8276 : valid_0_53; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9308 = 3'h5 == state ? _GEN_8277 : valid_0_54; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9309 = 3'h5 == state ? _GEN_8278 : valid_0_55; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9310 = 3'h5 == state ? _GEN_8279 : valid_0_56; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9311 = 3'h5 == state ? _GEN_8280 : valid_0_57; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9312 = 3'h5 == state ? _GEN_8281 : valid_0_58; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9313 = 3'h5 == state ? _GEN_8282 : valid_0_59; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9314 = 3'h5 == state ? _GEN_8283 : valid_0_60; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9315 = 3'h5 == state ? _GEN_8284 : valid_0_61; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9316 = 3'h5 == state ? _GEN_8285 : valid_0_62; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9317 = 3'h5 == state ? _GEN_8286 : valid_0_63; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9318 = 3'h5 == state ? _GEN_8287 : valid_0_64; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9319 = 3'h5 == state ? _GEN_8288 : valid_0_65; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9320 = 3'h5 == state ? _GEN_8289 : valid_0_66; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9321 = 3'h5 == state ? _GEN_8290 : valid_0_67; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9322 = 3'h5 == state ? _GEN_8291 : valid_0_68; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9323 = 3'h5 == state ? _GEN_8292 : valid_0_69; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9324 = 3'h5 == state ? _GEN_8293 : valid_0_70; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9325 = 3'h5 == state ? _GEN_8294 : valid_0_71; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9326 = 3'h5 == state ? _GEN_8295 : valid_0_72; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9327 = 3'h5 == state ? _GEN_8296 : valid_0_73; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9328 = 3'h5 == state ? _GEN_8297 : valid_0_74; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9329 = 3'h5 == state ? _GEN_8298 : valid_0_75; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9330 = 3'h5 == state ? _GEN_8299 : valid_0_76; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9331 = 3'h5 == state ? _GEN_8300 : valid_0_77; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9332 = 3'h5 == state ? _GEN_8301 : valid_0_78; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9333 = 3'h5 == state ? _GEN_8302 : valid_0_79; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9334 = 3'h5 == state ? _GEN_8303 : valid_0_80; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9335 = 3'h5 == state ? _GEN_8304 : valid_0_81; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9336 = 3'h5 == state ? _GEN_8305 : valid_0_82; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9337 = 3'h5 == state ? _GEN_8306 : valid_0_83; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9338 = 3'h5 == state ? _GEN_8307 : valid_0_84; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9339 = 3'h5 == state ? _GEN_8308 : valid_0_85; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9340 = 3'h5 == state ? _GEN_8309 : valid_0_86; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9341 = 3'h5 == state ? _GEN_8310 : valid_0_87; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9342 = 3'h5 == state ? _GEN_8311 : valid_0_88; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9343 = 3'h5 == state ? _GEN_8312 : valid_0_89; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9344 = 3'h5 == state ? _GEN_8313 : valid_0_90; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9345 = 3'h5 == state ? _GEN_8314 : valid_0_91; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9346 = 3'h5 == state ? _GEN_8315 : valid_0_92; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9347 = 3'h5 == state ? _GEN_8316 : valid_0_93; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9348 = 3'h5 == state ? _GEN_8317 : valid_0_94; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9349 = 3'h5 == state ? _GEN_8318 : valid_0_95; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9350 = 3'h5 == state ? _GEN_8319 : valid_0_96; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9351 = 3'h5 == state ? _GEN_8320 : valid_0_97; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9352 = 3'h5 == state ? _GEN_8321 : valid_0_98; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9353 = 3'h5 == state ? _GEN_8322 : valid_0_99; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9354 = 3'h5 == state ? _GEN_8323 : valid_0_100; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9355 = 3'h5 == state ? _GEN_8324 : valid_0_101; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9356 = 3'h5 == state ? _GEN_8325 : valid_0_102; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9357 = 3'h5 == state ? _GEN_8326 : valid_0_103; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9358 = 3'h5 == state ? _GEN_8327 : valid_0_104; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9359 = 3'h5 == state ? _GEN_8328 : valid_0_105; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9360 = 3'h5 == state ? _GEN_8329 : valid_0_106; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9361 = 3'h5 == state ? _GEN_8330 : valid_0_107; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9362 = 3'h5 == state ? _GEN_8331 : valid_0_108; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9363 = 3'h5 == state ? _GEN_8332 : valid_0_109; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9364 = 3'h5 == state ? _GEN_8333 : valid_0_110; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9365 = 3'h5 == state ? _GEN_8334 : valid_0_111; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9366 = 3'h5 == state ? _GEN_8335 : valid_0_112; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9367 = 3'h5 == state ? _GEN_8336 : valid_0_113; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9368 = 3'h5 == state ? _GEN_8337 : valid_0_114; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9369 = 3'h5 == state ? _GEN_8338 : valid_0_115; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9370 = 3'h5 == state ? _GEN_8339 : valid_0_116; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9371 = 3'h5 == state ? _GEN_8340 : valid_0_117; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9372 = 3'h5 == state ? _GEN_8341 : valid_0_118; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9373 = 3'h5 == state ? _GEN_8342 : valid_0_119; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9374 = 3'h5 == state ? _GEN_8343 : valid_0_120; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9375 = 3'h5 == state ? _GEN_8344 : valid_0_121; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9376 = 3'h5 == state ? _GEN_8345 : valid_0_122; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9377 = 3'h5 == state ? _GEN_8346 : valid_0_123; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9378 = 3'h5 == state ? _GEN_8347 : valid_0_124; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9379 = 3'h5 == state ? _GEN_8348 : valid_0_125; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9380 = 3'h5 == state ? _GEN_8349 : valid_0_126; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9381 = 3'h5 == state ? _GEN_8350 : valid_0_127; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_9382 = 3'h5 == state ? _GEN_8351 : quene; // @[d_cache.scala 64:18 35:24]
  wire [63:0] _GEN_9383 = 3'h5 == state ? _GEN_8352 : ram_1_0; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9384 = 3'h5 == state ? _GEN_8353 : ram_1_1; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9385 = 3'h5 == state ? _GEN_8354 : ram_1_2; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9386 = 3'h5 == state ? _GEN_8355 : ram_1_3; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9387 = 3'h5 == state ? _GEN_8356 : ram_1_4; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9388 = 3'h5 == state ? _GEN_8357 : ram_1_5; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9389 = 3'h5 == state ? _GEN_8358 : ram_1_6; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9390 = 3'h5 == state ? _GEN_8359 : ram_1_7; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9391 = 3'h5 == state ? _GEN_8360 : ram_1_8; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9392 = 3'h5 == state ? _GEN_8361 : ram_1_9; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9393 = 3'h5 == state ? _GEN_8362 : ram_1_10; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9394 = 3'h5 == state ? _GEN_8363 : ram_1_11; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9395 = 3'h5 == state ? _GEN_8364 : ram_1_12; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9396 = 3'h5 == state ? _GEN_8365 : ram_1_13; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9397 = 3'h5 == state ? _GEN_8366 : ram_1_14; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9398 = 3'h5 == state ? _GEN_8367 : ram_1_15; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9399 = 3'h5 == state ? _GEN_8368 : ram_1_16; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9400 = 3'h5 == state ? _GEN_8369 : ram_1_17; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9401 = 3'h5 == state ? _GEN_8370 : ram_1_18; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9402 = 3'h5 == state ? _GEN_8371 : ram_1_19; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9403 = 3'h5 == state ? _GEN_8372 : ram_1_20; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9404 = 3'h5 == state ? _GEN_8373 : ram_1_21; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9405 = 3'h5 == state ? _GEN_8374 : ram_1_22; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9406 = 3'h5 == state ? _GEN_8375 : ram_1_23; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9407 = 3'h5 == state ? _GEN_8376 : ram_1_24; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9408 = 3'h5 == state ? _GEN_8377 : ram_1_25; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9409 = 3'h5 == state ? _GEN_8378 : ram_1_26; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9410 = 3'h5 == state ? _GEN_8379 : ram_1_27; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9411 = 3'h5 == state ? _GEN_8380 : ram_1_28; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9412 = 3'h5 == state ? _GEN_8381 : ram_1_29; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9413 = 3'h5 == state ? _GEN_8382 : ram_1_30; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9414 = 3'h5 == state ? _GEN_8383 : ram_1_31; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9415 = 3'h5 == state ? _GEN_8384 : ram_1_32; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9416 = 3'h5 == state ? _GEN_8385 : ram_1_33; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9417 = 3'h5 == state ? _GEN_8386 : ram_1_34; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9418 = 3'h5 == state ? _GEN_8387 : ram_1_35; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9419 = 3'h5 == state ? _GEN_8388 : ram_1_36; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9420 = 3'h5 == state ? _GEN_8389 : ram_1_37; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9421 = 3'h5 == state ? _GEN_8390 : ram_1_38; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9422 = 3'h5 == state ? _GEN_8391 : ram_1_39; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9423 = 3'h5 == state ? _GEN_8392 : ram_1_40; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9424 = 3'h5 == state ? _GEN_8393 : ram_1_41; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9425 = 3'h5 == state ? _GEN_8394 : ram_1_42; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9426 = 3'h5 == state ? _GEN_8395 : ram_1_43; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9427 = 3'h5 == state ? _GEN_8396 : ram_1_44; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9428 = 3'h5 == state ? _GEN_8397 : ram_1_45; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9429 = 3'h5 == state ? _GEN_8398 : ram_1_46; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9430 = 3'h5 == state ? _GEN_8399 : ram_1_47; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9431 = 3'h5 == state ? _GEN_8400 : ram_1_48; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9432 = 3'h5 == state ? _GEN_8401 : ram_1_49; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9433 = 3'h5 == state ? _GEN_8402 : ram_1_50; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9434 = 3'h5 == state ? _GEN_8403 : ram_1_51; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9435 = 3'h5 == state ? _GEN_8404 : ram_1_52; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9436 = 3'h5 == state ? _GEN_8405 : ram_1_53; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9437 = 3'h5 == state ? _GEN_8406 : ram_1_54; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9438 = 3'h5 == state ? _GEN_8407 : ram_1_55; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9439 = 3'h5 == state ? _GEN_8408 : ram_1_56; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9440 = 3'h5 == state ? _GEN_8409 : ram_1_57; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9441 = 3'h5 == state ? _GEN_8410 : ram_1_58; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9442 = 3'h5 == state ? _GEN_8411 : ram_1_59; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9443 = 3'h5 == state ? _GEN_8412 : ram_1_60; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9444 = 3'h5 == state ? _GEN_8413 : ram_1_61; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9445 = 3'h5 == state ? _GEN_8414 : ram_1_62; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9446 = 3'h5 == state ? _GEN_8415 : ram_1_63; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9447 = 3'h5 == state ? _GEN_8416 : ram_1_64; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9448 = 3'h5 == state ? _GEN_8417 : ram_1_65; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9449 = 3'h5 == state ? _GEN_8418 : ram_1_66; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9450 = 3'h5 == state ? _GEN_8419 : ram_1_67; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9451 = 3'h5 == state ? _GEN_8420 : ram_1_68; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9452 = 3'h5 == state ? _GEN_8421 : ram_1_69; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9453 = 3'h5 == state ? _GEN_8422 : ram_1_70; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9454 = 3'h5 == state ? _GEN_8423 : ram_1_71; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9455 = 3'h5 == state ? _GEN_8424 : ram_1_72; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9456 = 3'h5 == state ? _GEN_8425 : ram_1_73; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9457 = 3'h5 == state ? _GEN_8426 : ram_1_74; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9458 = 3'h5 == state ? _GEN_8427 : ram_1_75; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9459 = 3'h5 == state ? _GEN_8428 : ram_1_76; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9460 = 3'h5 == state ? _GEN_8429 : ram_1_77; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9461 = 3'h5 == state ? _GEN_8430 : ram_1_78; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9462 = 3'h5 == state ? _GEN_8431 : ram_1_79; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9463 = 3'h5 == state ? _GEN_8432 : ram_1_80; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9464 = 3'h5 == state ? _GEN_8433 : ram_1_81; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9465 = 3'h5 == state ? _GEN_8434 : ram_1_82; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9466 = 3'h5 == state ? _GEN_8435 : ram_1_83; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9467 = 3'h5 == state ? _GEN_8436 : ram_1_84; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9468 = 3'h5 == state ? _GEN_8437 : ram_1_85; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9469 = 3'h5 == state ? _GEN_8438 : ram_1_86; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9470 = 3'h5 == state ? _GEN_8439 : ram_1_87; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9471 = 3'h5 == state ? _GEN_8440 : ram_1_88; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9472 = 3'h5 == state ? _GEN_8441 : ram_1_89; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9473 = 3'h5 == state ? _GEN_8442 : ram_1_90; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9474 = 3'h5 == state ? _GEN_8443 : ram_1_91; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9475 = 3'h5 == state ? _GEN_8444 : ram_1_92; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9476 = 3'h5 == state ? _GEN_8445 : ram_1_93; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9477 = 3'h5 == state ? _GEN_8446 : ram_1_94; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9478 = 3'h5 == state ? _GEN_8447 : ram_1_95; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9479 = 3'h5 == state ? _GEN_8448 : ram_1_96; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9480 = 3'h5 == state ? _GEN_8449 : ram_1_97; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9481 = 3'h5 == state ? _GEN_8450 : ram_1_98; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9482 = 3'h5 == state ? _GEN_8451 : ram_1_99; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9483 = 3'h5 == state ? _GEN_8452 : ram_1_100; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9484 = 3'h5 == state ? _GEN_8453 : ram_1_101; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9485 = 3'h5 == state ? _GEN_8454 : ram_1_102; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9486 = 3'h5 == state ? _GEN_8455 : ram_1_103; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9487 = 3'h5 == state ? _GEN_8456 : ram_1_104; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9488 = 3'h5 == state ? _GEN_8457 : ram_1_105; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9489 = 3'h5 == state ? _GEN_8458 : ram_1_106; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9490 = 3'h5 == state ? _GEN_8459 : ram_1_107; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9491 = 3'h5 == state ? _GEN_8460 : ram_1_108; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9492 = 3'h5 == state ? _GEN_8461 : ram_1_109; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9493 = 3'h5 == state ? _GEN_8462 : ram_1_110; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9494 = 3'h5 == state ? _GEN_8463 : ram_1_111; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9495 = 3'h5 == state ? _GEN_8464 : ram_1_112; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9496 = 3'h5 == state ? _GEN_8465 : ram_1_113; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9497 = 3'h5 == state ? _GEN_8466 : ram_1_114; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9498 = 3'h5 == state ? _GEN_8467 : ram_1_115; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9499 = 3'h5 == state ? _GEN_8468 : ram_1_116; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9500 = 3'h5 == state ? _GEN_8469 : ram_1_117; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9501 = 3'h5 == state ? _GEN_8470 : ram_1_118; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9502 = 3'h5 == state ? _GEN_8471 : ram_1_119; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9503 = 3'h5 == state ? _GEN_8472 : ram_1_120; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9504 = 3'h5 == state ? _GEN_8473 : ram_1_121; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9505 = 3'h5 == state ? _GEN_8474 : ram_1_122; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9506 = 3'h5 == state ? _GEN_8475 : ram_1_123; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9507 = 3'h5 == state ? _GEN_8476 : ram_1_124; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9508 = 3'h5 == state ? _GEN_8477 : ram_1_125; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9509 = 3'h5 == state ? _GEN_8478 : ram_1_126; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_9510 = 3'h5 == state ? _GEN_8479 : ram_1_127; // @[d_cache.scala 64:18 19:24]
  wire [31:0] _GEN_9511 = 3'h5 == state ? _GEN_8480 : tag_1_0; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9512 = 3'h5 == state ? _GEN_8481 : tag_1_1; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9513 = 3'h5 == state ? _GEN_8482 : tag_1_2; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9514 = 3'h5 == state ? _GEN_8483 : tag_1_3; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9515 = 3'h5 == state ? _GEN_8484 : tag_1_4; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9516 = 3'h5 == state ? _GEN_8485 : tag_1_5; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9517 = 3'h5 == state ? _GEN_8486 : tag_1_6; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9518 = 3'h5 == state ? _GEN_8487 : tag_1_7; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9519 = 3'h5 == state ? _GEN_8488 : tag_1_8; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9520 = 3'h5 == state ? _GEN_8489 : tag_1_9; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9521 = 3'h5 == state ? _GEN_8490 : tag_1_10; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9522 = 3'h5 == state ? _GEN_8491 : tag_1_11; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9523 = 3'h5 == state ? _GEN_8492 : tag_1_12; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9524 = 3'h5 == state ? _GEN_8493 : tag_1_13; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9525 = 3'h5 == state ? _GEN_8494 : tag_1_14; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9526 = 3'h5 == state ? _GEN_8495 : tag_1_15; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9527 = 3'h5 == state ? _GEN_8496 : tag_1_16; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9528 = 3'h5 == state ? _GEN_8497 : tag_1_17; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9529 = 3'h5 == state ? _GEN_8498 : tag_1_18; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9530 = 3'h5 == state ? _GEN_8499 : tag_1_19; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9531 = 3'h5 == state ? _GEN_8500 : tag_1_20; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9532 = 3'h5 == state ? _GEN_8501 : tag_1_21; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9533 = 3'h5 == state ? _GEN_8502 : tag_1_22; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9534 = 3'h5 == state ? _GEN_8503 : tag_1_23; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9535 = 3'h5 == state ? _GEN_8504 : tag_1_24; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9536 = 3'h5 == state ? _GEN_8505 : tag_1_25; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9537 = 3'h5 == state ? _GEN_8506 : tag_1_26; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9538 = 3'h5 == state ? _GEN_8507 : tag_1_27; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9539 = 3'h5 == state ? _GEN_8508 : tag_1_28; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9540 = 3'h5 == state ? _GEN_8509 : tag_1_29; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9541 = 3'h5 == state ? _GEN_8510 : tag_1_30; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9542 = 3'h5 == state ? _GEN_8511 : tag_1_31; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9543 = 3'h5 == state ? _GEN_8512 : tag_1_32; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9544 = 3'h5 == state ? _GEN_8513 : tag_1_33; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9545 = 3'h5 == state ? _GEN_8514 : tag_1_34; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9546 = 3'h5 == state ? _GEN_8515 : tag_1_35; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9547 = 3'h5 == state ? _GEN_8516 : tag_1_36; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9548 = 3'h5 == state ? _GEN_8517 : tag_1_37; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9549 = 3'h5 == state ? _GEN_8518 : tag_1_38; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9550 = 3'h5 == state ? _GEN_8519 : tag_1_39; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9551 = 3'h5 == state ? _GEN_8520 : tag_1_40; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9552 = 3'h5 == state ? _GEN_8521 : tag_1_41; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9553 = 3'h5 == state ? _GEN_8522 : tag_1_42; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9554 = 3'h5 == state ? _GEN_8523 : tag_1_43; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9555 = 3'h5 == state ? _GEN_8524 : tag_1_44; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9556 = 3'h5 == state ? _GEN_8525 : tag_1_45; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9557 = 3'h5 == state ? _GEN_8526 : tag_1_46; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9558 = 3'h5 == state ? _GEN_8527 : tag_1_47; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9559 = 3'h5 == state ? _GEN_8528 : tag_1_48; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9560 = 3'h5 == state ? _GEN_8529 : tag_1_49; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9561 = 3'h5 == state ? _GEN_8530 : tag_1_50; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9562 = 3'h5 == state ? _GEN_8531 : tag_1_51; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9563 = 3'h5 == state ? _GEN_8532 : tag_1_52; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9564 = 3'h5 == state ? _GEN_8533 : tag_1_53; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9565 = 3'h5 == state ? _GEN_8534 : tag_1_54; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9566 = 3'h5 == state ? _GEN_8535 : tag_1_55; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9567 = 3'h5 == state ? _GEN_8536 : tag_1_56; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9568 = 3'h5 == state ? _GEN_8537 : tag_1_57; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9569 = 3'h5 == state ? _GEN_8538 : tag_1_58; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9570 = 3'h5 == state ? _GEN_8539 : tag_1_59; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9571 = 3'h5 == state ? _GEN_8540 : tag_1_60; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9572 = 3'h5 == state ? _GEN_8541 : tag_1_61; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9573 = 3'h5 == state ? _GEN_8542 : tag_1_62; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9574 = 3'h5 == state ? _GEN_8543 : tag_1_63; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9575 = 3'h5 == state ? _GEN_8544 : tag_1_64; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9576 = 3'h5 == state ? _GEN_8545 : tag_1_65; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9577 = 3'h5 == state ? _GEN_8546 : tag_1_66; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9578 = 3'h5 == state ? _GEN_8547 : tag_1_67; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9579 = 3'h5 == state ? _GEN_8548 : tag_1_68; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9580 = 3'h5 == state ? _GEN_8549 : tag_1_69; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9581 = 3'h5 == state ? _GEN_8550 : tag_1_70; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9582 = 3'h5 == state ? _GEN_8551 : tag_1_71; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9583 = 3'h5 == state ? _GEN_8552 : tag_1_72; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9584 = 3'h5 == state ? _GEN_8553 : tag_1_73; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9585 = 3'h5 == state ? _GEN_8554 : tag_1_74; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9586 = 3'h5 == state ? _GEN_8555 : tag_1_75; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9587 = 3'h5 == state ? _GEN_8556 : tag_1_76; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9588 = 3'h5 == state ? _GEN_8557 : tag_1_77; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9589 = 3'h5 == state ? _GEN_8558 : tag_1_78; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9590 = 3'h5 == state ? _GEN_8559 : tag_1_79; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9591 = 3'h5 == state ? _GEN_8560 : tag_1_80; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9592 = 3'h5 == state ? _GEN_8561 : tag_1_81; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9593 = 3'h5 == state ? _GEN_8562 : tag_1_82; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9594 = 3'h5 == state ? _GEN_8563 : tag_1_83; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9595 = 3'h5 == state ? _GEN_8564 : tag_1_84; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9596 = 3'h5 == state ? _GEN_8565 : tag_1_85; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9597 = 3'h5 == state ? _GEN_8566 : tag_1_86; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9598 = 3'h5 == state ? _GEN_8567 : tag_1_87; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9599 = 3'h5 == state ? _GEN_8568 : tag_1_88; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9600 = 3'h5 == state ? _GEN_8569 : tag_1_89; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9601 = 3'h5 == state ? _GEN_8570 : tag_1_90; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9602 = 3'h5 == state ? _GEN_8571 : tag_1_91; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9603 = 3'h5 == state ? _GEN_8572 : tag_1_92; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9604 = 3'h5 == state ? _GEN_8573 : tag_1_93; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9605 = 3'h5 == state ? _GEN_8574 : tag_1_94; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9606 = 3'h5 == state ? _GEN_8575 : tag_1_95; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9607 = 3'h5 == state ? _GEN_8576 : tag_1_96; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9608 = 3'h5 == state ? _GEN_8577 : tag_1_97; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9609 = 3'h5 == state ? _GEN_8578 : tag_1_98; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9610 = 3'h5 == state ? _GEN_8579 : tag_1_99; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9611 = 3'h5 == state ? _GEN_8580 : tag_1_100; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9612 = 3'h5 == state ? _GEN_8581 : tag_1_101; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9613 = 3'h5 == state ? _GEN_8582 : tag_1_102; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9614 = 3'h5 == state ? _GEN_8583 : tag_1_103; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9615 = 3'h5 == state ? _GEN_8584 : tag_1_104; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9616 = 3'h5 == state ? _GEN_8585 : tag_1_105; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9617 = 3'h5 == state ? _GEN_8586 : tag_1_106; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9618 = 3'h5 == state ? _GEN_8587 : tag_1_107; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9619 = 3'h5 == state ? _GEN_8588 : tag_1_108; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9620 = 3'h5 == state ? _GEN_8589 : tag_1_109; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9621 = 3'h5 == state ? _GEN_8590 : tag_1_110; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9622 = 3'h5 == state ? _GEN_8591 : tag_1_111; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9623 = 3'h5 == state ? _GEN_8592 : tag_1_112; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9624 = 3'h5 == state ? _GEN_8593 : tag_1_113; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9625 = 3'h5 == state ? _GEN_8594 : tag_1_114; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9626 = 3'h5 == state ? _GEN_8595 : tag_1_115; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9627 = 3'h5 == state ? _GEN_8596 : tag_1_116; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9628 = 3'h5 == state ? _GEN_8597 : tag_1_117; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9629 = 3'h5 == state ? _GEN_8598 : tag_1_118; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9630 = 3'h5 == state ? _GEN_8599 : tag_1_119; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9631 = 3'h5 == state ? _GEN_8600 : tag_1_120; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9632 = 3'h5 == state ? _GEN_8601 : tag_1_121; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9633 = 3'h5 == state ? _GEN_8602 : tag_1_122; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9634 = 3'h5 == state ? _GEN_8603 : tag_1_123; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9635 = 3'h5 == state ? _GEN_8604 : tag_1_124; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9636 = 3'h5 == state ? _GEN_8605 : tag_1_125; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9637 = 3'h5 == state ? _GEN_8606 : tag_1_126; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_9638 = 3'h5 == state ? _GEN_8607 : tag_1_127; // @[d_cache.scala 64:18 21:24]
  wire  _GEN_9639 = 3'h5 == state ? _GEN_8608 : valid_1_0; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9640 = 3'h5 == state ? _GEN_8609 : valid_1_1; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9641 = 3'h5 == state ? _GEN_8610 : valid_1_2; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9642 = 3'h5 == state ? _GEN_8611 : valid_1_3; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9643 = 3'h5 == state ? _GEN_8612 : valid_1_4; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9644 = 3'h5 == state ? _GEN_8613 : valid_1_5; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9645 = 3'h5 == state ? _GEN_8614 : valid_1_6; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9646 = 3'h5 == state ? _GEN_8615 : valid_1_7; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9647 = 3'h5 == state ? _GEN_8616 : valid_1_8; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9648 = 3'h5 == state ? _GEN_8617 : valid_1_9; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9649 = 3'h5 == state ? _GEN_8618 : valid_1_10; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9650 = 3'h5 == state ? _GEN_8619 : valid_1_11; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9651 = 3'h5 == state ? _GEN_8620 : valid_1_12; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9652 = 3'h5 == state ? _GEN_8621 : valid_1_13; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9653 = 3'h5 == state ? _GEN_8622 : valid_1_14; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9654 = 3'h5 == state ? _GEN_8623 : valid_1_15; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9655 = 3'h5 == state ? _GEN_8624 : valid_1_16; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9656 = 3'h5 == state ? _GEN_8625 : valid_1_17; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9657 = 3'h5 == state ? _GEN_8626 : valid_1_18; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9658 = 3'h5 == state ? _GEN_8627 : valid_1_19; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9659 = 3'h5 == state ? _GEN_8628 : valid_1_20; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9660 = 3'h5 == state ? _GEN_8629 : valid_1_21; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9661 = 3'h5 == state ? _GEN_8630 : valid_1_22; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9662 = 3'h5 == state ? _GEN_8631 : valid_1_23; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9663 = 3'h5 == state ? _GEN_8632 : valid_1_24; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9664 = 3'h5 == state ? _GEN_8633 : valid_1_25; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9665 = 3'h5 == state ? _GEN_8634 : valid_1_26; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9666 = 3'h5 == state ? _GEN_8635 : valid_1_27; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9667 = 3'h5 == state ? _GEN_8636 : valid_1_28; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9668 = 3'h5 == state ? _GEN_8637 : valid_1_29; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9669 = 3'h5 == state ? _GEN_8638 : valid_1_30; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9670 = 3'h5 == state ? _GEN_8639 : valid_1_31; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9671 = 3'h5 == state ? _GEN_8640 : valid_1_32; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9672 = 3'h5 == state ? _GEN_8641 : valid_1_33; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9673 = 3'h5 == state ? _GEN_8642 : valid_1_34; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9674 = 3'h5 == state ? _GEN_8643 : valid_1_35; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9675 = 3'h5 == state ? _GEN_8644 : valid_1_36; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9676 = 3'h5 == state ? _GEN_8645 : valid_1_37; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9677 = 3'h5 == state ? _GEN_8646 : valid_1_38; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9678 = 3'h5 == state ? _GEN_8647 : valid_1_39; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9679 = 3'h5 == state ? _GEN_8648 : valid_1_40; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9680 = 3'h5 == state ? _GEN_8649 : valid_1_41; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9681 = 3'h5 == state ? _GEN_8650 : valid_1_42; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9682 = 3'h5 == state ? _GEN_8651 : valid_1_43; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9683 = 3'h5 == state ? _GEN_8652 : valid_1_44; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9684 = 3'h5 == state ? _GEN_8653 : valid_1_45; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9685 = 3'h5 == state ? _GEN_8654 : valid_1_46; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9686 = 3'h5 == state ? _GEN_8655 : valid_1_47; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9687 = 3'h5 == state ? _GEN_8656 : valid_1_48; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9688 = 3'h5 == state ? _GEN_8657 : valid_1_49; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9689 = 3'h5 == state ? _GEN_8658 : valid_1_50; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9690 = 3'h5 == state ? _GEN_8659 : valid_1_51; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9691 = 3'h5 == state ? _GEN_8660 : valid_1_52; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9692 = 3'h5 == state ? _GEN_8661 : valid_1_53; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9693 = 3'h5 == state ? _GEN_8662 : valid_1_54; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9694 = 3'h5 == state ? _GEN_8663 : valid_1_55; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9695 = 3'h5 == state ? _GEN_8664 : valid_1_56; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9696 = 3'h5 == state ? _GEN_8665 : valid_1_57; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9697 = 3'h5 == state ? _GEN_8666 : valid_1_58; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9698 = 3'h5 == state ? _GEN_8667 : valid_1_59; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9699 = 3'h5 == state ? _GEN_8668 : valid_1_60; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9700 = 3'h5 == state ? _GEN_8669 : valid_1_61; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9701 = 3'h5 == state ? _GEN_8670 : valid_1_62; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9702 = 3'h5 == state ? _GEN_8671 : valid_1_63; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9703 = 3'h5 == state ? _GEN_8672 : valid_1_64; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9704 = 3'h5 == state ? _GEN_8673 : valid_1_65; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9705 = 3'h5 == state ? _GEN_8674 : valid_1_66; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9706 = 3'h5 == state ? _GEN_8675 : valid_1_67; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9707 = 3'h5 == state ? _GEN_8676 : valid_1_68; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9708 = 3'h5 == state ? _GEN_8677 : valid_1_69; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9709 = 3'h5 == state ? _GEN_8678 : valid_1_70; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9710 = 3'h5 == state ? _GEN_8679 : valid_1_71; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9711 = 3'h5 == state ? _GEN_8680 : valid_1_72; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9712 = 3'h5 == state ? _GEN_8681 : valid_1_73; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9713 = 3'h5 == state ? _GEN_8682 : valid_1_74; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9714 = 3'h5 == state ? _GEN_8683 : valid_1_75; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9715 = 3'h5 == state ? _GEN_8684 : valid_1_76; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9716 = 3'h5 == state ? _GEN_8685 : valid_1_77; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9717 = 3'h5 == state ? _GEN_8686 : valid_1_78; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9718 = 3'h5 == state ? _GEN_8687 : valid_1_79; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9719 = 3'h5 == state ? _GEN_8688 : valid_1_80; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9720 = 3'h5 == state ? _GEN_8689 : valid_1_81; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9721 = 3'h5 == state ? _GEN_8690 : valid_1_82; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9722 = 3'h5 == state ? _GEN_8691 : valid_1_83; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9723 = 3'h5 == state ? _GEN_8692 : valid_1_84; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9724 = 3'h5 == state ? _GEN_8693 : valid_1_85; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9725 = 3'h5 == state ? _GEN_8694 : valid_1_86; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9726 = 3'h5 == state ? _GEN_8695 : valid_1_87; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9727 = 3'h5 == state ? _GEN_8696 : valid_1_88; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9728 = 3'h5 == state ? _GEN_8697 : valid_1_89; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9729 = 3'h5 == state ? _GEN_8698 : valid_1_90; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9730 = 3'h5 == state ? _GEN_8699 : valid_1_91; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9731 = 3'h5 == state ? _GEN_8700 : valid_1_92; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9732 = 3'h5 == state ? _GEN_8701 : valid_1_93; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9733 = 3'h5 == state ? _GEN_8702 : valid_1_94; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9734 = 3'h5 == state ? _GEN_8703 : valid_1_95; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9735 = 3'h5 == state ? _GEN_8704 : valid_1_96; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9736 = 3'h5 == state ? _GEN_8705 : valid_1_97; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9737 = 3'h5 == state ? _GEN_8706 : valid_1_98; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9738 = 3'h5 == state ? _GEN_8707 : valid_1_99; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9739 = 3'h5 == state ? _GEN_8708 : valid_1_100; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9740 = 3'h5 == state ? _GEN_8709 : valid_1_101; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9741 = 3'h5 == state ? _GEN_8710 : valid_1_102; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9742 = 3'h5 == state ? _GEN_8711 : valid_1_103; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9743 = 3'h5 == state ? _GEN_8712 : valid_1_104; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9744 = 3'h5 == state ? _GEN_8713 : valid_1_105; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9745 = 3'h5 == state ? _GEN_8714 : valid_1_106; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9746 = 3'h5 == state ? _GEN_8715 : valid_1_107; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9747 = 3'h5 == state ? _GEN_8716 : valid_1_108; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9748 = 3'h5 == state ? _GEN_8717 : valid_1_109; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9749 = 3'h5 == state ? _GEN_8718 : valid_1_110; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9750 = 3'h5 == state ? _GEN_8719 : valid_1_111; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9751 = 3'h5 == state ? _GEN_8720 : valid_1_112; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9752 = 3'h5 == state ? _GEN_8721 : valid_1_113; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9753 = 3'h5 == state ? _GEN_8722 : valid_1_114; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9754 = 3'h5 == state ? _GEN_8723 : valid_1_115; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9755 = 3'h5 == state ? _GEN_8724 : valid_1_116; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9756 = 3'h5 == state ? _GEN_8725 : valid_1_117; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9757 = 3'h5 == state ? _GEN_8726 : valid_1_118; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9758 = 3'h5 == state ? _GEN_8727 : valid_1_119; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9759 = 3'h5 == state ? _GEN_8728 : valid_1_120; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9760 = 3'h5 == state ? _GEN_8729 : valid_1_121; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9761 = 3'h5 == state ? _GEN_8730 : valid_1_122; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9762 = 3'h5 == state ? _GEN_8731 : valid_1_123; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9763 = 3'h5 == state ? _GEN_8732 : valid_1_124; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9764 = 3'h5 == state ? _GEN_8733 : valid_1_125; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9765 = 3'h5 == state ? _GEN_8734 : valid_1_126; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_9766 = 3'h5 == state ? _GEN_8735 : valid_1_127; // @[d_cache.scala 64:18 23:26]
  wire [63:0] _GEN_9767 = 3'h5 == state ? _GEN_8736 : write_back_data; // @[d_cache.scala 64:18 29:34]
  wire [38:0] _GEN_9768 = 3'h5 == state ? _GEN_8737 : {{7'd0}, write_back_addr}; // @[d_cache.scala 64:18 30:34]
  wire  _GEN_9769 = 3'h5 == state ? _GEN_8738 : dirty_0_0; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9770 = 3'h5 == state ? _GEN_8739 : dirty_0_1; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9771 = 3'h5 == state ? _GEN_8740 : dirty_0_2; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9772 = 3'h5 == state ? _GEN_8741 : dirty_0_3; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9773 = 3'h5 == state ? _GEN_8742 : dirty_0_4; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9774 = 3'h5 == state ? _GEN_8743 : dirty_0_5; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9775 = 3'h5 == state ? _GEN_8744 : dirty_0_6; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9776 = 3'h5 == state ? _GEN_8745 : dirty_0_7; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9777 = 3'h5 == state ? _GEN_8746 : dirty_0_8; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9778 = 3'h5 == state ? _GEN_8747 : dirty_0_9; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9779 = 3'h5 == state ? _GEN_8748 : dirty_0_10; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9780 = 3'h5 == state ? _GEN_8749 : dirty_0_11; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9781 = 3'h5 == state ? _GEN_8750 : dirty_0_12; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9782 = 3'h5 == state ? _GEN_8751 : dirty_0_13; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9783 = 3'h5 == state ? _GEN_8752 : dirty_0_14; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9784 = 3'h5 == state ? _GEN_8753 : dirty_0_15; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9785 = 3'h5 == state ? _GEN_8754 : dirty_0_16; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9786 = 3'h5 == state ? _GEN_8755 : dirty_0_17; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9787 = 3'h5 == state ? _GEN_8756 : dirty_0_18; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9788 = 3'h5 == state ? _GEN_8757 : dirty_0_19; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9789 = 3'h5 == state ? _GEN_8758 : dirty_0_20; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9790 = 3'h5 == state ? _GEN_8759 : dirty_0_21; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9791 = 3'h5 == state ? _GEN_8760 : dirty_0_22; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9792 = 3'h5 == state ? _GEN_8761 : dirty_0_23; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9793 = 3'h5 == state ? _GEN_8762 : dirty_0_24; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9794 = 3'h5 == state ? _GEN_8763 : dirty_0_25; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9795 = 3'h5 == state ? _GEN_8764 : dirty_0_26; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9796 = 3'h5 == state ? _GEN_8765 : dirty_0_27; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9797 = 3'h5 == state ? _GEN_8766 : dirty_0_28; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9798 = 3'h5 == state ? _GEN_8767 : dirty_0_29; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9799 = 3'h5 == state ? _GEN_8768 : dirty_0_30; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9800 = 3'h5 == state ? _GEN_8769 : dirty_0_31; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9801 = 3'h5 == state ? _GEN_8770 : dirty_0_32; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9802 = 3'h5 == state ? _GEN_8771 : dirty_0_33; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9803 = 3'h5 == state ? _GEN_8772 : dirty_0_34; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9804 = 3'h5 == state ? _GEN_8773 : dirty_0_35; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9805 = 3'h5 == state ? _GEN_8774 : dirty_0_36; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9806 = 3'h5 == state ? _GEN_8775 : dirty_0_37; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9807 = 3'h5 == state ? _GEN_8776 : dirty_0_38; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9808 = 3'h5 == state ? _GEN_8777 : dirty_0_39; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9809 = 3'h5 == state ? _GEN_8778 : dirty_0_40; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9810 = 3'h5 == state ? _GEN_8779 : dirty_0_41; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9811 = 3'h5 == state ? _GEN_8780 : dirty_0_42; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9812 = 3'h5 == state ? _GEN_8781 : dirty_0_43; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9813 = 3'h5 == state ? _GEN_8782 : dirty_0_44; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9814 = 3'h5 == state ? _GEN_8783 : dirty_0_45; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9815 = 3'h5 == state ? _GEN_8784 : dirty_0_46; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9816 = 3'h5 == state ? _GEN_8785 : dirty_0_47; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9817 = 3'h5 == state ? _GEN_8786 : dirty_0_48; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9818 = 3'h5 == state ? _GEN_8787 : dirty_0_49; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9819 = 3'h5 == state ? _GEN_8788 : dirty_0_50; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9820 = 3'h5 == state ? _GEN_8789 : dirty_0_51; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9821 = 3'h5 == state ? _GEN_8790 : dirty_0_52; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9822 = 3'h5 == state ? _GEN_8791 : dirty_0_53; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9823 = 3'h5 == state ? _GEN_8792 : dirty_0_54; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9824 = 3'h5 == state ? _GEN_8793 : dirty_0_55; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9825 = 3'h5 == state ? _GEN_8794 : dirty_0_56; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9826 = 3'h5 == state ? _GEN_8795 : dirty_0_57; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9827 = 3'h5 == state ? _GEN_8796 : dirty_0_58; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9828 = 3'h5 == state ? _GEN_8797 : dirty_0_59; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9829 = 3'h5 == state ? _GEN_8798 : dirty_0_60; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9830 = 3'h5 == state ? _GEN_8799 : dirty_0_61; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9831 = 3'h5 == state ? _GEN_8800 : dirty_0_62; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9832 = 3'h5 == state ? _GEN_8801 : dirty_0_63; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9833 = 3'h5 == state ? _GEN_8802 : dirty_0_64; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9834 = 3'h5 == state ? _GEN_8803 : dirty_0_65; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9835 = 3'h5 == state ? _GEN_8804 : dirty_0_66; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9836 = 3'h5 == state ? _GEN_8805 : dirty_0_67; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9837 = 3'h5 == state ? _GEN_8806 : dirty_0_68; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9838 = 3'h5 == state ? _GEN_8807 : dirty_0_69; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9839 = 3'h5 == state ? _GEN_8808 : dirty_0_70; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9840 = 3'h5 == state ? _GEN_8809 : dirty_0_71; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9841 = 3'h5 == state ? _GEN_8810 : dirty_0_72; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9842 = 3'h5 == state ? _GEN_8811 : dirty_0_73; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9843 = 3'h5 == state ? _GEN_8812 : dirty_0_74; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9844 = 3'h5 == state ? _GEN_8813 : dirty_0_75; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9845 = 3'h5 == state ? _GEN_8814 : dirty_0_76; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9846 = 3'h5 == state ? _GEN_8815 : dirty_0_77; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9847 = 3'h5 == state ? _GEN_8816 : dirty_0_78; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9848 = 3'h5 == state ? _GEN_8817 : dirty_0_79; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9849 = 3'h5 == state ? _GEN_8818 : dirty_0_80; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9850 = 3'h5 == state ? _GEN_8819 : dirty_0_81; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9851 = 3'h5 == state ? _GEN_8820 : dirty_0_82; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9852 = 3'h5 == state ? _GEN_8821 : dirty_0_83; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9853 = 3'h5 == state ? _GEN_8822 : dirty_0_84; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9854 = 3'h5 == state ? _GEN_8823 : dirty_0_85; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9855 = 3'h5 == state ? _GEN_8824 : dirty_0_86; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9856 = 3'h5 == state ? _GEN_8825 : dirty_0_87; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9857 = 3'h5 == state ? _GEN_8826 : dirty_0_88; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9858 = 3'h5 == state ? _GEN_8827 : dirty_0_89; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9859 = 3'h5 == state ? _GEN_8828 : dirty_0_90; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9860 = 3'h5 == state ? _GEN_8829 : dirty_0_91; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9861 = 3'h5 == state ? _GEN_8830 : dirty_0_92; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9862 = 3'h5 == state ? _GEN_8831 : dirty_0_93; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9863 = 3'h5 == state ? _GEN_8832 : dirty_0_94; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9864 = 3'h5 == state ? _GEN_8833 : dirty_0_95; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9865 = 3'h5 == state ? _GEN_8834 : dirty_0_96; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9866 = 3'h5 == state ? _GEN_8835 : dirty_0_97; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9867 = 3'h5 == state ? _GEN_8836 : dirty_0_98; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9868 = 3'h5 == state ? _GEN_8837 : dirty_0_99; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9869 = 3'h5 == state ? _GEN_8838 : dirty_0_100; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9870 = 3'h5 == state ? _GEN_8839 : dirty_0_101; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9871 = 3'h5 == state ? _GEN_8840 : dirty_0_102; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9872 = 3'h5 == state ? _GEN_8841 : dirty_0_103; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9873 = 3'h5 == state ? _GEN_8842 : dirty_0_104; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9874 = 3'h5 == state ? _GEN_8843 : dirty_0_105; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9875 = 3'h5 == state ? _GEN_8844 : dirty_0_106; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9876 = 3'h5 == state ? _GEN_8845 : dirty_0_107; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9877 = 3'h5 == state ? _GEN_8846 : dirty_0_108; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9878 = 3'h5 == state ? _GEN_8847 : dirty_0_109; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9879 = 3'h5 == state ? _GEN_8848 : dirty_0_110; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9880 = 3'h5 == state ? _GEN_8849 : dirty_0_111; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9881 = 3'h5 == state ? _GEN_8850 : dirty_0_112; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9882 = 3'h5 == state ? _GEN_8851 : dirty_0_113; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9883 = 3'h5 == state ? _GEN_8852 : dirty_0_114; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9884 = 3'h5 == state ? _GEN_8853 : dirty_0_115; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9885 = 3'h5 == state ? _GEN_8854 : dirty_0_116; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9886 = 3'h5 == state ? _GEN_8855 : dirty_0_117; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9887 = 3'h5 == state ? _GEN_8856 : dirty_0_118; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9888 = 3'h5 == state ? _GEN_8857 : dirty_0_119; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9889 = 3'h5 == state ? _GEN_8858 : dirty_0_120; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9890 = 3'h5 == state ? _GEN_8859 : dirty_0_121; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9891 = 3'h5 == state ? _GEN_8860 : dirty_0_122; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9892 = 3'h5 == state ? _GEN_8861 : dirty_0_123; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9893 = 3'h5 == state ? _GEN_8862 : dirty_0_124; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9894 = 3'h5 == state ? _GEN_8863 : dirty_0_125; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9895 = 3'h5 == state ? _GEN_8864 : dirty_0_126; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9896 = 3'h5 == state ? _GEN_8865 : dirty_0_127; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_9897 = 3'h5 == state ? _GEN_8866 : dirty_1_0; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9898 = 3'h5 == state ? _GEN_8867 : dirty_1_1; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9899 = 3'h5 == state ? _GEN_8868 : dirty_1_2; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9900 = 3'h5 == state ? _GEN_8869 : dirty_1_3; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9901 = 3'h5 == state ? _GEN_8870 : dirty_1_4; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9902 = 3'h5 == state ? _GEN_8871 : dirty_1_5; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9903 = 3'h5 == state ? _GEN_8872 : dirty_1_6; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9904 = 3'h5 == state ? _GEN_8873 : dirty_1_7; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9905 = 3'h5 == state ? _GEN_8874 : dirty_1_8; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9906 = 3'h5 == state ? _GEN_8875 : dirty_1_9; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9907 = 3'h5 == state ? _GEN_8876 : dirty_1_10; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9908 = 3'h5 == state ? _GEN_8877 : dirty_1_11; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9909 = 3'h5 == state ? _GEN_8878 : dirty_1_12; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9910 = 3'h5 == state ? _GEN_8879 : dirty_1_13; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9911 = 3'h5 == state ? _GEN_8880 : dirty_1_14; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9912 = 3'h5 == state ? _GEN_8881 : dirty_1_15; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9913 = 3'h5 == state ? _GEN_8882 : dirty_1_16; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9914 = 3'h5 == state ? _GEN_8883 : dirty_1_17; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9915 = 3'h5 == state ? _GEN_8884 : dirty_1_18; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9916 = 3'h5 == state ? _GEN_8885 : dirty_1_19; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9917 = 3'h5 == state ? _GEN_8886 : dirty_1_20; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9918 = 3'h5 == state ? _GEN_8887 : dirty_1_21; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9919 = 3'h5 == state ? _GEN_8888 : dirty_1_22; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9920 = 3'h5 == state ? _GEN_8889 : dirty_1_23; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9921 = 3'h5 == state ? _GEN_8890 : dirty_1_24; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9922 = 3'h5 == state ? _GEN_8891 : dirty_1_25; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9923 = 3'h5 == state ? _GEN_8892 : dirty_1_26; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9924 = 3'h5 == state ? _GEN_8893 : dirty_1_27; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9925 = 3'h5 == state ? _GEN_8894 : dirty_1_28; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9926 = 3'h5 == state ? _GEN_8895 : dirty_1_29; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9927 = 3'h5 == state ? _GEN_8896 : dirty_1_30; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9928 = 3'h5 == state ? _GEN_8897 : dirty_1_31; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9929 = 3'h5 == state ? _GEN_8898 : dirty_1_32; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9930 = 3'h5 == state ? _GEN_8899 : dirty_1_33; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9931 = 3'h5 == state ? _GEN_8900 : dirty_1_34; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9932 = 3'h5 == state ? _GEN_8901 : dirty_1_35; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9933 = 3'h5 == state ? _GEN_8902 : dirty_1_36; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9934 = 3'h5 == state ? _GEN_8903 : dirty_1_37; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9935 = 3'h5 == state ? _GEN_8904 : dirty_1_38; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9936 = 3'h5 == state ? _GEN_8905 : dirty_1_39; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9937 = 3'h5 == state ? _GEN_8906 : dirty_1_40; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9938 = 3'h5 == state ? _GEN_8907 : dirty_1_41; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9939 = 3'h5 == state ? _GEN_8908 : dirty_1_42; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9940 = 3'h5 == state ? _GEN_8909 : dirty_1_43; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9941 = 3'h5 == state ? _GEN_8910 : dirty_1_44; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9942 = 3'h5 == state ? _GEN_8911 : dirty_1_45; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9943 = 3'h5 == state ? _GEN_8912 : dirty_1_46; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9944 = 3'h5 == state ? _GEN_8913 : dirty_1_47; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9945 = 3'h5 == state ? _GEN_8914 : dirty_1_48; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9946 = 3'h5 == state ? _GEN_8915 : dirty_1_49; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9947 = 3'h5 == state ? _GEN_8916 : dirty_1_50; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9948 = 3'h5 == state ? _GEN_8917 : dirty_1_51; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9949 = 3'h5 == state ? _GEN_8918 : dirty_1_52; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9950 = 3'h5 == state ? _GEN_8919 : dirty_1_53; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9951 = 3'h5 == state ? _GEN_8920 : dirty_1_54; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9952 = 3'h5 == state ? _GEN_8921 : dirty_1_55; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9953 = 3'h5 == state ? _GEN_8922 : dirty_1_56; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9954 = 3'h5 == state ? _GEN_8923 : dirty_1_57; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9955 = 3'h5 == state ? _GEN_8924 : dirty_1_58; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9956 = 3'h5 == state ? _GEN_8925 : dirty_1_59; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9957 = 3'h5 == state ? _GEN_8926 : dirty_1_60; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9958 = 3'h5 == state ? _GEN_8927 : dirty_1_61; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9959 = 3'h5 == state ? _GEN_8928 : dirty_1_62; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9960 = 3'h5 == state ? _GEN_8929 : dirty_1_63; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9961 = 3'h5 == state ? _GEN_8930 : dirty_1_64; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9962 = 3'h5 == state ? _GEN_8931 : dirty_1_65; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9963 = 3'h5 == state ? _GEN_8932 : dirty_1_66; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9964 = 3'h5 == state ? _GEN_8933 : dirty_1_67; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9965 = 3'h5 == state ? _GEN_8934 : dirty_1_68; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9966 = 3'h5 == state ? _GEN_8935 : dirty_1_69; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9967 = 3'h5 == state ? _GEN_8936 : dirty_1_70; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9968 = 3'h5 == state ? _GEN_8937 : dirty_1_71; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9969 = 3'h5 == state ? _GEN_8938 : dirty_1_72; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9970 = 3'h5 == state ? _GEN_8939 : dirty_1_73; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9971 = 3'h5 == state ? _GEN_8940 : dirty_1_74; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9972 = 3'h5 == state ? _GEN_8941 : dirty_1_75; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9973 = 3'h5 == state ? _GEN_8942 : dirty_1_76; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9974 = 3'h5 == state ? _GEN_8943 : dirty_1_77; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9975 = 3'h5 == state ? _GEN_8944 : dirty_1_78; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9976 = 3'h5 == state ? _GEN_8945 : dirty_1_79; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9977 = 3'h5 == state ? _GEN_8946 : dirty_1_80; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9978 = 3'h5 == state ? _GEN_8947 : dirty_1_81; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9979 = 3'h5 == state ? _GEN_8948 : dirty_1_82; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9980 = 3'h5 == state ? _GEN_8949 : dirty_1_83; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9981 = 3'h5 == state ? _GEN_8950 : dirty_1_84; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9982 = 3'h5 == state ? _GEN_8951 : dirty_1_85; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9983 = 3'h5 == state ? _GEN_8952 : dirty_1_86; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9984 = 3'h5 == state ? _GEN_8953 : dirty_1_87; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9985 = 3'h5 == state ? _GEN_8954 : dirty_1_88; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9986 = 3'h5 == state ? _GEN_8955 : dirty_1_89; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9987 = 3'h5 == state ? _GEN_8956 : dirty_1_90; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9988 = 3'h5 == state ? _GEN_8957 : dirty_1_91; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9989 = 3'h5 == state ? _GEN_8958 : dirty_1_92; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9990 = 3'h5 == state ? _GEN_8959 : dirty_1_93; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9991 = 3'h5 == state ? _GEN_8960 : dirty_1_94; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9992 = 3'h5 == state ? _GEN_8961 : dirty_1_95; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9993 = 3'h5 == state ? _GEN_8962 : dirty_1_96; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9994 = 3'h5 == state ? _GEN_8963 : dirty_1_97; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9995 = 3'h5 == state ? _GEN_8964 : dirty_1_98; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9996 = 3'h5 == state ? _GEN_8965 : dirty_1_99; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9997 = 3'h5 == state ? _GEN_8966 : dirty_1_100; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9998 = 3'h5 == state ? _GEN_8967 : dirty_1_101; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_9999 = 3'h5 == state ? _GEN_8968 : dirty_1_102; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10000 = 3'h5 == state ? _GEN_8969 : dirty_1_103; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10001 = 3'h5 == state ? _GEN_8970 : dirty_1_104; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10002 = 3'h5 == state ? _GEN_8971 : dirty_1_105; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10003 = 3'h5 == state ? _GEN_8972 : dirty_1_106; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10004 = 3'h5 == state ? _GEN_8973 : dirty_1_107; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10005 = 3'h5 == state ? _GEN_8974 : dirty_1_108; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10006 = 3'h5 == state ? _GEN_8975 : dirty_1_109; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10007 = 3'h5 == state ? _GEN_8976 : dirty_1_110; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10008 = 3'h5 == state ? _GEN_8977 : dirty_1_111; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10009 = 3'h5 == state ? _GEN_8978 : dirty_1_112; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10010 = 3'h5 == state ? _GEN_8979 : dirty_1_113; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10011 = 3'h5 == state ? _GEN_8980 : dirty_1_114; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10012 = 3'h5 == state ? _GEN_8981 : dirty_1_115; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10013 = 3'h5 == state ? _GEN_8982 : dirty_1_116; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10014 = 3'h5 == state ? _GEN_8983 : dirty_1_117; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10015 = 3'h5 == state ? _GEN_8984 : dirty_1_118; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10016 = 3'h5 == state ? _GEN_8985 : dirty_1_119; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10017 = 3'h5 == state ? _GEN_8986 : dirty_1_120; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10018 = 3'h5 == state ? _GEN_8987 : dirty_1_121; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10019 = 3'h5 == state ? _GEN_8988 : dirty_1_122; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10020 = 3'h5 == state ? _GEN_8989 : dirty_1_123; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10021 = 3'h5 == state ? _GEN_8990 : dirty_1_124; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10022 = 3'h5 == state ? _GEN_8991 : dirty_1_125; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10023 = 3'h5 == state ? _GEN_8992 : dirty_1_126; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10024 = 3'h5 == state ? _GEN_8993 : dirty_1_127; // @[d_cache.scala 64:18 25:26]
  wire [2:0] _GEN_10025 = 3'h4 == state ? _GEN_2061 : _GEN_8997; // @[d_cache.scala 64:18]
  wire [63:0] _GEN_10026 = 3'h4 == state ? ram_0_0 : _GEN_8998; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10027 = 3'h4 == state ? ram_0_1 : _GEN_8999; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10028 = 3'h4 == state ? ram_0_2 : _GEN_9000; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10029 = 3'h4 == state ? ram_0_3 : _GEN_9001; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10030 = 3'h4 == state ? ram_0_4 : _GEN_9002; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10031 = 3'h4 == state ? ram_0_5 : _GEN_9003; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10032 = 3'h4 == state ? ram_0_6 : _GEN_9004; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10033 = 3'h4 == state ? ram_0_7 : _GEN_9005; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10034 = 3'h4 == state ? ram_0_8 : _GEN_9006; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10035 = 3'h4 == state ? ram_0_9 : _GEN_9007; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10036 = 3'h4 == state ? ram_0_10 : _GEN_9008; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10037 = 3'h4 == state ? ram_0_11 : _GEN_9009; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10038 = 3'h4 == state ? ram_0_12 : _GEN_9010; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10039 = 3'h4 == state ? ram_0_13 : _GEN_9011; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10040 = 3'h4 == state ? ram_0_14 : _GEN_9012; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10041 = 3'h4 == state ? ram_0_15 : _GEN_9013; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10042 = 3'h4 == state ? ram_0_16 : _GEN_9014; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10043 = 3'h4 == state ? ram_0_17 : _GEN_9015; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10044 = 3'h4 == state ? ram_0_18 : _GEN_9016; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10045 = 3'h4 == state ? ram_0_19 : _GEN_9017; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10046 = 3'h4 == state ? ram_0_20 : _GEN_9018; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10047 = 3'h4 == state ? ram_0_21 : _GEN_9019; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10048 = 3'h4 == state ? ram_0_22 : _GEN_9020; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10049 = 3'h4 == state ? ram_0_23 : _GEN_9021; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10050 = 3'h4 == state ? ram_0_24 : _GEN_9022; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10051 = 3'h4 == state ? ram_0_25 : _GEN_9023; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10052 = 3'h4 == state ? ram_0_26 : _GEN_9024; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10053 = 3'h4 == state ? ram_0_27 : _GEN_9025; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10054 = 3'h4 == state ? ram_0_28 : _GEN_9026; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10055 = 3'h4 == state ? ram_0_29 : _GEN_9027; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10056 = 3'h4 == state ? ram_0_30 : _GEN_9028; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10057 = 3'h4 == state ? ram_0_31 : _GEN_9029; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10058 = 3'h4 == state ? ram_0_32 : _GEN_9030; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10059 = 3'h4 == state ? ram_0_33 : _GEN_9031; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10060 = 3'h4 == state ? ram_0_34 : _GEN_9032; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10061 = 3'h4 == state ? ram_0_35 : _GEN_9033; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10062 = 3'h4 == state ? ram_0_36 : _GEN_9034; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10063 = 3'h4 == state ? ram_0_37 : _GEN_9035; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10064 = 3'h4 == state ? ram_0_38 : _GEN_9036; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10065 = 3'h4 == state ? ram_0_39 : _GEN_9037; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10066 = 3'h4 == state ? ram_0_40 : _GEN_9038; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10067 = 3'h4 == state ? ram_0_41 : _GEN_9039; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10068 = 3'h4 == state ? ram_0_42 : _GEN_9040; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10069 = 3'h4 == state ? ram_0_43 : _GEN_9041; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10070 = 3'h4 == state ? ram_0_44 : _GEN_9042; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10071 = 3'h4 == state ? ram_0_45 : _GEN_9043; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10072 = 3'h4 == state ? ram_0_46 : _GEN_9044; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10073 = 3'h4 == state ? ram_0_47 : _GEN_9045; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10074 = 3'h4 == state ? ram_0_48 : _GEN_9046; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10075 = 3'h4 == state ? ram_0_49 : _GEN_9047; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10076 = 3'h4 == state ? ram_0_50 : _GEN_9048; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10077 = 3'h4 == state ? ram_0_51 : _GEN_9049; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10078 = 3'h4 == state ? ram_0_52 : _GEN_9050; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10079 = 3'h4 == state ? ram_0_53 : _GEN_9051; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10080 = 3'h4 == state ? ram_0_54 : _GEN_9052; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10081 = 3'h4 == state ? ram_0_55 : _GEN_9053; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10082 = 3'h4 == state ? ram_0_56 : _GEN_9054; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10083 = 3'h4 == state ? ram_0_57 : _GEN_9055; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10084 = 3'h4 == state ? ram_0_58 : _GEN_9056; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10085 = 3'h4 == state ? ram_0_59 : _GEN_9057; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10086 = 3'h4 == state ? ram_0_60 : _GEN_9058; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10087 = 3'h4 == state ? ram_0_61 : _GEN_9059; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10088 = 3'h4 == state ? ram_0_62 : _GEN_9060; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10089 = 3'h4 == state ? ram_0_63 : _GEN_9061; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10090 = 3'h4 == state ? ram_0_64 : _GEN_9062; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10091 = 3'h4 == state ? ram_0_65 : _GEN_9063; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10092 = 3'h4 == state ? ram_0_66 : _GEN_9064; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10093 = 3'h4 == state ? ram_0_67 : _GEN_9065; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10094 = 3'h4 == state ? ram_0_68 : _GEN_9066; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10095 = 3'h4 == state ? ram_0_69 : _GEN_9067; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10096 = 3'h4 == state ? ram_0_70 : _GEN_9068; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10097 = 3'h4 == state ? ram_0_71 : _GEN_9069; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10098 = 3'h4 == state ? ram_0_72 : _GEN_9070; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10099 = 3'h4 == state ? ram_0_73 : _GEN_9071; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10100 = 3'h4 == state ? ram_0_74 : _GEN_9072; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10101 = 3'h4 == state ? ram_0_75 : _GEN_9073; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10102 = 3'h4 == state ? ram_0_76 : _GEN_9074; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10103 = 3'h4 == state ? ram_0_77 : _GEN_9075; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10104 = 3'h4 == state ? ram_0_78 : _GEN_9076; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10105 = 3'h4 == state ? ram_0_79 : _GEN_9077; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10106 = 3'h4 == state ? ram_0_80 : _GEN_9078; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10107 = 3'h4 == state ? ram_0_81 : _GEN_9079; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10108 = 3'h4 == state ? ram_0_82 : _GEN_9080; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10109 = 3'h4 == state ? ram_0_83 : _GEN_9081; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10110 = 3'h4 == state ? ram_0_84 : _GEN_9082; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10111 = 3'h4 == state ? ram_0_85 : _GEN_9083; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10112 = 3'h4 == state ? ram_0_86 : _GEN_9084; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10113 = 3'h4 == state ? ram_0_87 : _GEN_9085; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10114 = 3'h4 == state ? ram_0_88 : _GEN_9086; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10115 = 3'h4 == state ? ram_0_89 : _GEN_9087; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10116 = 3'h4 == state ? ram_0_90 : _GEN_9088; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10117 = 3'h4 == state ? ram_0_91 : _GEN_9089; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10118 = 3'h4 == state ? ram_0_92 : _GEN_9090; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10119 = 3'h4 == state ? ram_0_93 : _GEN_9091; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10120 = 3'h4 == state ? ram_0_94 : _GEN_9092; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10121 = 3'h4 == state ? ram_0_95 : _GEN_9093; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10122 = 3'h4 == state ? ram_0_96 : _GEN_9094; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10123 = 3'h4 == state ? ram_0_97 : _GEN_9095; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10124 = 3'h4 == state ? ram_0_98 : _GEN_9096; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10125 = 3'h4 == state ? ram_0_99 : _GEN_9097; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10126 = 3'h4 == state ? ram_0_100 : _GEN_9098; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10127 = 3'h4 == state ? ram_0_101 : _GEN_9099; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10128 = 3'h4 == state ? ram_0_102 : _GEN_9100; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10129 = 3'h4 == state ? ram_0_103 : _GEN_9101; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10130 = 3'h4 == state ? ram_0_104 : _GEN_9102; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10131 = 3'h4 == state ? ram_0_105 : _GEN_9103; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10132 = 3'h4 == state ? ram_0_106 : _GEN_9104; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10133 = 3'h4 == state ? ram_0_107 : _GEN_9105; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10134 = 3'h4 == state ? ram_0_108 : _GEN_9106; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10135 = 3'h4 == state ? ram_0_109 : _GEN_9107; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10136 = 3'h4 == state ? ram_0_110 : _GEN_9108; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10137 = 3'h4 == state ? ram_0_111 : _GEN_9109; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10138 = 3'h4 == state ? ram_0_112 : _GEN_9110; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10139 = 3'h4 == state ? ram_0_113 : _GEN_9111; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10140 = 3'h4 == state ? ram_0_114 : _GEN_9112; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10141 = 3'h4 == state ? ram_0_115 : _GEN_9113; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10142 = 3'h4 == state ? ram_0_116 : _GEN_9114; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10143 = 3'h4 == state ? ram_0_117 : _GEN_9115; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10144 = 3'h4 == state ? ram_0_118 : _GEN_9116; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10145 = 3'h4 == state ? ram_0_119 : _GEN_9117; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10146 = 3'h4 == state ? ram_0_120 : _GEN_9118; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10147 = 3'h4 == state ? ram_0_121 : _GEN_9119; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10148 = 3'h4 == state ? ram_0_122 : _GEN_9120; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10149 = 3'h4 == state ? ram_0_123 : _GEN_9121; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10150 = 3'h4 == state ? ram_0_124 : _GEN_9122; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10151 = 3'h4 == state ? ram_0_125 : _GEN_9123; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10152 = 3'h4 == state ? ram_0_126 : _GEN_9124; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_10153 = 3'h4 == state ? ram_0_127 : _GEN_9125; // @[d_cache.scala 64:18 18:24]
  wire [31:0] _GEN_10154 = 3'h4 == state ? tag_0_0 : _GEN_9126; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10155 = 3'h4 == state ? tag_0_1 : _GEN_9127; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10156 = 3'h4 == state ? tag_0_2 : _GEN_9128; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10157 = 3'h4 == state ? tag_0_3 : _GEN_9129; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10158 = 3'h4 == state ? tag_0_4 : _GEN_9130; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10159 = 3'h4 == state ? tag_0_5 : _GEN_9131; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10160 = 3'h4 == state ? tag_0_6 : _GEN_9132; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10161 = 3'h4 == state ? tag_0_7 : _GEN_9133; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10162 = 3'h4 == state ? tag_0_8 : _GEN_9134; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10163 = 3'h4 == state ? tag_0_9 : _GEN_9135; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10164 = 3'h4 == state ? tag_0_10 : _GEN_9136; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10165 = 3'h4 == state ? tag_0_11 : _GEN_9137; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10166 = 3'h4 == state ? tag_0_12 : _GEN_9138; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10167 = 3'h4 == state ? tag_0_13 : _GEN_9139; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10168 = 3'h4 == state ? tag_0_14 : _GEN_9140; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10169 = 3'h4 == state ? tag_0_15 : _GEN_9141; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10170 = 3'h4 == state ? tag_0_16 : _GEN_9142; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10171 = 3'h4 == state ? tag_0_17 : _GEN_9143; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10172 = 3'h4 == state ? tag_0_18 : _GEN_9144; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10173 = 3'h4 == state ? tag_0_19 : _GEN_9145; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10174 = 3'h4 == state ? tag_0_20 : _GEN_9146; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10175 = 3'h4 == state ? tag_0_21 : _GEN_9147; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10176 = 3'h4 == state ? tag_0_22 : _GEN_9148; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10177 = 3'h4 == state ? tag_0_23 : _GEN_9149; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10178 = 3'h4 == state ? tag_0_24 : _GEN_9150; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10179 = 3'h4 == state ? tag_0_25 : _GEN_9151; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10180 = 3'h4 == state ? tag_0_26 : _GEN_9152; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10181 = 3'h4 == state ? tag_0_27 : _GEN_9153; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10182 = 3'h4 == state ? tag_0_28 : _GEN_9154; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10183 = 3'h4 == state ? tag_0_29 : _GEN_9155; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10184 = 3'h4 == state ? tag_0_30 : _GEN_9156; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10185 = 3'h4 == state ? tag_0_31 : _GEN_9157; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10186 = 3'h4 == state ? tag_0_32 : _GEN_9158; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10187 = 3'h4 == state ? tag_0_33 : _GEN_9159; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10188 = 3'h4 == state ? tag_0_34 : _GEN_9160; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10189 = 3'h4 == state ? tag_0_35 : _GEN_9161; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10190 = 3'h4 == state ? tag_0_36 : _GEN_9162; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10191 = 3'h4 == state ? tag_0_37 : _GEN_9163; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10192 = 3'h4 == state ? tag_0_38 : _GEN_9164; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10193 = 3'h4 == state ? tag_0_39 : _GEN_9165; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10194 = 3'h4 == state ? tag_0_40 : _GEN_9166; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10195 = 3'h4 == state ? tag_0_41 : _GEN_9167; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10196 = 3'h4 == state ? tag_0_42 : _GEN_9168; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10197 = 3'h4 == state ? tag_0_43 : _GEN_9169; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10198 = 3'h4 == state ? tag_0_44 : _GEN_9170; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10199 = 3'h4 == state ? tag_0_45 : _GEN_9171; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10200 = 3'h4 == state ? tag_0_46 : _GEN_9172; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10201 = 3'h4 == state ? tag_0_47 : _GEN_9173; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10202 = 3'h4 == state ? tag_0_48 : _GEN_9174; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10203 = 3'h4 == state ? tag_0_49 : _GEN_9175; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10204 = 3'h4 == state ? tag_0_50 : _GEN_9176; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10205 = 3'h4 == state ? tag_0_51 : _GEN_9177; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10206 = 3'h4 == state ? tag_0_52 : _GEN_9178; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10207 = 3'h4 == state ? tag_0_53 : _GEN_9179; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10208 = 3'h4 == state ? tag_0_54 : _GEN_9180; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10209 = 3'h4 == state ? tag_0_55 : _GEN_9181; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10210 = 3'h4 == state ? tag_0_56 : _GEN_9182; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10211 = 3'h4 == state ? tag_0_57 : _GEN_9183; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10212 = 3'h4 == state ? tag_0_58 : _GEN_9184; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10213 = 3'h4 == state ? tag_0_59 : _GEN_9185; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10214 = 3'h4 == state ? tag_0_60 : _GEN_9186; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10215 = 3'h4 == state ? tag_0_61 : _GEN_9187; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10216 = 3'h4 == state ? tag_0_62 : _GEN_9188; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10217 = 3'h4 == state ? tag_0_63 : _GEN_9189; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10218 = 3'h4 == state ? tag_0_64 : _GEN_9190; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10219 = 3'h4 == state ? tag_0_65 : _GEN_9191; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10220 = 3'h4 == state ? tag_0_66 : _GEN_9192; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10221 = 3'h4 == state ? tag_0_67 : _GEN_9193; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10222 = 3'h4 == state ? tag_0_68 : _GEN_9194; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10223 = 3'h4 == state ? tag_0_69 : _GEN_9195; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10224 = 3'h4 == state ? tag_0_70 : _GEN_9196; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10225 = 3'h4 == state ? tag_0_71 : _GEN_9197; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10226 = 3'h4 == state ? tag_0_72 : _GEN_9198; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10227 = 3'h4 == state ? tag_0_73 : _GEN_9199; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10228 = 3'h4 == state ? tag_0_74 : _GEN_9200; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10229 = 3'h4 == state ? tag_0_75 : _GEN_9201; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10230 = 3'h4 == state ? tag_0_76 : _GEN_9202; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10231 = 3'h4 == state ? tag_0_77 : _GEN_9203; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10232 = 3'h4 == state ? tag_0_78 : _GEN_9204; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10233 = 3'h4 == state ? tag_0_79 : _GEN_9205; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10234 = 3'h4 == state ? tag_0_80 : _GEN_9206; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10235 = 3'h4 == state ? tag_0_81 : _GEN_9207; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10236 = 3'h4 == state ? tag_0_82 : _GEN_9208; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10237 = 3'h4 == state ? tag_0_83 : _GEN_9209; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10238 = 3'h4 == state ? tag_0_84 : _GEN_9210; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10239 = 3'h4 == state ? tag_0_85 : _GEN_9211; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10240 = 3'h4 == state ? tag_0_86 : _GEN_9212; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10241 = 3'h4 == state ? tag_0_87 : _GEN_9213; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10242 = 3'h4 == state ? tag_0_88 : _GEN_9214; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10243 = 3'h4 == state ? tag_0_89 : _GEN_9215; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10244 = 3'h4 == state ? tag_0_90 : _GEN_9216; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10245 = 3'h4 == state ? tag_0_91 : _GEN_9217; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10246 = 3'h4 == state ? tag_0_92 : _GEN_9218; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10247 = 3'h4 == state ? tag_0_93 : _GEN_9219; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10248 = 3'h4 == state ? tag_0_94 : _GEN_9220; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10249 = 3'h4 == state ? tag_0_95 : _GEN_9221; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10250 = 3'h4 == state ? tag_0_96 : _GEN_9222; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10251 = 3'h4 == state ? tag_0_97 : _GEN_9223; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10252 = 3'h4 == state ? tag_0_98 : _GEN_9224; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10253 = 3'h4 == state ? tag_0_99 : _GEN_9225; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10254 = 3'h4 == state ? tag_0_100 : _GEN_9226; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10255 = 3'h4 == state ? tag_0_101 : _GEN_9227; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10256 = 3'h4 == state ? tag_0_102 : _GEN_9228; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10257 = 3'h4 == state ? tag_0_103 : _GEN_9229; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10258 = 3'h4 == state ? tag_0_104 : _GEN_9230; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10259 = 3'h4 == state ? tag_0_105 : _GEN_9231; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10260 = 3'h4 == state ? tag_0_106 : _GEN_9232; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10261 = 3'h4 == state ? tag_0_107 : _GEN_9233; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10262 = 3'h4 == state ? tag_0_108 : _GEN_9234; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10263 = 3'h4 == state ? tag_0_109 : _GEN_9235; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10264 = 3'h4 == state ? tag_0_110 : _GEN_9236; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10265 = 3'h4 == state ? tag_0_111 : _GEN_9237; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10266 = 3'h4 == state ? tag_0_112 : _GEN_9238; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10267 = 3'h4 == state ? tag_0_113 : _GEN_9239; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10268 = 3'h4 == state ? tag_0_114 : _GEN_9240; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10269 = 3'h4 == state ? tag_0_115 : _GEN_9241; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10270 = 3'h4 == state ? tag_0_116 : _GEN_9242; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10271 = 3'h4 == state ? tag_0_117 : _GEN_9243; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10272 = 3'h4 == state ? tag_0_118 : _GEN_9244; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10273 = 3'h4 == state ? tag_0_119 : _GEN_9245; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10274 = 3'h4 == state ? tag_0_120 : _GEN_9246; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10275 = 3'h4 == state ? tag_0_121 : _GEN_9247; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10276 = 3'h4 == state ? tag_0_122 : _GEN_9248; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10277 = 3'h4 == state ? tag_0_123 : _GEN_9249; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10278 = 3'h4 == state ? tag_0_124 : _GEN_9250; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10279 = 3'h4 == state ? tag_0_125 : _GEN_9251; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10280 = 3'h4 == state ? tag_0_126 : _GEN_9252; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_10281 = 3'h4 == state ? tag_0_127 : _GEN_9253; // @[d_cache.scala 64:18 20:24]
  wire  _GEN_10282 = 3'h4 == state ? valid_0_0 : _GEN_9254; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10283 = 3'h4 == state ? valid_0_1 : _GEN_9255; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10284 = 3'h4 == state ? valid_0_2 : _GEN_9256; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10285 = 3'h4 == state ? valid_0_3 : _GEN_9257; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10286 = 3'h4 == state ? valid_0_4 : _GEN_9258; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10287 = 3'h4 == state ? valid_0_5 : _GEN_9259; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10288 = 3'h4 == state ? valid_0_6 : _GEN_9260; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10289 = 3'h4 == state ? valid_0_7 : _GEN_9261; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10290 = 3'h4 == state ? valid_0_8 : _GEN_9262; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10291 = 3'h4 == state ? valid_0_9 : _GEN_9263; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10292 = 3'h4 == state ? valid_0_10 : _GEN_9264; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10293 = 3'h4 == state ? valid_0_11 : _GEN_9265; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10294 = 3'h4 == state ? valid_0_12 : _GEN_9266; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10295 = 3'h4 == state ? valid_0_13 : _GEN_9267; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10296 = 3'h4 == state ? valid_0_14 : _GEN_9268; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10297 = 3'h4 == state ? valid_0_15 : _GEN_9269; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10298 = 3'h4 == state ? valid_0_16 : _GEN_9270; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10299 = 3'h4 == state ? valid_0_17 : _GEN_9271; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10300 = 3'h4 == state ? valid_0_18 : _GEN_9272; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10301 = 3'h4 == state ? valid_0_19 : _GEN_9273; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10302 = 3'h4 == state ? valid_0_20 : _GEN_9274; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10303 = 3'h4 == state ? valid_0_21 : _GEN_9275; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10304 = 3'h4 == state ? valid_0_22 : _GEN_9276; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10305 = 3'h4 == state ? valid_0_23 : _GEN_9277; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10306 = 3'h4 == state ? valid_0_24 : _GEN_9278; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10307 = 3'h4 == state ? valid_0_25 : _GEN_9279; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10308 = 3'h4 == state ? valid_0_26 : _GEN_9280; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10309 = 3'h4 == state ? valid_0_27 : _GEN_9281; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10310 = 3'h4 == state ? valid_0_28 : _GEN_9282; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10311 = 3'h4 == state ? valid_0_29 : _GEN_9283; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10312 = 3'h4 == state ? valid_0_30 : _GEN_9284; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10313 = 3'h4 == state ? valid_0_31 : _GEN_9285; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10314 = 3'h4 == state ? valid_0_32 : _GEN_9286; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10315 = 3'h4 == state ? valid_0_33 : _GEN_9287; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10316 = 3'h4 == state ? valid_0_34 : _GEN_9288; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10317 = 3'h4 == state ? valid_0_35 : _GEN_9289; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10318 = 3'h4 == state ? valid_0_36 : _GEN_9290; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10319 = 3'h4 == state ? valid_0_37 : _GEN_9291; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10320 = 3'h4 == state ? valid_0_38 : _GEN_9292; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10321 = 3'h4 == state ? valid_0_39 : _GEN_9293; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10322 = 3'h4 == state ? valid_0_40 : _GEN_9294; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10323 = 3'h4 == state ? valid_0_41 : _GEN_9295; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10324 = 3'h4 == state ? valid_0_42 : _GEN_9296; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10325 = 3'h4 == state ? valid_0_43 : _GEN_9297; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10326 = 3'h4 == state ? valid_0_44 : _GEN_9298; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10327 = 3'h4 == state ? valid_0_45 : _GEN_9299; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10328 = 3'h4 == state ? valid_0_46 : _GEN_9300; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10329 = 3'h4 == state ? valid_0_47 : _GEN_9301; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10330 = 3'h4 == state ? valid_0_48 : _GEN_9302; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10331 = 3'h4 == state ? valid_0_49 : _GEN_9303; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10332 = 3'h4 == state ? valid_0_50 : _GEN_9304; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10333 = 3'h4 == state ? valid_0_51 : _GEN_9305; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10334 = 3'h4 == state ? valid_0_52 : _GEN_9306; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10335 = 3'h4 == state ? valid_0_53 : _GEN_9307; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10336 = 3'h4 == state ? valid_0_54 : _GEN_9308; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10337 = 3'h4 == state ? valid_0_55 : _GEN_9309; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10338 = 3'h4 == state ? valid_0_56 : _GEN_9310; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10339 = 3'h4 == state ? valid_0_57 : _GEN_9311; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10340 = 3'h4 == state ? valid_0_58 : _GEN_9312; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10341 = 3'h4 == state ? valid_0_59 : _GEN_9313; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10342 = 3'h4 == state ? valid_0_60 : _GEN_9314; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10343 = 3'h4 == state ? valid_0_61 : _GEN_9315; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10344 = 3'h4 == state ? valid_0_62 : _GEN_9316; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10345 = 3'h4 == state ? valid_0_63 : _GEN_9317; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10346 = 3'h4 == state ? valid_0_64 : _GEN_9318; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10347 = 3'h4 == state ? valid_0_65 : _GEN_9319; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10348 = 3'h4 == state ? valid_0_66 : _GEN_9320; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10349 = 3'h4 == state ? valid_0_67 : _GEN_9321; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10350 = 3'h4 == state ? valid_0_68 : _GEN_9322; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10351 = 3'h4 == state ? valid_0_69 : _GEN_9323; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10352 = 3'h4 == state ? valid_0_70 : _GEN_9324; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10353 = 3'h4 == state ? valid_0_71 : _GEN_9325; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10354 = 3'h4 == state ? valid_0_72 : _GEN_9326; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10355 = 3'h4 == state ? valid_0_73 : _GEN_9327; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10356 = 3'h4 == state ? valid_0_74 : _GEN_9328; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10357 = 3'h4 == state ? valid_0_75 : _GEN_9329; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10358 = 3'h4 == state ? valid_0_76 : _GEN_9330; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10359 = 3'h4 == state ? valid_0_77 : _GEN_9331; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10360 = 3'h4 == state ? valid_0_78 : _GEN_9332; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10361 = 3'h4 == state ? valid_0_79 : _GEN_9333; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10362 = 3'h4 == state ? valid_0_80 : _GEN_9334; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10363 = 3'h4 == state ? valid_0_81 : _GEN_9335; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10364 = 3'h4 == state ? valid_0_82 : _GEN_9336; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10365 = 3'h4 == state ? valid_0_83 : _GEN_9337; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10366 = 3'h4 == state ? valid_0_84 : _GEN_9338; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10367 = 3'h4 == state ? valid_0_85 : _GEN_9339; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10368 = 3'h4 == state ? valid_0_86 : _GEN_9340; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10369 = 3'h4 == state ? valid_0_87 : _GEN_9341; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10370 = 3'h4 == state ? valid_0_88 : _GEN_9342; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10371 = 3'h4 == state ? valid_0_89 : _GEN_9343; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10372 = 3'h4 == state ? valid_0_90 : _GEN_9344; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10373 = 3'h4 == state ? valid_0_91 : _GEN_9345; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10374 = 3'h4 == state ? valid_0_92 : _GEN_9346; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10375 = 3'h4 == state ? valid_0_93 : _GEN_9347; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10376 = 3'h4 == state ? valid_0_94 : _GEN_9348; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10377 = 3'h4 == state ? valid_0_95 : _GEN_9349; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10378 = 3'h4 == state ? valid_0_96 : _GEN_9350; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10379 = 3'h4 == state ? valid_0_97 : _GEN_9351; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10380 = 3'h4 == state ? valid_0_98 : _GEN_9352; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10381 = 3'h4 == state ? valid_0_99 : _GEN_9353; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10382 = 3'h4 == state ? valid_0_100 : _GEN_9354; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10383 = 3'h4 == state ? valid_0_101 : _GEN_9355; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10384 = 3'h4 == state ? valid_0_102 : _GEN_9356; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10385 = 3'h4 == state ? valid_0_103 : _GEN_9357; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10386 = 3'h4 == state ? valid_0_104 : _GEN_9358; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10387 = 3'h4 == state ? valid_0_105 : _GEN_9359; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10388 = 3'h4 == state ? valid_0_106 : _GEN_9360; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10389 = 3'h4 == state ? valid_0_107 : _GEN_9361; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10390 = 3'h4 == state ? valid_0_108 : _GEN_9362; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10391 = 3'h4 == state ? valid_0_109 : _GEN_9363; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10392 = 3'h4 == state ? valid_0_110 : _GEN_9364; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10393 = 3'h4 == state ? valid_0_111 : _GEN_9365; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10394 = 3'h4 == state ? valid_0_112 : _GEN_9366; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10395 = 3'h4 == state ? valid_0_113 : _GEN_9367; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10396 = 3'h4 == state ? valid_0_114 : _GEN_9368; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10397 = 3'h4 == state ? valid_0_115 : _GEN_9369; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10398 = 3'h4 == state ? valid_0_116 : _GEN_9370; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10399 = 3'h4 == state ? valid_0_117 : _GEN_9371; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10400 = 3'h4 == state ? valid_0_118 : _GEN_9372; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10401 = 3'h4 == state ? valid_0_119 : _GEN_9373; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10402 = 3'h4 == state ? valid_0_120 : _GEN_9374; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10403 = 3'h4 == state ? valid_0_121 : _GEN_9375; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10404 = 3'h4 == state ? valid_0_122 : _GEN_9376; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10405 = 3'h4 == state ? valid_0_123 : _GEN_9377; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10406 = 3'h4 == state ? valid_0_124 : _GEN_9378; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10407 = 3'h4 == state ? valid_0_125 : _GEN_9379; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10408 = 3'h4 == state ? valid_0_126 : _GEN_9380; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10409 = 3'h4 == state ? valid_0_127 : _GEN_9381; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_10410 = 3'h4 == state ? quene : _GEN_9382; // @[d_cache.scala 64:18 35:24]
  wire [63:0] _GEN_10411 = 3'h4 == state ? ram_1_0 : _GEN_9383; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10412 = 3'h4 == state ? ram_1_1 : _GEN_9384; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10413 = 3'h4 == state ? ram_1_2 : _GEN_9385; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10414 = 3'h4 == state ? ram_1_3 : _GEN_9386; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10415 = 3'h4 == state ? ram_1_4 : _GEN_9387; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10416 = 3'h4 == state ? ram_1_5 : _GEN_9388; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10417 = 3'h4 == state ? ram_1_6 : _GEN_9389; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10418 = 3'h4 == state ? ram_1_7 : _GEN_9390; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10419 = 3'h4 == state ? ram_1_8 : _GEN_9391; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10420 = 3'h4 == state ? ram_1_9 : _GEN_9392; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10421 = 3'h4 == state ? ram_1_10 : _GEN_9393; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10422 = 3'h4 == state ? ram_1_11 : _GEN_9394; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10423 = 3'h4 == state ? ram_1_12 : _GEN_9395; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10424 = 3'h4 == state ? ram_1_13 : _GEN_9396; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10425 = 3'h4 == state ? ram_1_14 : _GEN_9397; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10426 = 3'h4 == state ? ram_1_15 : _GEN_9398; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10427 = 3'h4 == state ? ram_1_16 : _GEN_9399; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10428 = 3'h4 == state ? ram_1_17 : _GEN_9400; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10429 = 3'h4 == state ? ram_1_18 : _GEN_9401; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10430 = 3'h4 == state ? ram_1_19 : _GEN_9402; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10431 = 3'h4 == state ? ram_1_20 : _GEN_9403; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10432 = 3'h4 == state ? ram_1_21 : _GEN_9404; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10433 = 3'h4 == state ? ram_1_22 : _GEN_9405; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10434 = 3'h4 == state ? ram_1_23 : _GEN_9406; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10435 = 3'h4 == state ? ram_1_24 : _GEN_9407; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10436 = 3'h4 == state ? ram_1_25 : _GEN_9408; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10437 = 3'h4 == state ? ram_1_26 : _GEN_9409; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10438 = 3'h4 == state ? ram_1_27 : _GEN_9410; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10439 = 3'h4 == state ? ram_1_28 : _GEN_9411; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10440 = 3'h4 == state ? ram_1_29 : _GEN_9412; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10441 = 3'h4 == state ? ram_1_30 : _GEN_9413; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10442 = 3'h4 == state ? ram_1_31 : _GEN_9414; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10443 = 3'h4 == state ? ram_1_32 : _GEN_9415; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10444 = 3'h4 == state ? ram_1_33 : _GEN_9416; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10445 = 3'h4 == state ? ram_1_34 : _GEN_9417; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10446 = 3'h4 == state ? ram_1_35 : _GEN_9418; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10447 = 3'h4 == state ? ram_1_36 : _GEN_9419; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10448 = 3'h4 == state ? ram_1_37 : _GEN_9420; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10449 = 3'h4 == state ? ram_1_38 : _GEN_9421; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10450 = 3'h4 == state ? ram_1_39 : _GEN_9422; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10451 = 3'h4 == state ? ram_1_40 : _GEN_9423; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10452 = 3'h4 == state ? ram_1_41 : _GEN_9424; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10453 = 3'h4 == state ? ram_1_42 : _GEN_9425; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10454 = 3'h4 == state ? ram_1_43 : _GEN_9426; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10455 = 3'h4 == state ? ram_1_44 : _GEN_9427; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10456 = 3'h4 == state ? ram_1_45 : _GEN_9428; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10457 = 3'h4 == state ? ram_1_46 : _GEN_9429; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10458 = 3'h4 == state ? ram_1_47 : _GEN_9430; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10459 = 3'h4 == state ? ram_1_48 : _GEN_9431; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10460 = 3'h4 == state ? ram_1_49 : _GEN_9432; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10461 = 3'h4 == state ? ram_1_50 : _GEN_9433; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10462 = 3'h4 == state ? ram_1_51 : _GEN_9434; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10463 = 3'h4 == state ? ram_1_52 : _GEN_9435; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10464 = 3'h4 == state ? ram_1_53 : _GEN_9436; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10465 = 3'h4 == state ? ram_1_54 : _GEN_9437; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10466 = 3'h4 == state ? ram_1_55 : _GEN_9438; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10467 = 3'h4 == state ? ram_1_56 : _GEN_9439; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10468 = 3'h4 == state ? ram_1_57 : _GEN_9440; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10469 = 3'h4 == state ? ram_1_58 : _GEN_9441; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10470 = 3'h4 == state ? ram_1_59 : _GEN_9442; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10471 = 3'h4 == state ? ram_1_60 : _GEN_9443; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10472 = 3'h4 == state ? ram_1_61 : _GEN_9444; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10473 = 3'h4 == state ? ram_1_62 : _GEN_9445; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10474 = 3'h4 == state ? ram_1_63 : _GEN_9446; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10475 = 3'h4 == state ? ram_1_64 : _GEN_9447; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10476 = 3'h4 == state ? ram_1_65 : _GEN_9448; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10477 = 3'h4 == state ? ram_1_66 : _GEN_9449; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10478 = 3'h4 == state ? ram_1_67 : _GEN_9450; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10479 = 3'h4 == state ? ram_1_68 : _GEN_9451; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10480 = 3'h4 == state ? ram_1_69 : _GEN_9452; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10481 = 3'h4 == state ? ram_1_70 : _GEN_9453; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10482 = 3'h4 == state ? ram_1_71 : _GEN_9454; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10483 = 3'h4 == state ? ram_1_72 : _GEN_9455; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10484 = 3'h4 == state ? ram_1_73 : _GEN_9456; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10485 = 3'h4 == state ? ram_1_74 : _GEN_9457; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10486 = 3'h4 == state ? ram_1_75 : _GEN_9458; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10487 = 3'h4 == state ? ram_1_76 : _GEN_9459; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10488 = 3'h4 == state ? ram_1_77 : _GEN_9460; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10489 = 3'h4 == state ? ram_1_78 : _GEN_9461; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10490 = 3'h4 == state ? ram_1_79 : _GEN_9462; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10491 = 3'h4 == state ? ram_1_80 : _GEN_9463; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10492 = 3'h4 == state ? ram_1_81 : _GEN_9464; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10493 = 3'h4 == state ? ram_1_82 : _GEN_9465; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10494 = 3'h4 == state ? ram_1_83 : _GEN_9466; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10495 = 3'h4 == state ? ram_1_84 : _GEN_9467; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10496 = 3'h4 == state ? ram_1_85 : _GEN_9468; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10497 = 3'h4 == state ? ram_1_86 : _GEN_9469; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10498 = 3'h4 == state ? ram_1_87 : _GEN_9470; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10499 = 3'h4 == state ? ram_1_88 : _GEN_9471; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10500 = 3'h4 == state ? ram_1_89 : _GEN_9472; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10501 = 3'h4 == state ? ram_1_90 : _GEN_9473; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10502 = 3'h4 == state ? ram_1_91 : _GEN_9474; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10503 = 3'h4 == state ? ram_1_92 : _GEN_9475; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10504 = 3'h4 == state ? ram_1_93 : _GEN_9476; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10505 = 3'h4 == state ? ram_1_94 : _GEN_9477; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10506 = 3'h4 == state ? ram_1_95 : _GEN_9478; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10507 = 3'h4 == state ? ram_1_96 : _GEN_9479; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10508 = 3'h4 == state ? ram_1_97 : _GEN_9480; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10509 = 3'h4 == state ? ram_1_98 : _GEN_9481; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10510 = 3'h4 == state ? ram_1_99 : _GEN_9482; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10511 = 3'h4 == state ? ram_1_100 : _GEN_9483; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10512 = 3'h4 == state ? ram_1_101 : _GEN_9484; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10513 = 3'h4 == state ? ram_1_102 : _GEN_9485; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10514 = 3'h4 == state ? ram_1_103 : _GEN_9486; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10515 = 3'h4 == state ? ram_1_104 : _GEN_9487; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10516 = 3'h4 == state ? ram_1_105 : _GEN_9488; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10517 = 3'h4 == state ? ram_1_106 : _GEN_9489; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10518 = 3'h4 == state ? ram_1_107 : _GEN_9490; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10519 = 3'h4 == state ? ram_1_108 : _GEN_9491; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10520 = 3'h4 == state ? ram_1_109 : _GEN_9492; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10521 = 3'h4 == state ? ram_1_110 : _GEN_9493; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10522 = 3'h4 == state ? ram_1_111 : _GEN_9494; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10523 = 3'h4 == state ? ram_1_112 : _GEN_9495; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10524 = 3'h4 == state ? ram_1_113 : _GEN_9496; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10525 = 3'h4 == state ? ram_1_114 : _GEN_9497; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10526 = 3'h4 == state ? ram_1_115 : _GEN_9498; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10527 = 3'h4 == state ? ram_1_116 : _GEN_9499; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10528 = 3'h4 == state ? ram_1_117 : _GEN_9500; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10529 = 3'h4 == state ? ram_1_118 : _GEN_9501; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10530 = 3'h4 == state ? ram_1_119 : _GEN_9502; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10531 = 3'h4 == state ? ram_1_120 : _GEN_9503; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10532 = 3'h4 == state ? ram_1_121 : _GEN_9504; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10533 = 3'h4 == state ? ram_1_122 : _GEN_9505; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10534 = 3'h4 == state ? ram_1_123 : _GEN_9506; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10535 = 3'h4 == state ? ram_1_124 : _GEN_9507; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10536 = 3'h4 == state ? ram_1_125 : _GEN_9508; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10537 = 3'h4 == state ? ram_1_126 : _GEN_9509; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_10538 = 3'h4 == state ? ram_1_127 : _GEN_9510; // @[d_cache.scala 64:18 19:24]
  wire [31:0] _GEN_10539 = 3'h4 == state ? tag_1_0 : _GEN_9511; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10540 = 3'h4 == state ? tag_1_1 : _GEN_9512; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10541 = 3'h4 == state ? tag_1_2 : _GEN_9513; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10542 = 3'h4 == state ? tag_1_3 : _GEN_9514; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10543 = 3'h4 == state ? tag_1_4 : _GEN_9515; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10544 = 3'h4 == state ? tag_1_5 : _GEN_9516; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10545 = 3'h4 == state ? tag_1_6 : _GEN_9517; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10546 = 3'h4 == state ? tag_1_7 : _GEN_9518; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10547 = 3'h4 == state ? tag_1_8 : _GEN_9519; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10548 = 3'h4 == state ? tag_1_9 : _GEN_9520; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10549 = 3'h4 == state ? tag_1_10 : _GEN_9521; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10550 = 3'h4 == state ? tag_1_11 : _GEN_9522; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10551 = 3'h4 == state ? tag_1_12 : _GEN_9523; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10552 = 3'h4 == state ? tag_1_13 : _GEN_9524; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10553 = 3'h4 == state ? tag_1_14 : _GEN_9525; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10554 = 3'h4 == state ? tag_1_15 : _GEN_9526; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10555 = 3'h4 == state ? tag_1_16 : _GEN_9527; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10556 = 3'h4 == state ? tag_1_17 : _GEN_9528; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10557 = 3'h4 == state ? tag_1_18 : _GEN_9529; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10558 = 3'h4 == state ? tag_1_19 : _GEN_9530; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10559 = 3'h4 == state ? tag_1_20 : _GEN_9531; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10560 = 3'h4 == state ? tag_1_21 : _GEN_9532; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10561 = 3'h4 == state ? tag_1_22 : _GEN_9533; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10562 = 3'h4 == state ? tag_1_23 : _GEN_9534; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10563 = 3'h4 == state ? tag_1_24 : _GEN_9535; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10564 = 3'h4 == state ? tag_1_25 : _GEN_9536; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10565 = 3'h4 == state ? tag_1_26 : _GEN_9537; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10566 = 3'h4 == state ? tag_1_27 : _GEN_9538; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10567 = 3'h4 == state ? tag_1_28 : _GEN_9539; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10568 = 3'h4 == state ? tag_1_29 : _GEN_9540; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10569 = 3'h4 == state ? tag_1_30 : _GEN_9541; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10570 = 3'h4 == state ? tag_1_31 : _GEN_9542; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10571 = 3'h4 == state ? tag_1_32 : _GEN_9543; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10572 = 3'h4 == state ? tag_1_33 : _GEN_9544; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10573 = 3'h4 == state ? tag_1_34 : _GEN_9545; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10574 = 3'h4 == state ? tag_1_35 : _GEN_9546; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10575 = 3'h4 == state ? tag_1_36 : _GEN_9547; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10576 = 3'h4 == state ? tag_1_37 : _GEN_9548; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10577 = 3'h4 == state ? tag_1_38 : _GEN_9549; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10578 = 3'h4 == state ? tag_1_39 : _GEN_9550; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10579 = 3'h4 == state ? tag_1_40 : _GEN_9551; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10580 = 3'h4 == state ? tag_1_41 : _GEN_9552; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10581 = 3'h4 == state ? tag_1_42 : _GEN_9553; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10582 = 3'h4 == state ? tag_1_43 : _GEN_9554; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10583 = 3'h4 == state ? tag_1_44 : _GEN_9555; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10584 = 3'h4 == state ? tag_1_45 : _GEN_9556; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10585 = 3'h4 == state ? tag_1_46 : _GEN_9557; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10586 = 3'h4 == state ? tag_1_47 : _GEN_9558; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10587 = 3'h4 == state ? tag_1_48 : _GEN_9559; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10588 = 3'h4 == state ? tag_1_49 : _GEN_9560; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10589 = 3'h4 == state ? tag_1_50 : _GEN_9561; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10590 = 3'h4 == state ? tag_1_51 : _GEN_9562; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10591 = 3'h4 == state ? tag_1_52 : _GEN_9563; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10592 = 3'h4 == state ? tag_1_53 : _GEN_9564; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10593 = 3'h4 == state ? tag_1_54 : _GEN_9565; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10594 = 3'h4 == state ? tag_1_55 : _GEN_9566; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10595 = 3'h4 == state ? tag_1_56 : _GEN_9567; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10596 = 3'h4 == state ? tag_1_57 : _GEN_9568; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10597 = 3'h4 == state ? tag_1_58 : _GEN_9569; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10598 = 3'h4 == state ? tag_1_59 : _GEN_9570; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10599 = 3'h4 == state ? tag_1_60 : _GEN_9571; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10600 = 3'h4 == state ? tag_1_61 : _GEN_9572; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10601 = 3'h4 == state ? tag_1_62 : _GEN_9573; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10602 = 3'h4 == state ? tag_1_63 : _GEN_9574; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10603 = 3'h4 == state ? tag_1_64 : _GEN_9575; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10604 = 3'h4 == state ? tag_1_65 : _GEN_9576; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10605 = 3'h4 == state ? tag_1_66 : _GEN_9577; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10606 = 3'h4 == state ? tag_1_67 : _GEN_9578; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10607 = 3'h4 == state ? tag_1_68 : _GEN_9579; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10608 = 3'h4 == state ? tag_1_69 : _GEN_9580; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10609 = 3'h4 == state ? tag_1_70 : _GEN_9581; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10610 = 3'h4 == state ? tag_1_71 : _GEN_9582; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10611 = 3'h4 == state ? tag_1_72 : _GEN_9583; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10612 = 3'h4 == state ? tag_1_73 : _GEN_9584; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10613 = 3'h4 == state ? tag_1_74 : _GEN_9585; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10614 = 3'h4 == state ? tag_1_75 : _GEN_9586; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10615 = 3'h4 == state ? tag_1_76 : _GEN_9587; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10616 = 3'h4 == state ? tag_1_77 : _GEN_9588; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10617 = 3'h4 == state ? tag_1_78 : _GEN_9589; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10618 = 3'h4 == state ? tag_1_79 : _GEN_9590; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10619 = 3'h4 == state ? tag_1_80 : _GEN_9591; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10620 = 3'h4 == state ? tag_1_81 : _GEN_9592; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10621 = 3'h4 == state ? tag_1_82 : _GEN_9593; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10622 = 3'h4 == state ? tag_1_83 : _GEN_9594; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10623 = 3'h4 == state ? tag_1_84 : _GEN_9595; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10624 = 3'h4 == state ? tag_1_85 : _GEN_9596; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10625 = 3'h4 == state ? tag_1_86 : _GEN_9597; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10626 = 3'h4 == state ? tag_1_87 : _GEN_9598; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10627 = 3'h4 == state ? tag_1_88 : _GEN_9599; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10628 = 3'h4 == state ? tag_1_89 : _GEN_9600; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10629 = 3'h4 == state ? tag_1_90 : _GEN_9601; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10630 = 3'h4 == state ? tag_1_91 : _GEN_9602; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10631 = 3'h4 == state ? tag_1_92 : _GEN_9603; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10632 = 3'h4 == state ? tag_1_93 : _GEN_9604; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10633 = 3'h4 == state ? tag_1_94 : _GEN_9605; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10634 = 3'h4 == state ? tag_1_95 : _GEN_9606; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10635 = 3'h4 == state ? tag_1_96 : _GEN_9607; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10636 = 3'h4 == state ? tag_1_97 : _GEN_9608; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10637 = 3'h4 == state ? tag_1_98 : _GEN_9609; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10638 = 3'h4 == state ? tag_1_99 : _GEN_9610; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10639 = 3'h4 == state ? tag_1_100 : _GEN_9611; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10640 = 3'h4 == state ? tag_1_101 : _GEN_9612; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10641 = 3'h4 == state ? tag_1_102 : _GEN_9613; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10642 = 3'h4 == state ? tag_1_103 : _GEN_9614; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10643 = 3'h4 == state ? tag_1_104 : _GEN_9615; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10644 = 3'h4 == state ? tag_1_105 : _GEN_9616; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10645 = 3'h4 == state ? tag_1_106 : _GEN_9617; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10646 = 3'h4 == state ? tag_1_107 : _GEN_9618; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10647 = 3'h4 == state ? tag_1_108 : _GEN_9619; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10648 = 3'h4 == state ? tag_1_109 : _GEN_9620; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10649 = 3'h4 == state ? tag_1_110 : _GEN_9621; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10650 = 3'h4 == state ? tag_1_111 : _GEN_9622; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10651 = 3'h4 == state ? tag_1_112 : _GEN_9623; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10652 = 3'h4 == state ? tag_1_113 : _GEN_9624; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10653 = 3'h4 == state ? tag_1_114 : _GEN_9625; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10654 = 3'h4 == state ? tag_1_115 : _GEN_9626; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10655 = 3'h4 == state ? tag_1_116 : _GEN_9627; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10656 = 3'h4 == state ? tag_1_117 : _GEN_9628; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10657 = 3'h4 == state ? tag_1_118 : _GEN_9629; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10658 = 3'h4 == state ? tag_1_119 : _GEN_9630; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10659 = 3'h4 == state ? tag_1_120 : _GEN_9631; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10660 = 3'h4 == state ? tag_1_121 : _GEN_9632; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10661 = 3'h4 == state ? tag_1_122 : _GEN_9633; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10662 = 3'h4 == state ? tag_1_123 : _GEN_9634; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10663 = 3'h4 == state ? tag_1_124 : _GEN_9635; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10664 = 3'h4 == state ? tag_1_125 : _GEN_9636; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10665 = 3'h4 == state ? tag_1_126 : _GEN_9637; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_10666 = 3'h4 == state ? tag_1_127 : _GEN_9638; // @[d_cache.scala 64:18 21:24]
  wire  _GEN_10667 = 3'h4 == state ? valid_1_0 : _GEN_9639; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10668 = 3'h4 == state ? valid_1_1 : _GEN_9640; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10669 = 3'h4 == state ? valid_1_2 : _GEN_9641; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10670 = 3'h4 == state ? valid_1_3 : _GEN_9642; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10671 = 3'h4 == state ? valid_1_4 : _GEN_9643; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10672 = 3'h4 == state ? valid_1_5 : _GEN_9644; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10673 = 3'h4 == state ? valid_1_6 : _GEN_9645; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10674 = 3'h4 == state ? valid_1_7 : _GEN_9646; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10675 = 3'h4 == state ? valid_1_8 : _GEN_9647; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10676 = 3'h4 == state ? valid_1_9 : _GEN_9648; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10677 = 3'h4 == state ? valid_1_10 : _GEN_9649; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10678 = 3'h4 == state ? valid_1_11 : _GEN_9650; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10679 = 3'h4 == state ? valid_1_12 : _GEN_9651; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10680 = 3'h4 == state ? valid_1_13 : _GEN_9652; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10681 = 3'h4 == state ? valid_1_14 : _GEN_9653; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10682 = 3'h4 == state ? valid_1_15 : _GEN_9654; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10683 = 3'h4 == state ? valid_1_16 : _GEN_9655; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10684 = 3'h4 == state ? valid_1_17 : _GEN_9656; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10685 = 3'h4 == state ? valid_1_18 : _GEN_9657; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10686 = 3'h4 == state ? valid_1_19 : _GEN_9658; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10687 = 3'h4 == state ? valid_1_20 : _GEN_9659; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10688 = 3'h4 == state ? valid_1_21 : _GEN_9660; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10689 = 3'h4 == state ? valid_1_22 : _GEN_9661; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10690 = 3'h4 == state ? valid_1_23 : _GEN_9662; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10691 = 3'h4 == state ? valid_1_24 : _GEN_9663; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10692 = 3'h4 == state ? valid_1_25 : _GEN_9664; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10693 = 3'h4 == state ? valid_1_26 : _GEN_9665; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10694 = 3'h4 == state ? valid_1_27 : _GEN_9666; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10695 = 3'h4 == state ? valid_1_28 : _GEN_9667; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10696 = 3'h4 == state ? valid_1_29 : _GEN_9668; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10697 = 3'h4 == state ? valid_1_30 : _GEN_9669; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10698 = 3'h4 == state ? valid_1_31 : _GEN_9670; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10699 = 3'h4 == state ? valid_1_32 : _GEN_9671; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10700 = 3'h4 == state ? valid_1_33 : _GEN_9672; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10701 = 3'h4 == state ? valid_1_34 : _GEN_9673; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10702 = 3'h4 == state ? valid_1_35 : _GEN_9674; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10703 = 3'h4 == state ? valid_1_36 : _GEN_9675; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10704 = 3'h4 == state ? valid_1_37 : _GEN_9676; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10705 = 3'h4 == state ? valid_1_38 : _GEN_9677; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10706 = 3'h4 == state ? valid_1_39 : _GEN_9678; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10707 = 3'h4 == state ? valid_1_40 : _GEN_9679; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10708 = 3'h4 == state ? valid_1_41 : _GEN_9680; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10709 = 3'h4 == state ? valid_1_42 : _GEN_9681; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10710 = 3'h4 == state ? valid_1_43 : _GEN_9682; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10711 = 3'h4 == state ? valid_1_44 : _GEN_9683; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10712 = 3'h4 == state ? valid_1_45 : _GEN_9684; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10713 = 3'h4 == state ? valid_1_46 : _GEN_9685; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10714 = 3'h4 == state ? valid_1_47 : _GEN_9686; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10715 = 3'h4 == state ? valid_1_48 : _GEN_9687; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10716 = 3'h4 == state ? valid_1_49 : _GEN_9688; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10717 = 3'h4 == state ? valid_1_50 : _GEN_9689; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10718 = 3'h4 == state ? valid_1_51 : _GEN_9690; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10719 = 3'h4 == state ? valid_1_52 : _GEN_9691; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10720 = 3'h4 == state ? valid_1_53 : _GEN_9692; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10721 = 3'h4 == state ? valid_1_54 : _GEN_9693; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10722 = 3'h4 == state ? valid_1_55 : _GEN_9694; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10723 = 3'h4 == state ? valid_1_56 : _GEN_9695; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10724 = 3'h4 == state ? valid_1_57 : _GEN_9696; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10725 = 3'h4 == state ? valid_1_58 : _GEN_9697; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10726 = 3'h4 == state ? valid_1_59 : _GEN_9698; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10727 = 3'h4 == state ? valid_1_60 : _GEN_9699; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10728 = 3'h4 == state ? valid_1_61 : _GEN_9700; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10729 = 3'h4 == state ? valid_1_62 : _GEN_9701; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10730 = 3'h4 == state ? valid_1_63 : _GEN_9702; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10731 = 3'h4 == state ? valid_1_64 : _GEN_9703; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10732 = 3'h4 == state ? valid_1_65 : _GEN_9704; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10733 = 3'h4 == state ? valid_1_66 : _GEN_9705; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10734 = 3'h4 == state ? valid_1_67 : _GEN_9706; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10735 = 3'h4 == state ? valid_1_68 : _GEN_9707; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10736 = 3'h4 == state ? valid_1_69 : _GEN_9708; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10737 = 3'h4 == state ? valid_1_70 : _GEN_9709; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10738 = 3'h4 == state ? valid_1_71 : _GEN_9710; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10739 = 3'h4 == state ? valid_1_72 : _GEN_9711; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10740 = 3'h4 == state ? valid_1_73 : _GEN_9712; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10741 = 3'h4 == state ? valid_1_74 : _GEN_9713; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10742 = 3'h4 == state ? valid_1_75 : _GEN_9714; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10743 = 3'h4 == state ? valid_1_76 : _GEN_9715; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10744 = 3'h4 == state ? valid_1_77 : _GEN_9716; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10745 = 3'h4 == state ? valid_1_78 : _GEN_9717; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10746 = 3'h4 == state ? valid_1_79 : _GEN_9718; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10747 = 3'h4 == state ? valid_1_80 : _GEN_9719; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10748 = 3'h4 == state ? valid_1_81 : _GEN_9720; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10749 = 3'h4 == state ? valid_1_82 : _GEN_9721; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10750 = 3'h4 == state ? valid_1_83 : _GEN_9722; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10751 = 3'h4 == state ? valid_1_84 : _GEN_9723; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10752 = 3'h4 == state ? valid_1_85 : _GEN_9724; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10753 = 3'h4 == state ? valid_1_86 : _GEN_9725; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10754 = 3'h4 == state ? valid_1_87 : _GEN_9726; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10755 = 3'h4 == state ? valid_1_88 : _GEN_9727; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10756 = 3'h4 == state ? valid_1_89 : _GEN_9728; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10757 = 3'h4 == state ? valid_1_90 : _GEN_9729; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10758 = 3'h4 == state ? valid_1_91 : _GEN_9730; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10759 = 3'h4 == state ? valid_1_92 : _GEN_9731; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10760 = 3'h4 == state ? valid_1_93 : _GEN_9732; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10761 = 3'h4 == state ? valid_1_94 : _GEN_9733; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10762 = 3'h4 == state ? valid_1_95 : _GEN_9734; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10763 = 3'h4 == state ? valid_1_96 : _GEN_9735; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10764 = 3'h4 == state ? valid_1_97 : _GEN_9736; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10765 = 3'h4 == state ? valid_1_98 : _GEN_9737; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10766 = 3'h4 == state ? valid_1_99 : _GEN_9738; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10767 = 3'h4 == state ? valid_1_100 : _GEN_9739; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10768 = 3'h4 == state ? valid_1_101 : _GEN_9740; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10769 = 3'h4 == state ? valid_1_102 : _GEN_9741; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10770 = 3'h4 == state ? valid_1_103 : _GEN_9742; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10771 = 3'h4 == state ? valid_1_104 : _GEN_9743; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10772 = 3'h4 == state ? valid_1_105 : _GEN_9744; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10773 = 3'h4 == state ? valid_1_106 : _GEN_9745; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10774 = 3'h4 == state ? valid_1_107 : _GEN_9746; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10775 = 3'h4 == state ? valid_1_108 : _GEN_9747; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10776 = 3'h4 == state ? valid_1_109 : _GEN_9748; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10777 = 3'h4 == state ? valid_1_110 : _GEN_9749; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10778 = 3'h4 == state ? valid_1_111 : _GEN_9750; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10779 = 3'h4 == state ? valid_1_112 : _GEN_9751; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10780 = 3'h4 == state ? valid_1_113 : _GEN_9752; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10781 = 3'h4 == state ? valid_1_114 : _GEN_9753; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10782 = 3'h4 == state ? valid_1_115 : _GEN_9754; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10783 = 3'h4 == state ? valid_1_116 : _GEN_9755; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10784 = 3'h4 == state ? valid_1_117 : _GEN_9756; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10785 = 3'h4 == state ? valid_1_118 : _GEN_9757; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10786 = 3'h4 == state ? valid_1_119 : _GEN_9758; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10787 = 3'h4 == state ? valid_1_120 : _GEN_9759; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10788 = 3'h4 == state ? valid_1_121 : _GEN_9760; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10789 = 3'h4 == state ? valid_1_122 : _GEN_9761; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10790 = 3'h4 == state ? valid_1_123 : _GEN_9762; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10791 = 3'h4 == state ? valid_1_124 : _GEN_9763; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10792 = 3'h4 == state ? valid_1_125 : _GEN_9764; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10793 = 3'h4 == state ? valid_1_126 : _GEN_9765; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_10794 = 3'h4 == state ? valid_1_127 : _GEN_9766; // @[d_cache.scala 64:18 23:26]
  wire [63:0] _GEN_10795 = 3'h4 == state ? write_back_data : _GEN_9767; // @[d_cache.scala 64:18 29:34]
  wire [38:0] _GEN_10796 = 3'h4 == state ? {{7'd0}, write_back_addr} : _GEN_9768; // @[d_cache.scala 64:18 30:34]
  wire  _GEN_10797 = 3'h4 == state ? dirty_0_0 : _GEN_9769; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10798 = 3'h4 == state ? dirty_0_1 : _GEN_9770; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10799 = 3'h4 == state ? dirty_0_2 : _GEN_9771; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10800 = 3'h4 == state ? dirty_0_3 : _GEN_9772; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10801 = 3'h4 == state ? dirty_0_4 : _GEN_9773; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10802 = 3'h4 == state ? dirty_0_5 : _GEN_9774; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10803 = 3'h4 == state ? dirty_0_6 : _GEN_9775; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10804 = 3'h4 == state ? dirty_0_7 : _GEN_9776; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10805 = 3'h4 == state ? dirty_0_8 : _GEN_9777; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10806 = 3'h4 == state ? dirty_0_9 : _GEN_9778; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10807 = 3'h4 == state ? dirty_0_10 : _GEN_9779; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10808 = 3'h4 == state ? dirty_0_11 : _GEN_9780; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10809 = 3'h4 == state ? dirty_0_12 : _GEN_9781; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10810 = 3'h4 == state ? dirty_0_13 : _GEN_9782; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10811 = 3'h4 == state ? dirty_0_14 : _GEN_9783; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10812 = 3'h4 == state ? dirty_0_15 : _GEN_9784; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10813 = 3'h4 == state ? dirty_0_16 : _GEN_9785; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10814 = 3'h4 == state ? dirty_0_17 : _GEN_9786; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10815 = 3'h4 == state ? dirty_0_18 : _GEN_9787; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10816 = 3'h4 == state ? dirty_0_19 : _GEN_9788; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10817 = 3'h4 == state ? dirty_0_20 : _GEN_9789; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10818 = 3'h4 == state ? dirty_0_21 : _GEN_9790; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10819 = 3'h4 == state ? dirty_0_22 : _GEN_9791; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10820 = 3'h4 == state ? dirty_0_23 : _GEN_9792; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10821 = 3'h4 == state ? dirty_0_24 : _GEN_9793; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10822 = 3'h4 == state ? dirty_0_25 : _GEN_9794; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10823 = 3'h4 == state ? dirty_0_26 : _GEN_9795; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10824 = 3'h4 == state ? dirty_0_27 : _GEN_9796; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10825 = 3'h4 == state ? dirty_0_28 : _GEN_9797; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10826 = 3'h4 == state ? dirty_0_29 : _GEN_9798; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10827 = 3'h4 == state ? dirty_0_30 : _GEN_9799; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10828 = 3'h4 == state ? dirty_0_31 : _GEN_9800; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10829 = 3'h4 == state ? dirty_0_32 : _GEN_9801; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10830 = 3'h4 == state ? dirty_0_33 : _GEN_9802; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10831 = 3'h4 == state ? dirty_0_34 : _GEN_9803; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10832 = 3'h4 == state ? dirty_0_35 : _GEN_9804; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10833 = 3'h4 == state ? dirty_0_36 : _GEN_9805; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10834 = 3'h4 == state ? dirty_0_37 : _GEN_9806; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10835 = 3'h4 == state ? dirty_0_38 : _GEN_9807; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10836 = 3'h4 == state ? dirty_0_39 : _GEN_9808; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10837 = 3'h4 == state ? dirty_0_40 : _GEN_9809; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10838 = 3'h4 == state ? dirty_0_41 : _GEN_9810; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10839 = 3'h4 == state ? dirty_0_42 : _GEN_9811; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10840 = 3'h4 == state ? dirty_0_43 : _GEN_9812; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10841 = 3'h4 == state ? dirty_0_44 : _GEN_9813; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10842 = 3'h4 == state ? dirty_0_45 : _GEN_9814; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10843 = 3'h4 == state ? dirty_0_46 : _GEN_9815; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10844 = 3'h4 == state ? dirty_0_47 : _GEN_9816; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10845 = 3'h4 == state ? dirty_0_48 : _GEN_9817; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10846 = 3'h4 == state ? dirty_0_49 : _GEN_9818; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10847 = 3'h4 == state ? dirty_0_50 : _GEN_9819; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10848 = 3'h4 == state ? dirty_0_51 : _GEN_9820; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10849 = 3'h4 == state ? dirty_0_52 : _GEN_9821; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10850 = 3'h4 == state ? dirty_0_53 : _GEN_9822; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10851 = 3'h4 == state ? dirty_0_54 : _GEN_9823; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10852 = 3'h4 == state ? dirty_0_55 : _GEN_9824; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10853 = 3'h4 == state ? dirty_0_56 : _GEN_9825; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10854 = 3'h4 == state ? dirty_0_57 : _GEN_9826; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10855 = 3'h4 == state ? dirty_0_58 : _GEN_9827; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10856 = 3'h4 == state ? dirty_0_59 : _GEN_9828; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10857 = 3'h4 == state ? dirty_0_60 : _GEN_9829; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10858 = 3'h4 == state ? dirty_0_61 : _GEN_9830; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10859 = 3'h4 == state ? dirty_0_62 : _GEN_9831; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10860 = 3'h4 == state ? dirty_0_63 : _GEN_9832; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10861 = 3'h4 == state ? dirty_0_64 : _GEN_9833; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10862 = 3'h4 == state ? dirty_0_65 : _GEN_9834; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10863 = 3'h4 == state ? dirty_0_66 : _GEN_9835; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10864 = 3'h4 == state ? dirty_0_67 : _GEN_9836; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10865 = 3'h4 == state ? dirty_0_68 : _GEN_9837; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10866 = 3'h4 == state ? dirty_0_69 : _GEN_9838; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10867 = 3'h4 == state ? dirty_0_70 : _GEN_9839; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10868 = 3'h4 == state ? dirty_0_71 : _GEN_9840; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10869 = 3'h4 == state ? dirty_0_72 : _GEN_9841; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10870 = 3'h4 == state ? dirty_0_73 : _GEN_9842; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10871 = 3'h4 == state ? dirty_0_74 : _GEN_9843; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10872 = 3'h4 == state ? dirty_0_75 : _GEN_9844; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10873 = 3'h4 == state ? dirty_0_76 : _GEN_9845; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10874 = 3'h4 == state ? dirty_0_77 : _GEN_9846; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10875 = 3'h4 == state ? dirty_0_78 : _GEN_9847; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10876 = 3'h4 == state ? dirty_0_79 : _GEN_9848; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10877 = 3'h4 == state ? dirty_0_80 : _GEN_9849; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10878 = 3'h4 == state ? dirty_0_81 : _GEN_9850; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10879 = 3'h4 == state ? dirty_0_82 : _GEN_9851; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10880 = 3'h4 == state ? dirty_0_83 : _GEN_9852; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10881 = 3'h4 == state ? dirty_0_84 : _GEN_9853; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10882 = 3'h4 == state ? dirty_0_85 : _GEN_9854; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10883 = 3'h4 == state ? dirty_0_86 : _GEN_9855; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10884 = 3'h4 == state ? dirty_0_87 : _GEN_9856; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10885 = 3'h4 == state ? dirty_0_88 : _GEN_9857; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10886 = 3'h4 == state ? dirty_0_89 : _GEN_9858; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10887 = 3'h4 == state ? dirty_0_90 : _GEN_9859; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10888 = 3'h4 == state ? dirty_0_91 : _GEN_9860; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10889 = 3'h4 == state ? dirty_0_92 : _GEN_9861; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10890 = 3'h4 == state ? dirty_0_93 : _GEN_9862; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10891 = 3'h4 == state ? dirty_0_94 : _GEN_9863; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10892 = 3'h4 == state ? dirty_0_95 : _GEN_9864; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10893 = 3'h4 == state ? dirty_0_96 : _GEN_9865; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10894 = 3'h4 == state ? dirty_0_97 : _GEN_9866; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10895 = 3'h4 == state ? dirty_0_98 : _GEN_9867; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10896 = 3'h4 == state ? dirty_0_99 : _GEN_9868; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10897 = 3'h4 == state ? dirty_0_100 : _GEN_9869; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10898 = 3'h4 == state ? dirty_0_101 : _GEN_9870; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10899 = 3'h4 == state ? dirty_0_102 : _GEN_9871; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10900 = 3'h4 == state ? dirty_0_103 : _GEN_9872; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10901 = 3'h4 == state ? dirty_0_104 : _GEN_9873; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10902 = 3'h4 == state ? dirty_0_105 : _GEN_9874; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10903 = 3'h4 == state ? dirty_0_106 : _GEN_9875; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10904 = 3'h4 == state ? dirty_0_107 : _GEN_9876; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10905 = 3'h4 == state ? dirty_0_108 : _GEN_9877; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10906 = 3'h4 == state ? dirty_0_109 : _GEN_9878; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10907 = 3'h4 == state ? dirty_0_110 : _GEN_9879; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10908 = 3'h4 == state ? dirty_0_111 : _GEN_9880; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10909 = 3'h4 == state ? dirty_0_112 : _GEN_9881; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10910 = 3'h4 == state ? dirty_0_113 : _GEN_9882; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10911 = 3'h4 == state ? dirty_0_114 : _GEN_9883; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10912 = 3'h4 == state ? dirty_0_115 : _GEN_9884; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10913 = 3'h4 == state ? dirty_0_116 : _GEN_9885; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10914 = 3'h4 == state ? dirty_0_117 : _GEN_9886; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10915 = 3'h4 == state ? dirty_0_118 : _GEN_9887; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10916 = 3'h4 == state ? dirty_0_119 : _GEN_9888; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10917 = 3'h4 == state ? dirty_0_120 : _GEN_9889; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10918 = 3'h4 == state ? dirty_0_121 : _GEN_9890; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10919 = 3'h4 == state ? dirty_0_122 : _GEN_9891; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10920 = 3'h4 == state ? dirty_0_123 : _GEN_9892; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10921 = 3'h4 == state ? dirty_0_124 : _GEN_9893; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10922 = 3'h4 == state ? dirty_0_125 : _GEN_9894; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10923 = 3'h4 == state ? dirty_0_126 : _GEN_9895; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10924 = 3'h4 == state ? dirty_0_127 : _GEN_9896; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_10925 = 3'h4 == state ? dirty_1_0 : _GEN_9897; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10926 = 3'h4 == state ? dirty_1_1 : _GEN_9898; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10927 = 3'h4 == state ? dirty_1_2 : _GEN_9899; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10928 = 3'h4 == state ? dirty_1_3 : _GEN_9900; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10929 = 3'h4 == state ? dirty_1_4 : _GEN_9901; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10930 = 3'h4 == state ? dirty_1_5 : _GEN_9902; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10931 = 3'h4 == state ? dirty_1_6 : _GEN_9903; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10932 = 3'h4 == state ? dirty_1_7 : _GEN_9904; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10933 = 3'h4 == state ? dirty_1_8 : _GEN_9905; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10934 = 3'h4 == state ? dirty_1_9 : _GEN_9906; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10935 = 3'h4 == state ? dirty_1_10 : _GEN_9907; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10936 = 3'h4 == state ? dirty_1_11 : _GEN_9908; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10937 = 3'h4 == state ? dirty_1_12 : _GEN_9909; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10938 = 3'h4 == state ? dirty_1_13 : _GEN_9910; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10939 = 3'h4 == state ? dirty_1_14 : _GEN_9911; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10940 = 3'h4 == state ? dirty_1_15 : _GEN_9912; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10941 = 3'h4 == state ? dirty_1_16 : _GEN_9913; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10942 = 3'h4 == state ? dirty_1_17 : _GEN_9914; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10943 = 3'h4 == state ? dirty_1_18 : _GEN_9915; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10944 = 3'h4 == state ? dirty_1_19 : _GEN_9916; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10945 = 3'h4 == state ? dirty_1_20 : _GEN_9917; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10946 = 3'h4 == state ? dirty_1_21 : _GEN_9918; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10947 = 3'h4 == state ? dirty_1_22 : _GEN_9919; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10948 = 3'h4 == state ? dirty_1_23 : _GEN_9920; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10949 = 3'h4 == state ? dirty_1_24 : _GEN_9921; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10950 = 3'h4 == state ? dirty_1_25 : _GEN_9922; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10951 = 3'h4 == state ? dirty_1_26 : _GEN_9923; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10952 = 3'h4 == state ? dirty_1_27 : _GEN_9924; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10953 = 3'h4 == state ? dirty_1_28 : _GEN_9925; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10954 = 3'h4 == state ? dirty_1_29 : _GEN_9926; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10955 = 3'h4 == state ? dirty_1_30 : _GEN_9927; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10956 = 3'h4 == state ? dirty_1_31 : _GEN_9928; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10957 = 3'h4 == state ? dirty_1_32 : _GEN_9929; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10958 = 3'h4 == state ? dirty_1_33 : _GEN_9930; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10959 = 3'h4 == state ? dirty_1_34 : _GEN_9931; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10960 = 3'h4 == state ? dirty_1_35 : _GEN_9932; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10961 = 3'h4 == state ? dirty_1_36 : _GEN_9933; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10962 = 3'h4 == state ? dirty_1_37 : _GEN_9934; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10963 = 3'h4 == state ? dirty_1_38 : _GEN_9935; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10964 = 3'h4 == state ? dirty_1_39 : _GEN_9936; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10965 = 3'h4 == state ? dirty_1_40 : _GEN_9937; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10966 = 3'h4 == state ? dirty_1_41 : _GEN_9938; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10967 = 3'h4 == state ? dirty_1_42 : _GEN_9939; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10968 = 3'h4 == state ? dirty_1_43 : _GEN_9940; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10969 = 3'h4 == state ? dirty_1_44 : _GEN_9941; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10970 = 3'h4 == state ? dirty_1_45 : _GEN_9942; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10971 = 3'h4 == state ? dirty_1_46 : _GEN_9943; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10972 = 3'h4 == state ? dirty_1_47 : _GEN_9944; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10973 = 3'h4 == state ? dirty_1_48 : _GEN_9945; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10974 = 3'h4 == state ? dirty_1_49 : _GEN_9946; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10975 = 3'h4 == state ? dirty_1_50 : _GEN_9947; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10976 = 3'h4 == state ? dirty_1_51 : _GEN_9948; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10977 = 3'h4 == state ? dirty_1_52 : _GEN_9949; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10978 = 3'h4 == state ? dirty_1_53 : _GEN_9950; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10979 = 3'h4 == state ? dirty_1_54 : _GEN_9951; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10980 = 3'h4 == state ? dirty_1_55 : _GEN_9952; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10981 = 3'h4 == state ? dirty_1_56 : _GEN_9953; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10982 = 3'h4 == state ? dirty_1_57 : _GEN_9954; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10983 = 3'h4 == state ? dirty_1_58 : _GEN_9955; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10984 = 3'h4 == state ? dirty_1_59 : _GEN_9956; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10985 = 3'h4 == state ? dirty_1_60 : _GEN_9957; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10986 = 3'h4 == state ? dirty_1_61 : _GEN_9958; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10987 = 3'h4 == state ? dirty_1_62 : _GEN_9959; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10988 = 3'h4 == state ? dirty_1_63 : _GEN_9960; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10989 = 3'h4 == state ? dirty_1_64 : _GEN_9961; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10990 = 3'h4 == state ? dirty_1_65 : _GEN_9962; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10991 = 3'h4 == state ? dirty_1_66 : _GEN_9963; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10992 = 3'h4 == state ? dirty_1_67 : _GEN_9964; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10993 = 3'h4 == state ? dirty_1_68 : _GEN_9965; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10994 = 3'h4 == state ? dirty_1_69 : _GEN_9966; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10995 = 3'h4 == state ? dirty_1_70 : _GEN_9967; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10996 = 3'h4 == state ? dirty_1_71 : _GEN_9968; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10997 = 3'h4 == state ? dirty_1_72 : _GEN_9969; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10998 = 3'h4 == state ? dirty_1_73 : _GEN_9970; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_10999 = 3'h4 == state ? dirty_1_74 : _GEN_9971; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11000 = 3'h4 == state ? dirty_1_75 : _GEN_9972; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11001 = 3'h4 == state ? dirty_1_76 : _GEN_9973; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11002 = 3'h4 == state ? dirty_1_77 : _GEN_9974; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11003 = 3'h4 == state ? dirty_1_78 : _GEN_9975; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11004 = 3'h4 == state ? dirty_1_79 : _GEN_9976; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11005 = 3'h4 == state ? dirty_1_80 : _GEN_9977; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11006 = 3'h4 == state ? dirty_1_81 : _GEN_9978; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11007 = 3'h4 == state ? dirty_1_82 : _GEN_9979; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11008 = 3'h4 == state ? dirty_1_83 : _GEN_9980; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11009 = 3'h4 == state ? dirty_1_84 : _GEN_9981; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11010 = 3'h4 == state ? dirty_1_85 : _GEN_9982; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11011 = 3'h4 == state ? dirty_1_86 : _GEN_9983; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11012 = 3'h4 == state ? dirty_1_87 : _GEN_9984; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11013 = 3'h4 == state ? dirty_1_88 : _GEN_9985; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11014 = 3'h4 == state ? dirty_1_89 : _GEN_9986; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11015 = 3'h4 == state ? dirty_1_90 : _GEN_9987; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11016 = 3'h4 == state ? dirty_1_91 : _GEN_9988; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11017 = 3'h4 == state ? dirty_1_92 : _GEN_9989; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11018 = 3'h4 == state ? dirty_1_93 : _GEN_9990; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11019 = 3'h4 == state ? dirty_1_94 : _GEN_9991; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11020 = 3'h4 == state ? dirty_1_95 : _GEN_9992; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11021 = 3'h4 == state ? dirty_1_96 : _GEN_9993; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11022 = 3'h4 == state ? dirty_1_97 : _GEN_9994; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11023 = 3'h4 == state ? dirty_1_98 : _GEN_9995; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11024 = 3'h4 == state ? dirty_1_99 : _GEN_9996; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11025 = 3'h4 == state ? dirty_1_100 : _GEN_9997; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11026 = 3'h4 == state ? dirty_1_101 : _GEN_9998; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11027 = 3'h4 == state ? dirty_1_102 : _GEN_9999; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11028 = 3'h4 == state ? dirty_1_103 : _GEN_10000; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11029 = 3'h4 == state ? dirty_1_104 : _GEN_10001; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11030 = 3'h4 == state ? dirty_1_105 : _GEN_10002; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11031 = 3'h4 == state ? dirty_1_106 : _GEN_10003; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11032 = 3'h4 == state ? dirty_1_107 : _GEN_10004; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11033 = 3'h4 == state ? dirty_1_108 : _GEN_10005; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11034 = 3'h4 == state ? dirty_1_109 : _GEN_10006; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11035 = 3'h4 == state ? dirty_1_110 : _GEN_10007; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11036 = 3'h4 == state ? dirty_1_111 : _GEN_10008; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11037 = 3'h4 == state ? dirty_1_112 : _GEN_10009; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11038 = 3'h4 == state ? dirty_1_113 : _GEN_10010; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11039 = 3'h4 == state ? dirty_1_114 : _GEN_10011; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11040 = 3'h4 == state ? dirty_1_115 : _GEN_10012; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11041 = 3'h4 == state ? dirty_1_116 : _GEN_10013; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11042 = 3'h4 == state ? dirty_1_117 : _GEN_10014; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11043 = 3'h4 == state ? dirty_1_118 : _GEN_10015; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11044 = 3'h4 == state ? dirty_1_119 : _GEN_10016; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11045 = 3'h4 == state ? dirty_1_120 : _GEN_10017; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11046 = 3'h4 == state ? dirty_1_121 : _GEN_10018; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11047 = 3'h4 == state ? dirty_1_122 : _GEN_10019; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11048 = 3'h4 == state ? dirty_1_123 : _GEN_10020; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11049 = 3'h4 == state ? dirty_1_124 : _GEN_10021; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11050 = 3'h4 == state ? dirty_1_125 : _GEN_10022; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11051 = 3'h4 == state ? dirty_1_126 : _GEN_10023; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11052 = 3'h4 == state ? dirty_1_127 : _GEN_10024; // @[d_cache.scala 64:18 25:26]
  wire [2:0] _GEN_11053 = 3'h3 == state ? _GEN_2059 : _GEN_10025; // @[d_cache.scala 64:18]
  wire [63:0] _GEN_11054 = 3'h3 == state ? _GEN_2060 : receive_data; // @[d_cache.scala 64:18 34:31]
  wire [63:0] _GEN_11055 = 3'h3 == state ? ram_0_0 : _GEN_10026; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11056 = 3'h3 == state ? ram_0_1 : _GEN_10027; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11057 = 3'h3 == state ? ram_0_2 : _GEN_10028; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11058 = 3'h3 == state ? ram_0_3 : _GEN_10029; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11059 = 3'h3 == state ? ram_0_4 : _GEN_10030; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11060 = 3'h3 == state ? ram_0_5 : _GEN_10031; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11061 = 3'h3 == state ? ram_0_6 : _GEN_10032; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11062 = 3'h3 == state ? ram_0_7 : _GEN_10033; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11063 = 3'h3 == state ? ram_0_8 : _GEN_10034; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11064 = 3'h3 == state ? ram_0_9 : _GEN_10035; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11065 = 3'h3 == state ? ram_0_10 : _GEN_10036; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11066 = 3'h3 == state ? ram_0_11 : _GEN_10037; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11067 = 3'h3 == state ? ram_0_12 : _GEN_10038; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11068 = 3'h3 == state ? ram_0_13 : _GEN_10039; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11069 = 3'h3 == state ? ram_0_14 : _GEN_10040; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11070 = 3'h3 == state ? ram_0_15 : _GEN_10041; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11071 = 3'h3 == state ? ram_0_16 : _GEN_10042; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11072 = 3'h3 == state ? ram_0_17 : _GEN_10043; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11073 = 3'h3 == state ? ram_0_18 : _GEN_10044; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11074 = 3'h3 == state ? ram_0_19 : _GEN_10045; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11075 = 3'h3 == state ? ram_0_20 : _GEN_10046; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11076 = 3'h3 == state ? ram_0_21 : _GEN_10047; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11077 = 3'h3 == state ? ram_0_22 : _GEN_10048; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11078 = 3'h3 == state ? ram_0_23 : _GEN_10049; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11079 = 3'h3 == state ? ram_0_24 : _GEN_10050; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11080 = 3'h3 == state ? ram_0_25 : _GEN_10051; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11081 = 3'h3 == state ? ram_0_26 : _GEN_10052; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11082 = 3'h3 == state ? ram_0_27 : _GEN_10053; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11083 = 3'h3 == state ? ram_0_28 : _GEN_10054; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11084 = 3'h3 == state ? ram_0_29 : _GEN_10055; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11085 = 3'h3 == state ? ram_0_30 : _GEN_10056; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11086 = 3'h3 == state ? ram_0_31 : _GEN_10057; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11087 = 3'h3 == state ? ram_0_32 : _GEN_10058; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11088 = 3'h3 == state ? ram_0_33 : _GEN_10059; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11089 = 3'h3 == state ? ram_0_34 : _GEN_10060; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11090 = 3'h3 == state ? ram_0_35 : _GEN_10061; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11091 = 3'h3 == state ? ram_0_36 : _GEN_10062; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11092 = 3'h3 == state ? ram_0_37 : _GEN_10063; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11093 = 3'h3 == state ? ram_0_38 : _GEN_10064; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11094 = 3'h3 == state ? ram_0_39 : _GEN_10065; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11095 = 3'h3 == state ? ram_0_40 : _GEN_10066; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11096 = 3'h3 == state ? ram_0_41 : _GEN_10067; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11097 = 3'h3 == state ? ram_0_42 : _GEN_10068; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11098 = 3'h3 == state ? ram_0_43 : _GEN_10069; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11099 = 3'h3 == state ? ram_0_44 : _GEN_10070; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11100 = 3'h3 == state ? ram_0_45 : _GEN_10071; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11101 = 3'h3 == state ? ram_0_46 : _GEN_10072; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11102 = 3'h3 == state ? ram_0_47 : _GEN_10073; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11103 = 3'h3 == state ? ram_0_48 : _GEN_10074; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11104 = 3'h3 == state ? ram_0_49 : _GEN_10075; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11105 = 3'h3 == state ? ram_0_50 : _GEN_10076; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11106 = 3'h3 == state ? ram_0_51 : _GEN_10077; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11107 = 3'h3 == state ? ram_0_52 : _GEN_10078; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11108 = 3'h3 == state ? ram_0_53 : _GEN_10079; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11109 = 3'h3 == state ? ram_0_54 : _GEN_10080; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11110 = 3'h3 == state ? ram_0_55 : _GEN_10081; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11111 = 3'h3 == state ? ram_0_56 : _GEN_10082; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11112 = 3'h3 == state ? ram_0_57 : _GEN_10083; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11113 = 3'h3 == state ? ram_0_58 : _GEN_10084; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11114 = 3'h3 == state ? ram_0_59 : _GEN_10085; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11115 = 3'h3 == state ? ram_0_60 : _GEN_10086; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11116 = 3'h3 == state ? ram_0_61 : _GEN_10087; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11117 = 3'h3 == state ? ram_0_62 : _GEN_10088; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11118 = 3'h3 == state ? ram_0_63 : _GEN_10089; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11119 = 3'h3 == state ? ram_0_64 : _GEN_10090; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11120 = 3'h3 == state ? ram_0_65 : _GEN_10091; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11121 = 3'h3 == state ? ram_0_66 : _GEN_10092; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11122 = 3'h3 == state ? ram_0_67 : _GEN_10093; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11123 = 3'h3 == state ? ram_0_68 : _GEN_10094; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11124 = 3'h3 == state ? ram_0_69 : _GEN_10095; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11125 = 3'h3 == state ? ram_0_70 : _GEN_10096; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11126 = 3'h3 == state ? ram_0_71 : _GEN_10097; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11127 = 3'h3 == state ? ram_0_72 : _GEN_10098; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11128 = 3'h3 == state ? ram_0_73 : _GEN_10099; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11129 = 3'h3 == state ? ram_0_74 : _GEN_10100; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11130 = 3'h3 == state ? ram_0_75 : _GEN_10101; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11131 = 3'h3 == state ? ram_0_76 : _GEN_10102; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11132 = 3'h3 == state ? ram_0_77 : _GEN_10103; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11133 = 3'h3 == state ? ram_0_78 : _GEN_10104; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11134 = 3'h3 == state ? ram_0_79 : _GEN_10105; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11135 = 3'h3 == state ? ram_0_80 : _GEN_10106; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11136 = 3'h3 == state ? ram_0_81 : _GEN_10107; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11137 = 3'h3 == state ? ram_0_82 : _GEN_10108; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11138 = 3'h3 == state ? ram_0_83 : _GEN_10109; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11139 = 3'h3 == state ? ram_0_84 : _GEN_10110; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11140 = 3'h3 == state ? ram_0_85 : _GEN_10111; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11141 = 3'h3 == state ? ram_0_86 : _GEN_10112; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11142 = 3'h3 == state ? ram_0_87 : _GEN_10113; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11143 = 3'h3 == state ? ram_0_88 : _GEN_10114; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11144 = 3'h3 == state ? ram_0_89 : _GEN_10115; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11145 = 3'h3 == state ? ram_0_90 : _GEN_10116; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11146 = 3'h3 == state ? ram_0_91 : _GEN_10117; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11147 = 3'h3 == state ? ram_0_92 : _GEN_10118; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11148 = 3'h3 == state ? ram_0_93 : _GEN_10119; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11149 = 3'h3 == state ? ram_0_94 : _GEN_10120; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11150 = 3'h3 == state ? ram_0_95 : _GEN_10121; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11151 = 3'h3 == state ? ram_0_96 : _GEN_10122; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11152 = 3'h3 == state ? ram_0_97 : _GEN_10123; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11153 = 3'h3 == state ? ram_0_98 : _GEN_10124; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11154 = 3'h3 == state ? ram_0_99 : _GEN_10125; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11155 = 3'h3 == state ? ram_0_100 : _GEN_10126; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11156 = 3'h3 == state ? ram_0_101 : _GEN_10127; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11157 = 3'h3 == state ? ram_0_102 : _GEN_10128; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11158 = 3'h3 == state ? ram_0_103 : _GEN_10129; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11159 = 3'h3 == state ? ram_0_104 : _GEN_10130; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11160 = 3'h3 == state ? ram_0_105 : _GEN_10131; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11161 = 3'h3 == state ? ram_0_106 : _GEN_10132; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11162 = 3'h3 == state ? ram_0_107 : _GEN_10133; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11163 = 3'h3 == state ? ram_0_108 : _GEN_10134; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11164 = 3'h3 == state ? ram_0_109 : _GEN_10135; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11165 = 3'h3 == state ? ram_0_110 : _GEN_10136; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11166 = 3'h3 == state ? ram_0_111 : _GEN_10137; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11167 = 3'h3 == state ? ram_0_112 : _GEN_10138; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11168 = 3'h3 == state ? ram_0_113 : _GEN_10139; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11169 = 3'h3 == state ? ram_0_114 : _GEN_10140; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11170 = 3'h3 == state ? ram_0_115 : _GEN_10141; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11171 = 3'h3 == state ? ram_0_116 : _GEN_10142; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11172 = 3'h3 == state ? ram_0_117 : _GEN_10143; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11173 = 3'h3 == state ? ram_0_118 : _GEN_10144; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11174 = 3'h3 == state ? ram_0_119 : _GEN_10145; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11175 = 3'h3 == state ? ram_0_120 : _GEN_10146; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11176 = 3'h3 == state ? ram_0_121 : _GEN_10147; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11177 = 3'h3 == state ? ram_0_122 : _GEN_10148; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11178 = 3'h3 == state ? ram_0_123 : _GEN_10149; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11179 = 3'h3 == state ? ram_0_124 : _GEN_10150; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11180 = 3'h3 == state ? ram_0_125 : _GEN_10151; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11181 = 3'h3 == state ? ram_0_126 : _GEN_10152; // @[d_cache.scala 64:18 18:24]
  wire [63:0] _GEN_11182 = 3'h3 == state ? ram_0_127 : _GEN_10153; // @[d_cache.scala 64:18 18:24]
  wire [31:0] _GEN_11183 = 3'h3 == state ? tag_0_0 : _GEN_10154; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11184 = 3'h3 == state ? tag_0_1 : _GEN_10155; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11185 = 3'h3 == state ? tag_0_2 : _GEN_10156; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11186 = 3'h3 == state ? tag_0_3 : _GEN_10157; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11187 = 3'h3 == state ? tag_0_4 : _GEN_10158; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11188 = 3'h3 == state ? tag_0_5 : _GEN_10159; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11189 = 3'h3 == state ? tag_0_6 : _GEN_10160; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11190 = 3'h3 == state ? tag_0_7 : _GEN_10161; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11191 = 3'h3 == state ? tag_0_8 : _GEN_10162; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11192 = 3'h3 == state ? tag_0_9 : _GEN_10163; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11193 = 3'h3 == state ? tag_0_10 : _GEN_10164; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11194 = 3'h3 == state ? tag_0_11 : _GEN_10165; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11195 = 3'h3 == state ? tag_0_12 : _GEN_10166; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11196 = 3'h3 == state ? tag_0_13 : _GEN_10167; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11197 = 3'h3 == state ? tag_0_14 : _GEN_10168; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11198 = 3'h3 == state ? tag_0_15 : _GEN_10169; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11199 = 3'h3 == state ? tag_0_16 : _GEN_10170; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11200 = 3'h3 == state ? tag_0_17 : _GEN_10171; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11201 = 3'h3 == state ? tag_0_18 : _GEN_10172; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11202 = 3'h3 == state ? tag_0_19 : _GEN_10173; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11203 = 3'h3 == state ? tag_0_20 : _GEN_10174; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11204 = 3'h3 == state ? tag_0_21 : _GEN_10175; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11205 = 3'h3 == state ? tag_0_22 : _GEN_10176; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11206 = 3'h3 == state ? tag_0_23 : _GEN_10177; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11207 = 3'h3 == state ? tag_0_24 : _GEN_10178; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11208 = 3'h3 == state ? tag_0_25 : _GEN_10179; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11209 = 3'h3 == state ? tag_0_26 : _GEN_10180; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11210 = 3'h3 == state ? tag_0_27 : _GEN_10181; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11211 = 3'h3 == state ? tag_0_28 : _GEN_10182; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11212 = 3'h3 == state ? tag_0_29 : _GEN_10183; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11213 = 3'h3 == state ? tag_0_30 : _GEN_10184; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11214 = 3'h3 == state ? tag_0_31 : _GEN_10185; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11215 = 3'h3 == state ? tag_0_32 : _GEN_10186; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11216 = 3'h3 == state ? tag_0_33 : _GEN_10187; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11217 = 3'h3 == state ? tag_0_34 : _GEN_10188; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11218 = 3'h3 == state ? tag_0_35 : _GEN_10189; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11219 = 3'h3 == state ? tag_0_36 : _GEN_10190; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11220 = 3'h3 == state ? tag_0_37 : _GEN_10191; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11221 = 3'h3 == state ? tag_0_38 : _GEN_10192; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11222 = 3'h3 == state ? tag_0_39 : _GEN_10193; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11223 = 3'h3 == state ? tag_0_40 : _GEN_10194; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11224 = 3'h3 == state ? tag_0_41 : _GEN_10195; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11225 = 3'h3 == state ? tag_0_42 : _GEN_10196; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11226 = 3'h3 == state ? tag_0_43 : _GEN_10197; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11227 = 3'h3 == state ? tag_0_44 : _GEN_10198; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11228 = 3'h3 == state ? tag_0_45 : _GEN_10199; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11229 = 3'h3 == state ? tag_0_46 : _GEN_10200; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11230 = 3'h3 == state ? tag_0_47 : _GEN_10201; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11231 = 3'h3 == state ? tag_0_48 : _GEN_10202; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11232 = 3'h3 == state ? tag_0_49 : _GEN_10203; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11233 = 3'h3 == state ? tag_0_50 : _GEN_10204; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11234 = 3'h3 == state ? tag_0_51 : _GEN_10205; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11235 = 3'h3 == state ? tag_0_52 : _GEN_10206; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11236 = 3'h3 == state ? tag_0_53 : _GEN_10207; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11237 = 3'h3 == state ? tag_0_54 : _GEN_10208; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11238 = 3'h3 == state ? tag_0_55 : _GEN_10209; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11239 = 3'h3 == state ? tag_0_56 : _GEN_10210; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11240 = 3'h3 == state ? tag_0_57 : _GEN_10211; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11241 = 3'h3 == state ? tag_0_58 : _GEN_10212; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11242 = 3'h3 == state ? tag_0_59 : _GEN_10213; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11243 = 3'h3 == state ? tag_0_60 : _GEN_10214; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11244 = 3'h3 == state ? tag_0_61 : _GEN_10215; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11245 = 3'h3 == state ? tag_0_62 : _GEN_10216; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11246 = 3'h3 == state ? tag_0_63 : _GEN_10217; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11247 = 3'h3 == state ? tag_0_64 : _GEN_10218; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11248 = 3'h3 == state ? tag_0_65 : _GEN_10219; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11249 = 3'h3 == state ? tag_0_66 : _GEN_10220; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11250 = 3'h3 == state ? tag_0_67 : _GEN_10221; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11251 = 3'h3 == state ? tag_0_68 : _GEN_10222; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11252 = 3'h3 == state ? tag_0_69 : _GEN_10223; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11253 = 3'h3 == state ? tag_0_70 : _GEN_10224; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11254 = 3'h3 == state ? tag_0_71 : _GEN_10225; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11255 = 3'h3 == state ? tag_0_72 : _GEN_10226; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11256 = 3'h3 == state ? tag_0_73 : _GEN_10227; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11257 = 3'h3 == state ? tag_0_74 : _GEN_10228; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11258 = 3'h3 == state ? tag_0_75 : _GEN_10229; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11259 = 3'h3 == state ? tag_0_76 : _GEN_10230; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11260 = 3'h3 == state ? tag_0_77 : _GEN_10231; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11261 = 3'h3 == state ? tag_0_78 : _GEN_10232; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11262 = 3'h3 == state ? tag_0_79 : _GEN_10233; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11263 = 3'h3 == state ? tag_0_80 : _GEN_10234; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11264 = 3'h3 == state ? tag_0_81 : _GEN_10235; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11265 = 3'h3 == state ? tag_0_82 : _GEN_10236; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11266 = 3'h3 == state ? tag_0_83 : _GEN_10237; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11267 = 3'h3 == state ? tag_0_84 : _GEN_10238; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11268 = 3'h3 == state ? tag_0_85 : _GEN_10239; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11269 = 3'h3 == state ? tag_0_86 : _GEN_10240; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11270 = 3'h3 == state ? tag_0_87 : _GEN_10241; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11271 = 3'h3 == state ? tag_0_88 : _GEN_10242; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11272 = 3'h3 == state ? tag_0_89 : _GEN_10243; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11273 = 3'h3 == state ? tag_0_90 : _GEN_10244; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11274 = 3'h3 == state ? tag_0_91 : _GEN_10245; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11275 = 3'h3 == state ? tag_0_92 : _GEN_10246; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11276 = 3'h3 == state ? tag_0_93 : _GEN_10247; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11277 = 3'h3 == state ? tag_0_94 : _GEN_10248; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11278 = 3'h3 == state ? tag_0_95 : _GEN_10249; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11279 = 3'h3 == state ? tag_0_96 : _GEN_10250; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11280 = 3'h3 == state ? tag_0_97 : _GEN_10251; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11281 = 3'h3 == state ? tag_0_98 : _GEN_10252; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11282 = 3'h3 == state ? tag_0_99 : _GEN_10253; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11283 = 3'h3 == state ? tag_0_100 : _GEN_10254; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11284 = 3'h3 == state ? tag_0_101 : _GEN_10255; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11285 = 3'h3 == state ? tag_0_102 : _GEN_10256; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11286 = 3'h3 == state ? tag_0_103 : _GEN_10257; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11287 = 3'h3 == state ? tag_0_104 : _GEN_10258; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11288 = 3'h3 == state ? tag_0_105 : _GEN_10259; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11289 = 3'h3 == state ? tag_0_106 : _GEN_10260; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11290 = 3'h3 == state ? tag_0_107 : _GEN_10261; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11291 = 3'h3 == state ? tag_0_108 : _GEN_10262; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11292 = 3'h3 == state ? tag_0_109 : _GEN_10263; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11293 = 3'h3 == state ? tag_0_110 : _GEN_10264; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11294 = 3'h3 == state ? tag_0_111 : _GEN_10265; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11295 = 3'h3 == state ? tag_0_112 : _GEN_10266; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11296 = 3'h3 == state ? tag_0_113 : _GEN_10267; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11297 = 3'h3 == state ? tag_0_114 : _GEN_10268; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11298 = 3'h3 == state ? tag_0_115 : _GEN_10269; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11299 = 3'h3 == state ? tag_0_116 : _GEN_10270; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11300 = 3'h3 == state ? tag_0_117 : _GEN_10271; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11301 = 3'h3 == state ? tag_0_118 : _GEN_10272; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11302 = 3'h3 == state ? tag_0_119 : _GEN_10273; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11303 = 3'h3 == state ? tag_0_120 : _GEN_10274; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11304 = 3'h3 == state ? tag_0_121 : _GEN_10275; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11305 = 3'h3 == state ? tag_0_122 : _GEN_10276; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11306 = 3'h3 == state ? tag_0_123 : _GEN_10277; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11307 = 3'h3 == state ? tag_0_124 : _GEN_10278; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11308 = 3'h3 == state ? tag_0_125 : _GEN_10279; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11309 = 3'h3 == state ? tag_0_126 : _GEN_10280; // @[d_cache.scala 64:18 20:24]
  wire [31:0] _GEN_11310 = 3'h3 == state ? tag_0_127 : _GEN_10281; // @[d_cache.scala 64:18 20:24]
  wire  _GEN_11311 = 3'h3 == state ? valid_0_0 : _GEN_10282; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11312 = 3'h3 == state ? valid_0_1 : _GEN_10283; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11313 = 3'h3 == state ? valid_0_2 : _GEN_10284; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11314 = 3'h3 == state ? valid_0_3 : _GEN_10285; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11315 = 3'h3 == state ? valid_0_4 : _GEN_10286; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11316 = 3'h3 == state ? valid_0_5 : _GEN_10287; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11317 = 3'h3 == state ? valid_0_6 : _GEN_10288; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11318 = 3'h3 == state ? valid_0_7 : _GEN_10289; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11319 = 3'h3 == state ? valid_0_8 : _GEN_10290; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11320 = 3'h3 == state ? valid_0_9 : _GEN_10291; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11321 = 3'h3 == state ? valid_0_10 : _GEN_10292; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11322 = 3'h3 == state ? valid_0_11 : _GEN_10293; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11323 = 3'h3 == state ? valid_0_12 : _GEN_10294; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11324 = 3'h3 == state ? valid_0_13 : _GEN_10295; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11325 = 3'h3 == state ? valid_0_14 : _GEN_10296; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11326 = 3'h3 == state ? valid_0_15 : _GEN_10297; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11327 = 3'h3 == state ? valid_0_16 : _GEN_10298; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11328 = 3'h3 == state ? valid_0_17 : _GEN_10299; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11329 = 3'h3 == state ? valid_0_18 : _GEN_10300; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11330 = 3'h3 == state ? valid_0_19 : _GEN_10301; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11331 = 3'h3 == state ? valid_0_20 : _GEN_10302; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11332 = 3'h3 == state ? valid_0_21 : _GEN_10303; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11333 = 3'h3 == state ? valid_0_22 : _GEN_10304; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11334 = 3'h3 == state ? valid_0_23 : _GEN_10305; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11335 = 3'h3 == state ? valid_0_24 : _GEN_10306; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11336 = 3'h3 == state ? valid_0_25 : _GEN_10307; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11337 = 3'h3 == state ? valid_0_26 : _GEN_10308; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11338 = 3'h3 == state ? valid_0_27 : _GEN_10309; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11339 = 3'h3 == state ? valid_0_28 : _GEN_10310; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11340 = 3'h3 == state ? valid_0_29 : _GEN_10311; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11341 = 3'h3 == state ? valid_0_30 : _GEN_10312; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11342 = 3'h3 == state ? valid_0_31 : _GEN_10313; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11343 = 3'h3 == state ? valid_0_32 : _GEN_10314; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11344 = 3'h3 == state ? valid_0_33 : _GEN_10315; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11345 = 3'h3 == state ? valid_0_34 : _GEN_10316; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11346 = 3'h3 == state ? valid_0_35 : _GEN_10317; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11347 = 3'h3 == state ? valid_0_36 : _GEN_10318; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11348 = 3'h3 == state ? valid_0_37 : _GEN_10319; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11349 = 3'h3 == state ? valid_0_38 : _GEN_10320; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11350 = 3'h3 == state ? valid_0_39 : _GEN_10321; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11351 = 3'h3 == state ? valid_0_40 : _GEN_10322; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11352 = 3'h3 == state ? valid_0_41 : _GEN_10323; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11353 = 3'h3 == state ? valid_0_42 : _GEN_10324; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11354 = 3'h3 == state ? valid_0_43 : _GEN_10325; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11355 = 3'h3 == state ? valid_0_44 : _GEN_10326; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11356 = 3'h3 == state ? valid_0_45 : _GEN_10327; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11357 = 3'h3 == state ? valid_0_46 : _GEN_10328; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11358 = 3'h3 == state ? valid_0_47 : _GEN_10329; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11359 = 3'h3 == state ? valid_0_48 : _GEN_10330; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11360 = 3'h3 == state ? valid_0_49 : _GEN_10331; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11361 = 3'h3 == state ? valid_0_50 : _GEN_10332; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11362 = 3'h3 == state ? valid_0_51 : _GEN_10333; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11363 = 3'h3 == state ? valid_0_52 : _GEN_10334; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11364 = 3'h3 == state ? valid_0_53 : _GEN_10335; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11365 = 3'h3 == state ? valid_0_54 : _GEN_10336; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11366 = 3'h3 == state ? valid_0_55 : _GEN_10337; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11367 = 3'h3 == state ? valid_0_56 : _GEN_10338; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11368 = 3'h3 == state ? valid_0_57 : _GEN_10339; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11369 = 3'h3 == state ? valid_0_58 : _GEN_10340; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11370 = 3'h3 == state ? valid_0_59 : _GEN_10341; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11371 = 3'h3 == state ? valid_0_60 : _GEN_10342; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11372 = 3'h3 == state ? valid_0_61 : _GEN_10343; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11373 = 3'h3 == state ? valid_0_62 : _GEN_10344; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11374 = 3'h3 == state ? valid_0_63 : _GEN_10345; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11375 = 3'h3 == state ? valid_0_64 : _GEN_10346; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11376 = 3'h3 == state ? valid_0_65 : _GEN_10347; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11377 = 3'h3 == state ? valid_0_66 : _GEN_10348; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11378 = 3'h3 == state ? valid_0_67 : _GEN_10349; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11379 = 3'h3 == state ? valid_0_68 : _GEN_10350; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11380 = 3'h3 == state ? valid_0_69 : _GEN_10351; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11381 = 3'h3 == state ? valid_0_70 : _GEN_10352; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11382 = 3'h3 == state ? valid_0_71 : _GEN_10353; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11383 = 3'h3 == state ? valid_0_72 : _GEN_10354; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11384 = 3'h3 == state ? valid_0_73 : _GEN_10355; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11385 = 3'h3 == state ? valid_0_74 : _GEN_10356; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11386 = 3'h3 == state ? valid_0_75 : _GEN_10357; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11387 = 3'h3 == state ? valid_0_76 : _GEN_10358; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11388 = 3'h3 == state ? valid_0_77 : _GEN_10359; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11389 = 3'h3 == state ? valid_0_78 : _GEN_10360; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11390 = 3'h3 == state ? valid_0_79 : _GEN_10361; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11391 = 3'h3 == state ? valid_0_80 : _GEN_10362; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11392 = 3'h3 == state ? valid_0_81 : _GEN_10363; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11393 = 3'h3 == state ? valid_0_82 : _GEN_10364; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11394 = 3'h3 == state ? valid_0_83 : _GEN_10365; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11395 = 3'h3 == state ? valid_0_84 : _GEN_10366; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11396 = 3'h3 == state ? valid_0_85 : _GEN_10367; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11397 = 3'h3 == state ? valid_0_86 : _GEN_10368; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11398 = 3'h3 == state ? valid_0_87 : _GEN_10369; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11399 = 3'h3 == state ? valid_0_88 : _GEN_10370; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11400 = 3'h3 == state ? valid_0_89 : _GEN_10371; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11401 = 3'h3 == state ? valid_0_90 : _GEN_10372; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11402 = 3'h3 == state ? valid_0_91 : _GEN_10373; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11403 = 3'h3 == state ? valid_0_92 : _GEN_10374; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11404 = 3'h3 == state ? valid_0_93 : _GEN_10375; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11405 = 3'h3 == state ? valid_0_94 : _GEN_10376; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11406 = 3'h3 == state ? valid_0_95 : _GEN_10377; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11407 = 3'h3 == state ? valid_0_96 : _GEN_10378; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11408 = 3'h3 == state ? valid_0_97 : _GEN_10379; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11409 = 3'h3 == state ? valid_0_98 : _GEN_10380; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11410 = 3'h3 == state ? valid_0_99 : _GEN_10381; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11411 = 3'h3 == state ? valid_0_100 : _GEN_10382; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11412 = 3'h3 == state ? valid_0_101 : _GEN_10383; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11413 = 3'h3 == state ? valid_0_102 : _GEN_10384; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11414 = 3'h3 == state ? valid_0_103 : _GEN_10385; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11415 = 3'h3 == state ? valid_0_104 : _GEN_10386; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11416 = 3'h3 == state ? valid_0_105 : _GEN_10387; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11417 = 3'h3 == state ? valid_0_106 : _GEN_10388; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11418 = 3'h3 == state ? valid_0_107 : _GEN_10389; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11419 = 3'h3 == state ? valid_0_108 : _GEN_10390; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11420 = 3'h3 == state ? valid_0_109 : _GEN_10391; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11421 = 3'h3 == state ? valid_0_110 : _GEN_10392; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11422 = 3'h3 == state ? valid_0_111 : _GEN_10393; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11423 = 3'h3 == state ? valid_0_112 : _GEN_10394; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11424 = 3'h3 == state ? valid_0_113 : _GEN_10395; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11425 = 3'h3 == state ? valid_0_114 : _GEN_10396; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11426 = 3'h3 == state ? valid_0_115 : _GEN_10397; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11427 = 3'h3 == state ? valid_0_116 : _GEN_10398; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11428 = 3'h3 == state ? valid_0_117 : _GEN_10399; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11429 = 3'h3 == state ? valid_0_118 : _GEN_10400; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11430 = 3'h3 == state ? valid_0_119 : _GEN_10401; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11431 = 3'h3 == state ? valid_0_120 : _GEN_10402; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11432 = 3'h3 == state ? valid_0_121 : _GEN_10403; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11433 = 3'h3 == state ? valid_0_122 : _GEN_10404; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11434 = 3'h3 == state ? valid_0_123 : _GEN_10405; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11435 = 3'h3 == state ? valid_0_124 : _GEN_10406; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11436 = 3'h3 == state ? valid_0_125 : _GEN_10407; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11437 = 3'h3 == state ? valid_0_126 : _GEN_10408; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11438 = 3'h3 == state ? valid_0_127 : _GEN_10409; // @[d_cache.scala 64:18 22:26]
  wire  _GEN_11439 = 3'h3 == state ? quene : _GEN_10410; // @[d_cache.scala 64:18 35:24]
  wire [63:0] _GEN_11440 = 3'h3 == state ? ram_1_0 : _GEN_10411; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11441 = 3'h3 == state ? ram_1_1 : _GEN_10412; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11442 = 3'h3 == state ? ram_1_2 : _GEN_10413; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11443 = 3'h3 == state ? ram_1_3 : _GEN_10414; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11444 = 3'h3 == state ? ram_1_4 : _GEN_10415; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11445 = 3'h3 == state ? ram_1_5 : _GEN_10416; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11446 = 3'h3 == state ? ram_1_6 : _GEN_10417; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11447 = 3'h3 == state ? ram_1_7 : _GEN_10418; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11448 = 3'h3 == state ? ram_1_8 : _GEN_10419; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11449 = 3'h3 == state ? ram_1_9 : _GEN_10420; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11450 = 3'h3 == state ? ram_1_10 : _GEN_10421; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11451 = 3'h3 == state ? ram_1_11 : _GEN_10422; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11452 = 3'h3 == state ? ram_1_12 : _GEN_10423; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11453 = 3'h3 == state ? ram_1_13 : _GEN_10424; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11454 = 3'h3 == state ? ram_1_14 : _GEN_10425; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11455 = 3'h3 == state ? ram_1_15 : _GEN_10426; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11456 = 3'h3 == state ? ram_1_16 : _GEN_10427; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11457 = 3'h3 == state ? ram_1_17 : _GEN_10428; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11458 = 3'h3 == state ? ram_1_18 : _GEN_10429; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11459 = 3'h3 == state ? ram_1_19 : _GEN_10430; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11460 = 3'h3 == state ? ram_1_20 : _GEN_10431; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11461 = 3'h3 == state ? ram_1_21 : _GEN_10432; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11462 = 3'h3 == state ? ram_1_22 : _GEN_10433; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11463 = 3'h3 == state ? ram_1_23 : _GEN_10434; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11464 = 3'h3 == state ? ram_1_24 : _GEN_10435; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11465 = 3'h3 == state ? ram_1_25 : _GEN_10436; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11466 = 3'h3 == state ? ram_1_26 : _GEN_10437; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11467 = 3'h3 == state ? ram_1_27 : _GEN_10438; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11468 = 3'h3 == state ? ram_1_28 : _GEN_10439; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11469 = 3'h3 == state ? ram_1_29 : _GEN_10440; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11470 = 3'h3 == state ? ram_1_30 : _GEN_10441; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11471 = 3'h3 == state ? ram_1_31 : _GEN_10442; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11472 = 3'h3 == state ? ram_1_32 : _GEN_10443; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11473 = 3'h3 == state ? ram_1_33 : _GEN_10444; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11474 = 3'h3 == state ? ram_1_34 : _GEN_10445; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11475 = 3'h3 == state ? ram_1_35 : _GEN_10446; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11476 = 3'h3 == state ? ram_1_36 : _GEN_10447; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11477 = 3'h3 == state ? ram_1_37 : _GEN_10448; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11478 = 3'h3 == state ? ram_1_38 : _GEN_10449; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11479 = 3'h3 == state ? ram_1_39 : _GEN_10450; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11480 = 3'h3 == state ? ram_1_40 : _GEN_10451; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11481 = 3'h3 == state ? ram_1_41 : _GEN_10452; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11482 = 3'h3 == state ? ram_1_42 : _GEN_10453; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11483 = 3'h3 == state ? ram_1_43 : _GEN_10454; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11484 = 3'h3 == state ? ram_1_44 : _GEN_10455; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11485 = 3'h3 == state ? ram_1_45 : _GEN_10456; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11486 = 3'h3 == state ? ram_1_46 : _GEN_10457; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11487 = 3'h3 == state ? ram_1_47 : _GEN_10458; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11488 = 3'h3 == state ? ram_1_48 : _GEN_10459; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11489 = 3'h3 == state ? ram_1_49 : _GEN_10460; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11490 = 3'h3 == state ? ram_1_50 : _GEN_10461; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11491 = 3'h3 == state ? ram_1_51 : _GEN_10462; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11492 = 3'h3 == state ? ram_1_52 : _GEN_10463; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11493 = 3'h3 == state ? ram_1_53 : _GEN_10464; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11494 = 3'h3 == state ? ram_1_54 : _GEN_10465; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11495 = 3'h3 == state ? ram_1_55 : _GEN_10466; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11496 = 3'h3 == state ? ram_1_56 : _GEN_10467; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11497 = 3'h3 == state ? ram_1_57 : _GEN_10468; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11498 = 3'h3 == state ? ram_1_58 : _GEN_10469; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11499 = 3'h3 == state ? ram_1_59 : _GEN_10470; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11500 = 3'h3 == state ? ram_1_60 : _GEN_10471; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11501 = 3'h3 == state ? ram_1_61 : _GEN_10472; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11502 = 3'h3 == state ? ram_1_62 : _GEN_10473; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11503 = 3'h3 == state ? ram_1_63 : _GEN_10474; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11504 = 3'h3 == state ? ram_1_64 : _GEN_10475; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11505 = 3'h3 == state ? ram_1_65 : _GEN_10476; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11506 = 3'h3 == state ? ram_1_66 : _GEN_10477; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11507 = 3'h3 == state ? ram_1_67 : _GEN_10478; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11508 = 3'h3 == state ? ram_1_68 : _GEN_10479; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11509 = 3'h3 == state ? ram_1_69 : _GEN_10480; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11510 = 3'h3 == state ? ram_1_70 : _GEN_10481; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11511 = 3'h3 == state ? ram_1_71 : _GEN_10482; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11512 = 3'h3 == state ? ram_1_72 : _GEN_10483; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11513 = 3'h3 == state ? ram_1_73 : _GEN_10484; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11514 = 3'h3 == state ? ram_1_74 : _GEN_10485; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11515 = 3'h3 == state ? ram_1_75 : _GEN_10486; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11516 = 3'h3 == state ? ram_1_76 : _GEN_10487; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11517 = 3'h3 == state ? ram_1_77 : _GEN_10488; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11518 = 3'h3 == state ? ram_1_78 : _GEN_10489; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11519 = 3'h3 == state ? ram_1_79 : _GEN_10490; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11520 = 3'h3 == state ? ram_1_80 : _GEN_10491; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11521 = 3'h3 == state ? ram_1_81 : _GEN_10492; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11522 = 3'h3 == state ? ram_1_82 : _GEN_10493; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11523 = 3'h3 == state ? ram_1_83 : _GEN_10494; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11524 = 3'h3 == state ? ram_1_84 : _GEN_10495; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11525 = 3'h3 == state ? ram_1_85 : _GEN_10496; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11526 = 3'h3 == state ? ram_1_86 : _GEN_10497; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11527 = 3'h3 == state ? ram_1_87 : _GEN_10498; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11528 = 3'h3 == state ? ram_1_88 : _GEN_10499; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11529 = 3'h3 == state ? ram_1_89 : _GEN_10500; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11530 = 3'h3 == state ? ram_1_90 : _GEN_10501; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11531 = 3'h3 == state ? ram_1_91 : _GEN_10502; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11532 = 3'h3 == state ? ram_1_92 : _GEN_10503; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11533 = 3'h3 == state ? ram_1_93 : _GEN_10504; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11534 = 3'h3 == state ? ram_1_94 : _GEN_10505; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11535 = 3'h3 == state ? ram_1_95 : _GEN_10506; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11536 = 3'h3 == state ? ram_1_96 : _GEN_10507; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11537 = 3'h3 == state ? ram_1_97 : _GEN_10508; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11538 = 3'h3 == state ? ram_1_98 : _GEN_10509; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11539 = 3'h3 == state ? ram_1_99 : _GEN_10510; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11540 = 3'h3 == state ? ram_1_100 : _GEN_10511; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11541 = 3'h3 == state ? ram_1_101 : _GEN_10512; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11542 = 3'h3 == state ? ram_1_102 : _GEN_10513; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11543 = 3'h3 == state ? ram_1_103 : _GEN_10514; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11544 = 3'h3 == state ? ram_1_104 : _GEN_10515; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11545 = 3'h3 == state ? ram_1_105 : _GEN_10516; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11546 = 3'h3 == state ? ram_1_106 : _GEN_10517; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11547 = 3'h3 == state ? ram_1_107 : _GEN_10518; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11548 = 3'h3 == state ? ram_1_108 : _GEN_10519; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11549 = 3'h3 == state ? ram_1_109 : _GEN_10520; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11550 = 3'h3 == state ? ram_1_110 : _GEN_10521; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11551 = 3'h3 == state ? ram_1_111 : _GEN_10522; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11552 = 3'h3 == state ? ram_1_112 : _GEN_10523; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11553 = 3'h3 == state ? ram_1_113 : _GEN_10524; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11554 = 3'h3 == state ? ram_1_114 : _GEN_10525; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11555 = 3'h3 == state ? ram_1_115 : _GEN_10526; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11556 = 3'h3 == state ? ram_1_116 : _GEN_10527; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11557 = 3'h3 == state ? ram_1_117 : _GEN_10528; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11558 = 3'h3 == state ? ram_1_118 : _GEN_10529; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11559 = 3'h3 == state ? ram_1_119 : _GEN_10530; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11560 = 3'h3 == state ? ram_1_120 : _GEN_10531; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11561 = 3'h3 == state ? ram_1_121 : _GEN_10532; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11562 = 3'h3 == state ? ram_1_122 : _GEN_10533; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11563 = 3'h3 == state ? ram_1_123 : _GEN_10534; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11564 = 3'h3 == state ? ram_1_124 : _GEN_10535; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11565 = 3'h3 == state ? ram_1_125 : _GEN_10536; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11566 = 3'h3 == state ? ram_1_126 : _GEN_10537; // @[d_cache.scala 64:18 19:24]
  wire [63:0] _GEN_11567 = 3'h3 == state ? ram_1_127 : _GEN_10538; // @[d_cache.scala 64:18 19:24]
  wire [31:0] _GEN_11568 = 3'h3 == state ? tag_1_0 : _GEN_10539; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11569 = 3'h3 == state ? tag_1_1 : _GEN_10540; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11570 = 3'h3 == state ? tag_1_2 : _GEN_10541; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11571 = 3'h3 == state ? tag_1_3 : _GEN_10542; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11572 = 3'h3 == state ? tag_1_4 : _GEN_10543; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11573 = 3'h3 == state ? tag_1_5 : _GEN_10544; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11574 = 3'h3 == state ? tag_1_6 : _GEN_10545; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11575 = 3'h3 == state ? tag_1_7 : _GEN_10546; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11576 = 3'h3 == state ? tag_1_8 : _GEN_10547; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11577 = 3'h3 == state ? tag_1_9 : _GEN_10548; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11578 = 3'h3 == state ? tag_1_10 : _GEN_10549; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11579 = 3'h3 == state ? tag_1_11 : _GEN_10550; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11580 = 3'h3 == state ? tag_1_12 : _GEN_10551; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11581 = 3'h3 == state ? tag_1_13 : _GEN_10552; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11582 = 3'h3 == state ? tag_1_14 : _GEN_10553; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11583 = 3'h3 == state ? tag_1_15 : _GEN_10554; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11584 = 3'h3 == state ? tag_1_16 : _GEN_10555; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11585 = 3'h3 == state ? tag_1_17 : _GEN_10556; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11586 = 3'h3 == state ? tag_1_18 : _GEN_10557; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11587 = 3'h3 == state ? tag_1_19 : _GEN_10558; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11588 = 3'h3 == state ? tag_1_20 : _GEN_10559; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11589 = 3'h3 == state ? tag_1_21 : _GEN_10560; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11590 = 3'h3 == state ? tag_1_22 : _GEN_10561; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11591 = 3'h3 == state ? tag_1_23 : _GEN_10562; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11592 = 3'h3 == state ? tag_1_24 : _GEN_10563; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11593 = 3'h3 == state ? tag_1_25 : _GEN_10564; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11594 = 3'h3 == state ? tag_1_26 : _GEN_10565; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11595 = 3'h3 == state ? tag_1_27 : _GEN_10566; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11596 = 3'h3 == state ? tag_1_28 : _GEN_10567; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11597 = 3'h3 == state ? tag_1_29 : _GEN_10568; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11598 = 3'h3 == state ? tag_1_30 : _GEN_10569; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11599 = 3'h3 == state ? tag_1_31 : _GEN_10570; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11600 = 3'h3 == state ? tag_1_32 : _GEN_10571; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11601 = 3'h3 == state ? tag_1_33 : _GEN_10572; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11602 = 3'h3 == state ? tag_1_34 : _GEN_10573; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11603 = 3'h3 == state ? tag_1_35 : _GEN_10574; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11604 = 3'h3 == state ? tag_1_36 : _GEN_10575; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11605 = 3'h3 == state ? tag_1_37 : _GEN_10576; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11606 = 3'h3 == state ? tag_1_38 : _GEN_10577; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11607 = 3'h3 == state ? tag_1_39 : _GEN_10578; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11608 = 3'h3 == state ? tag_1_40 : _GEN_10579; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11609 = 3'h3 == state ? tag_1_41 : _GEN_10580; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11610 = 3'h3 == state ? tag_1_42 : _GEN_10581; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11611 = 3'h3 == state ? tag_1_43 : _GEN_10582; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11612 = 3'h3 == state ? tag_1_44 : _GEN_10583; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11613 = 3'h3 == state ? tag_1_45 : _GEN_10584; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11614 = 3'h3 == state ? tag_1_46 : _GEN_10585; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11615 = 3'h3 == state ? tag_1_47 : _GEN_10586; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11616 = 3'h3 == state ? tag_1_48 : _GEN_10587; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11617 = 3'h3 == state ? tag_1_49 : _GEN_10588; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11618 = 3'h3 == state ? tag_1_50 : _GEN_10589; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11619 = 3'h3 == state ? tag_1_51 : _GEN_10590; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11620 = 3'h3 == state ? tag_1_52 : _GEN_10591; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11621 = 3'h3 == state ? tag_1_53 : _GEN_10592; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11622 = 3'h3 == state ? tag_1_54 : _GEN_10593; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11623 = 3'h3 == state ? tag_1_55 : _GEN_10594; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11624 = 3'h3 == state ? tag_1_56 : _GEN_10595; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11625 = 3'h3 == state ? tag_1_57 : _GEN_10596; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11626 = 3'h3 == state ? tag_1_58 : _GEN_10597; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11627 = 3'h3 == state ? tag_1_59 : _GEN_10598; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11628 = 3'h3 == state ? tag_1_60 : _GEN_10599; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11629 = 3'h3 == state ? tag_1_61 : _GEN_10600; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11630 = 3'h3 == state ? tag_1_62 : _GEN_10601; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11631 = 3'h3 == state ? tag_1_63 : _GEN_10602; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11632 = 3'h3 == state ? tag_1_64 : _GEN_10603; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11633 = 3'h3 == state ? tag_1_65 : _GEN_10604; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11634 = 3'h3 == state ? tag_1_66 : _GEN_10605; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11635 = 3'h3 == state ? tag_1_67 : _GEN_10606; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11636 = 3'h3 == state ? tag_1_68 : _GEN_10607; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11637 = 3'h3 == state ? tag_1_69 : _GEN_10608; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11638 = 3'h3 == state ? tag_1_70 : _GEN_10609; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11639 = 3'h3 == state ? tag_1_71 : _GEN_10610; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11640 = 3'h3 == state ? tag_1_72 : _GEN_10611; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11641 = 3'h3 == state ? tag_1_73 : _GEN_10612; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11642 = 3'h3 == state ? tag_1_74 : _GEN_10613; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11643 = 3'h3 == state ? tag_1_75 : _GEN_10614; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11644 = 3'h3 == state ? tag_1_76 : _GEN_10615; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11645 = 3'h3 == state ? tag_1_77 : _GEN_10616; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11646 = 3'h3 == state ? tag_1_78 : _GEN_10617; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11647 = 3'h3 == state ? tag_1_79 : _GEN_10618; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11648 = 3'h3 == state ? tag_1_80 : _GEN_10619; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11649 = 3'h3 == state ? tag_1_81 : _GEN_10620; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11650 = 3'h3 == state ? tag_1_82 : _GEN_10621; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11651 = 3'h3 == state ? tag_1_83 : _GEN_10622; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11652 = 3'h3 == state ? tag_1_84 : _GEN_10623; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11653 = 3'h3 == state ? tag_1_85 : _GEN_10624; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11654 = 3'h3 == state ? tag_1_86 : _GEN_10625; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11655 = 3'h3 == state ? tag_1_87 : _GEN_10626; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11656 = 3'h3 == state ? tag_1_88 : _GEN_10627; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11657 = 3'h3 == state ? tag_1_89 : _GEN_10628; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11658 = 3'h3 == state ? tag_1_90 : _GEN_10629; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11659 = 3'h3 == state ? tag_1_91 : _GEN_10630; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11660 = 3'h3 == state ? tag_1_92 : _GEN_10631; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11661 = 3'h3 == state ? tag_1_93 : _GEN_10632; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11662 = 3'h3 == state ? tag_1_94 : _GEN_10633; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11663 = 3'h3 == state ? tag_1_95 : _GEN_10634; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11664 = 3'h3 == state ? tag_1_96 : _GEN_10635; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11665 = 3'h3 == state ? tag_1_97 : _GEN_10636; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11666 = 3'h3 == state ? tag_1_98 : _GEN_10637; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11667 = 3'h3 == state ? tag_1_99 : _GEN_10638; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11668 = 3'h3 == state ? tag_1_100 : _GEN_10639; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11669 = 3'h3 == state ? tag_1_101 : _GEN_10640; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11670 = 3'h3 == state ? tag_1_102 : _GEN_10641; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11671 = 3'h3 == state ? tag_1_103 : _GEN_10642; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11672 = 3'h3 == state ? tag_1_104 : _GEN_10643; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11673 = 3'h3 == state ? tag_1_105 : _GEN_10644; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11674 = 3'h3 == state ? tag_1_106 : _GEN_10645; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11675 = 3'h3 == state ? tag_1_107 : _GEN_10646; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11676 = 3'h3 == state ? tag_1_108 : _GEN_10647; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11677 = 3'h3 == state ? tag_1_109 : _GEN_10648; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11678 = 3'h3 == state ? tag_1_110 : _GEN_10649; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11679 = 3'h3 == state ? tag_1_111 : _GEN_10650; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11680 = 3'h3 == state ? tag_1_112 : _GEN_10651; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11681 = 3'h3 == state ? tag_1_113 : _GEN_10652; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11682 = 3'h3 == state ? tag_1_114 : _GEN_10653; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11683 = 3'h3 == state ? tag_1_115 : _GEN_10654; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11684 = 3'h3 == state ? tag_1_116 : _GEN_10655; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11685 = 3'h3 == state ? tag_1_117 : _GEN_10656; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11686 = 3'h3 == state ? tag_1_118 : _GEN_10657; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11687 = 3'h3 == state ? tag_1_119 : _GEN_10658; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11688 = 3'h3 == state ? tag_1_120 : _GEN_10659; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11689 = 3'h3 == state ? tag_1_121 : _GEN_10660; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11690 = 3'h3 == state ? tag_1_122 : _GEN_10661; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11691 = 3'h3 == state ? tag_1_123 : _GEN_10662; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11692 = 3'h3 == state ? tag_1_124 : _GEN_10663; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11693 = 3'h3 == state ? tag_1_125 : _GEN_10664; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11694 = 3'h3 == state ? tag_1_126 : _GEN_10665; // @[d_cache.scala 64:18 21:24]
  wire [31:0] _GEN_11695 = 3'h3 == state ? tag_1_127 : _GEN_10666; // @[d_cache.scala 64:18 21:24]
  wire  _GEN_11696 = 3'h3 == state ? valid_1_0 : _GEN_10667; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11697 = 3'h3 == state ? valid_1_1 : _GEN_10668; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11698 = 3'h3 == state ? valid_1_2 : _GEN_10669; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11699 = 3'h3 == state ? valid_1_3 : _GEN_10670; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11700 = 3'h3 == state ? valid_1_4 : _GEN_10671; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11701 = 3'h3 == state ? valid_1_5 : _GEN_10672; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11702 = 3'h3 == state ? valid_1_6 : _GEN_10673; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11703 = 3'h3 == state ? valid_1_7 : _GEN_10674; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11704 = 3'h3 == state ? valid_1_8 : _GEN_10675; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11705 = 3'h3 == state ? valid_1_9 : _GEN_10676; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11706 = 3'h3 == state ? valid_1_10 : _GEN_10677; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11707 = 3'h3 == state ? valid_1_11 : _GEN_10678; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11708 = 3'h3 == state ? valid_1_12 : _GEN_10679; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11709 = 3'h3 == state ? valid_1_13 : _GEN_10680; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11710 = 3'h3 == state ? valid_1_14 : _GEN_10681; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11711 = 3'h3 == state ? valid_1_15 : _GEN_10682; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11712 = 3'h3 == state ? valid_1_16 : _GEN_10683; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11713 = 3'h3 == state ? valid_1_17 : _GEN_10684; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11714 = 3'h3 == state ? valid_1_18 : _GEN_10685; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11715 = 3'h3 == state ? valid_1_19 : _GEN_10686; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11716 = 3'h3 == state ? valid_1_20 : _GEN_10687; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11717 = 3'h3 == state ? valid_1_21 : _GEN_10688; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11718 = 3'h3 == state ? valid_1_22 : _GEN_10689; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11719 = 3'h3 == state ? valid_1_23 : _GEN_10690; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11720 = 3'h3 == state ? valid_1_24 : _GEN_10691; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11721 = 3'h3 == state ? valid_1_25 : _GEN_10692; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11722 = 3'h3 == state ? valid_1_26 : _GEN_10693; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11723 = 3'h3 == state ? valid_1_27 : _GEN_10694; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11724 = 3'h3 == state ? valid_1_28 : _GEN_10695; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11725 = 3'h3 == state ? valid_1_29 : _GEN_10696; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11726 = 3'h3 == state ? valid_1_30 : _GEN_10697; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11727 = 3'h3 == state ? valid_1_31 : _GEN_10698; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11728 = 3'h3 == state ? valid_1_32 : _GEN_10699; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11729 = 3'h3 == state ? valid_1_33 : _GEN_10700; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11730 = 3'h3 == state ? valid_1_34 : _GEN_10701; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11731 = 3'h3 == state ? valid_1_35 : _GEN_10702; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11732 = 3'h3 == state ? valid_1_36 : _GEN_10703; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11733 = 3'h3 == state ? valid_1_37 : _GEN_10704; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11734 = 3'h3 == state ? valid_1_38 : _GEN_10705; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11735 = 3'h3 == state ? valid_1_39 : _GEN_10706; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11736 = 3'h3 == state ? valid_1_40 : _GEN_10707; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11737 = 3'h3 == state ? valid_1_41 : _GEN_10708; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11738 = 3'h3 == state ? valid_1_42 : _GEN_10709; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11739 = 3'h3 == state ? valid_1_43 : _GEN_10710; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11740 = 3'h3 == state ? valid_1_44 : _GEN_10711; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11741 = 3'h3 == state ? valid_1_45 : _GEN_10712; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11742 = 3'h3 == state ? valid_1_46 : _GEN_10713; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11743 = 3'h3 == state ? valid_1_47 : _GEN_10714; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11744 = 3'h3 == state ? valid_1_48 : _GEN_10715; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11745 = 3'h3 == state ? valid_1_49 : _GEN_10716; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11746 = 3'h3 == state ? valid_1_50 : _GEN_10717; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11747 = 3'h3 == state ? valid_1_51 : _GEN_10718; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11748 = 3'h3 == state ? valid_1_52 : _GEN_10719; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11749 = 3'h3 == state ? valid_1_53 : _GEN_10720; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11750 = 3'h3 == state ? valid_1_54 : _GEN_10721; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11751 = 3'h3 == state ? valid_1_55 : _GEN_10722; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11752 = 3'h3 == state ? valid_1_56 : _GEN_10723; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11753 = 3'h3 == state ? valid_1_57 : _GEN_10724; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11754 = 3'h3 == state ? valid_1_58 : _GEN_10725; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11755 = 3'h3 == state ? valid_1_59 : _GEN_10726; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11756 = 3'h3 == state ? valid_1_60 : _GEN_10727; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11757 = 3'h3 == state ? valid_1_61 : _GEN_10728; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11758 = 3'h3 == state ? valid_1_62 : _GEN_10729; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11759 = 3'h3 == state ? valid_1_63 : _GEN_10730; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11760 = 3'h3 == state ? valid_1_64 : _GEN_10731; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11761 = 3'h3 == state ? valid_1_65 : _GEN_10732; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11762 = 3'h3 == state ? valid_1_66 : _GEN_10733; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11763 = 3'h3 == state ? valid_1_67 : _GEN_10734; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11764 = 3'h3 == state ? valid_1_68 : _GEN_10735; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11765 = 3'h3 == state ? valid_1_69 : _GEN_10736; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11766 = 3'h3 == state ? valid_1_70 : _GEN_10737; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11767 = 3'h3 == state ? valid_1_71 : _GEN_10738; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11768 = 3'h3 == state ? valid_1_72 : _GEN_10739; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11769 = 3'h3 == state ? valid_1_73 : _GEN_10740; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11770 = 3'h3 == state ? valid_1_74 : _GEN_10741; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11771 = 3'h3 == state ? valid_1_75 : _GEN_10742; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11772 = 3'h3 == state ? valid_1_76 : _GEN_10743; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11773 = 3'h3 == state ? valid_1_77 : _GEN_10744; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11774 = 3'h3 == state ? valid_1_78 : _GEN_10745; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11775 = 3'h3 == state ? valid_1_79 : _GEN_10746; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11776 = 3'h3 == state ? valid_1_80 : _GEN_10747; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11777 = 3'h3 == state ? valid_1_81 : _GEN_10748; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11778 = 3'h3 == state ? valid_1_82 : _GEN_10749; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11779 = 3'h3 == state ? valid_1_83 : _GEN_10750; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11780 = 3'h3 == state ? valid_1_84 : _GEN_10751; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11781 = 3'h3 == state ? valid_1_85 : _GEN_10752; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11782 = 3'h3 == state ? valid_1_86 : _GEN_10753; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11783 = 3'h3 == state ? valid_1_87 : _GEN_10754; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11784 = 3'h3 == state ? valid_1_88 : _GEN_10755; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11785 = 3'h3 == state ? valid_1_89 : _GEN_10756; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11786 = 3'h3 == state ? valid_1_90 : _GEN_10757; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11787 = 3'h3 == state ? valid_1_91 : _GEN_10758; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11788 = 3'h3 == state ? valid_1_92 : _GEN_10759; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11789 = 3'h3 == state ? valid_1_93 : _GEN_10760; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11790 = 3'h3 == state ? valid_1_94 : _GEN_10761; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11791 = 3'h3 == state ? valid_1_95 : _GEN_10762; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11792 = 3'h3 == state ? valid_1_96 : _GEN_10763; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11793 = 3'h3 == state ? valid_1_97 : _GEN_10764; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11794 = 3'h3 == state ? valid_1_98 : _GEN_10765; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11795 = 3'h3 == state ? valid_1_99 : _GEN_10766; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11796 = 3'h3 == state ? valid_1_100 : _GEN_10767; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11797 = 3'h3 == state ? valid_1_101 : _GEN_10768; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11798 = 3'h3 == state ? valid_1_102 : _GEN_10769; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11799 = 3'h3 == state ? valid_1_103 : _GEN_10770; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11800 = 3'h3 == state ? valid_1_104 : _GEN_10771; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11801 = 3'h3 == state ? valid_1_105 : _GEN_10772; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11802 = 3'h3 == state ? valid_1_106 : _GEN_10773; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11803 = 3'h3 == state ? valid_1_107 : _GEN_10774; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11804 = 3'h3 == state ? valid_1_108 : _GEN_10775; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11805 = 3'h3 == state ? valid_1_109 : _GEN_10776; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11806 = 3'h3 == state ? valid_1_110 : _GEN_10777; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11807 = 3'h3 == state ? valid_1_111 : _GEN_10778; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11808 = 3'h3 == state ? valid_1_112 : _GEN_10779; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11809 = 3'h3 == state ? valid_1_113 : _GEN_10780; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11810 = 3'h3 == state ? valid_1_114 : _GEN_10781; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11811 = 3'h3 == state ? valid_1_115 : _GEN_10782; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11812 = 3'h3 == state ? valid_1_116 : _GEN_10783; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11813 = 3'h3 == state ? valid_1_117 : _GEN_10784; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11814 = 3'h3 == state ? valid_1_118 : _GEN_10785; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11815 = 3'h3 == state ? valid_1_119 : _GEN_10786; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11816 = 3'h3 == state ? valid_1_120 : _GEN_10787; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11817 = 3'h3 == state ? valid_1_121 : _GEN_10788; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11818 = 3'h3 == state ? valid_1_122 : _GEN_10789; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11819 = 3'h3 == state ? valid_1_123 : _GEN_10790; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11820 = 3'h3 == state ? valid_1_124 : _GEN_10791; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11821 = 3'h3 == state ? valid_1_125 : _GEN_10792; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11822 = 3'h3 == state ? valid_1_126 : _GEN_10793; // @[d_cache.scala 64:18 23:26]
  wire  _GEN_11823 = 3'h3 == state ? valid_1_127 : _GEN_10794; // @[d_cache.scala 64:18 23:26]
  wire [63:0] _GEN_11824 = 3'h3 == state ? write_back_data : _GEN_10795; // @[d_cache.scala 64:18 29:34]
  wire [38:0] _GEN_11825 = 3'h3 == state ? {{7'd0}, write_back_addr} : _GEN_10796; // @[d_cache.scala 64:18 30:34]
  wire  _GEN_11826 = 3'h3 == state ? dirty_0_0 : _GEN_10797; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11827 = 3'h3 == state ? dirty_0_1 : _GEN_10798; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11828 = 3'h3 == state ? dirty_0_2 : _GEN_10799; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11829 = 3'h3 == state ? dirty_0_3 : _GEN_10800; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11830 = 3'h3 == state ? dirty_0_4 : _GEN_10801; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11831 = 3'h3 == state ? dirty_0_5 : _GEN_10802; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11832 = 3'h3 == state ? dirty_0_6 : _GEN_10803; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11833 = 3'h3 == state ? dirty_0_7 : _GEN_10804; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11834 = 3'h3 == state ? dirty_0_8 : _GEN_10805; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11835 = 3'h3 == state ? dirty_0_9 : _GEN_10806; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11836 = 3'h3 == state ? dirty_0_10 : _GEN_10807; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11837 = 3'h3 == state ? dirty_0_11 : _GEN_10808; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11838 = 3'h3 == state ? dirty_0_12 : _GEN_10809; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11839 = 3'h3 == state ? dirty_0_13 : _GEN_10810; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11840 = 3'h3 == state ? dirty_0_14 : _GEN_10811; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11841 = 3'h3 == state ? dirty_0_15 : _GEN_10812; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11842 = 3'h3 == state ? dirty_0_16 : _GEN_10813; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11843 = 3'h3 == state ? dirty_0_17 : _GEN_10814; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11844 = 3'h3 == state ? dirty_0_18 : _GEN_10815; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11845 = 3'h3 == state ? dirty_0_19 : _GEN_10816; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11846 = 3'h3 == state ? dirty_0_20 : _GEN_10817; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11847 = 3'h3 == state ? dirty_0_21 : _GEN_10818; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11848 = 3'h3 == state ? dirty_0_22 : _GEN_10819; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11849 = 3'h3 == state ? dirty_0_23 : _GEN_10820; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11850 = 3'h3 == state ? dirty_0_24 : _GEN_10821; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11851 = 3'h3 == state ? dirty_0_25 : _GEN_10822; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11852 = 3'h3 == state ? dirty_0_26 : _GEN_10823; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11853 = 3'h3 == state ? dirty_0_27 : _GEN_10824; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11854 = 3'h3 == state ? dirty_0_28 : _GEN_10825; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11855 = 3'h3 == state ? dirty_0_29 : _GEN_10826; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11856 = 3'h3 == state ? dirty_0_30 : _GEN_10827; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11857 = 3'h3 == state ? dirty_0_31 : _GEN_10828; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11858 = 3'h3 == state ? dirty_0_32 : _GEN_10829; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11859 = 3'h3 == state ? dirty_0_33 : _GEN_10830; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11860 = 3'h3 == state ? dirty_0_34 : _GEN_10831; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11861 = 3'h3 == state ? dirty_0_35 : _GEN_10832; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11862 = 3'h3 == state ? dirty_0_36 : _GEN_10833; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11863 = 3'h3 == state ? dirty_0_37 : _GEN_10834; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11864 = 3'h3 == state ? dirty_0_38 : _GEN_10835; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11865 = 3'h3 == state ? dirty_0_39 : _GEN_10836; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11866 = 3'h3 == state ? dirty_0_40 : _GEN_10837; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11867 = 3'h3 == state ? dirty_0_41 : _GEN_10838; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11868 = 3'h3 == state ? dirty_0_42 : _GEN_10839; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11869 = 3'h3 == state ? dirty_0_43 : _GEN_10840; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11870 = 3'h3 == state ? dirty_0_44 : _GEN_10841; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11871 = 3'h3 == state ? dirty_0_45 : _GEN_10842; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11872 = 3'h3 == state ? dirty_0_46 : _GEN_10843; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11873 = 3'h3 == state ? dirty_0_47 : _GEN_10844; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11874 = 3'h3 == state ? dirty_0_48 : _GEN_10845; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11875 = 3'h3 == state ? dirty_0_49 : _GEN_10846; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11876 = 3'h3 == state ? dirty_0_50 : _GEN_10847; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11877 = 3'h3 == state ? dirty_0_51 : _GEN_10848; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11878 = 3'h3 == state ? dirty_0_52 : _GEN_10849; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11879 = 3'h3 == state ? dirty_0_53 : _GEN_10850; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11880 = 3'h3 == state ? dirty_0_54 : _GEN_10851; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11881 = 3'h3 == state ? dirty_0_55 : _GEN_10852; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11882 = 3'h3 == state ? dirty_0_56 : _GEN_10853; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11883 = 3'h3 == state ? dirty_0_57 : _GEN_10854; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11884 = 3'h3 == state ? dirty_0_58 : _GEN_10855; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11885 = 3'h3 == state ? dirty_0_59 : _GEN_10856; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11886 = 3'h3 == state ? dirty_0_60 : _GEN_10857; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11887 = 3'h3 == state ? dirty_0_61 : _GEN_10858; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11888 = 3'h3 == state ? dirty_0_62 : _GEN_10859; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11889 = 3'h3 == state ? dirty_0_63 : _GEN_10860; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11890 = 3'h3 == state ? dirty_0_64 : _GEN_10861; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11891 = 3'h3 == state ? dirty_0_65 : _GEN_10862; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11892 = 3'h3 == state ? dirty_0_66 : _GEN_10863; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11893 = 3'h3 == state ? dirty_0_67 : _GEN_10864; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11894 = 3'h3 == state ? dirty_0_68 : _GEN_10865; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11895 = 3'h3 == state ? dirty_0_69 : _GEN_10866; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11896 = 3'h3 == state ? dirty_0_70 : _GEN_10867; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11897 = 3'h3 == state ? dirty_0_71 : _GEN_10868; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11898 = 3'h3 == state ? dirty_0_72 : _GEN_10869; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11899 = 3'h3 == state ? dirty_0_73 : _GEN_10870; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11900 = 3'h3 == state ? dirty_0_74 : _GEN_10871; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11901 = 3'h3 == state ? dirty_0_75 : _GEN_10872; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11902 = 3'h3 == state ? dirty_0_76 : _GEN_10873; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11903 = 3'h3 == state ? dirty_0_77 : _GEN_10874; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11904 = 3'h3 == state ? dirty_0_78 : _GEN_10875; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11905 = 3'h3 == state ? dirty_0_79 : _GEN_10876; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11906 = 3'h3 == state ? dirty_0_80 : _GEN_10877; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11907 = 3'h3 == state ? dirty_0_81 : _GEN_10878; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11908 = 3'h3 == state ? dirty_0_82 : _GEN_10879; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11909 = 3'h3 == state ? dirty_0_83 : _GEN_10880; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11910 = 3'h3 == state ? dirty_0_84 : _GEN_10881; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11911 = 3'h3 == state ? dirty_0_85 : _GEN_10882; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11912 = 3'h3 == state ? dirty_0_86 : _GEN_10883; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11913 = 3'h3 == state ? dirty_0_87 : _GEN_10884; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11914 = 3'h3 == state ? dirty_0_88 : _GEN_10885; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11915 = 3'h3 == state ? dirty_0_89 : _GEN_10886; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11916 = 3'h3 == state ? dirty_0_90 : _GEN_10887; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11917 = 3'h3 == state ? dirty_0_91 : _GEN_10888; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11918 = 3'h3 == state ? dirty_0_92 : _GEN_10889; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11919 = 3'h3 == state ? dirty_0_93 : _GEN_10890; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11920 = 3'h3 == state ? dirty_0_94 : _GEN_10891; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11921 = 3'h3 == state ? dirty_0_95 : _GEN_10892; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11922 = 3'h3 == state ? dirty_0_96 : _GEN_10893; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11923 = 3'h3 == state ? dirty_0_97 : _GEN_10894; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11924 = 3'h3 == state ? dirty_0_98 : _GEN_10895; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11925 = 3'h3 == state ? dirty_0_99 : _GEN_10896; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11926 = 3'h3 == state ? dirty_0_100 : _GEN_10897; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11927 = 3'h3 == state ? dirty_0_101 : _GEN_10898; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11928 = 3'h3 == state ? dirty_0_102 : _GEN_10899; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11929 = 3'h3 == state ? dirty_0_103 : _GEN_10900; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11930 = 3'h3 == state ? dirty_0_104 : _GEN_10901; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11931 = 3'h3 == state ? dirty_0_105 : _GEN_10902; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11932 = 3'h3 == state ? dirty_0_106 : _GEN_10903; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11933 = 3'h3 == state ? dirty_0_107 : _GEN_10904; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11934 = 3'h3 == state ? dirty_0_108 : _GEN_10905; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11935 = 3'h3 == state ? dirty_0_109 : _GEN_10906; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11936 = 3'h3 == state ? dirty_0_110 : _GEN_10907; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11937 = 3'h3 == state ? dirty_0_111 : _GEN_10908; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11938 = 3'h3 == state ? dirty_0_112 : _GEN_10909; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11939 = 3'h3 == state ? dirty_0_113 : _GEN_10910; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11940 = 3'h3 == state ? dirty_0_114 : _GEN_10911; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11941 = 3'h3 == state ? dirty_0_115 : _GEN_10912; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11942 = 3'h3 == state ? dirty_0_116 : _GEN_10913; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11943 = 3'h3 == state ? dirty_0_117 : _GEN_10914; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11944 = 3'h3 == state ? dirty_0_118 : _GEN_10915; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11945 = 3'h3 == state ? dirty_0_119 : _GEN_10916; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11946 = 3'h3 == state ? dirty_0_120 : _GEN_10917; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11947 = 3'h3 == state ? dirty_0_121 : _GEN_10918; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11948 = 3'h3 == state ? dirty_0_122 : _GEN_10919; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11949 = 3'h3 == state ? dirty_0_123 : _GEN_10920; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11950 = 3'h3 == state ? dirty_0_124 : _GEN_10921; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11951 = 3'h3 == state ? dirty_0_125 : _GEN_10922; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11952 = 3'h3 == state ? dirty_0_126 : _GEN_10923; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11953 = 3'h3 == state ? dirty_0_127 : _GEN_10924; // @[d_cache.scala 64:18 24:26]
  wire  _GEN_11954 = 3'h3 == state ? dirty_1_0 : _GEN_10925; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11955 = 3'h3 == state ? dirty_1_1 : _GEN_10926; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11956 = 3'h3 == state ? dirty_1_2 : _GEN_10927; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11957 = 3'h3 == state ? dirty_1_3 : _GEN_10928; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11958 = 3'h3 == state ? dirty_1_4 : _GEN_10929; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11959 = 3'h3 == state ? dirty_1_5 : _GEN_10930; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11960 = 3'h3 == state ? dirty_1_6 : _GEN_10931; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11961 = 3'h3 == state ? dirty_1_7 : _GEN_10932; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11962 = 3'h3 == state ? dirty_1_8 : _GEN_10933; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11963 = 3'h3 == state ? dirty_1_9 : _GEN_10934; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11964 = 3'h3 == state ? dirty_1_10 : _GEN_10935; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11965 = 3'h3 == state ? dirty_1_11 : _GEN_10936; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11966 = 3'h3 == state ? dirty_1_12 : _GEN_10937; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11967 = 3'h3 == state ? dirty_1_13 : _GEN_10938; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11968 = 3'h3 == state ? dirty_1_14 : _GEN_10939; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11969 = 3'h3 == state ? dirty_1_15 : _GEN_10940; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11970 = 3'h3 == state ? dirty_1_16 : _GEN_10941; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11971 = 3'h3 == state ? dirty_1_17 : _GEN_10942; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11972 = 3'h3 == state ? dirty_1_18 : _GEN_10943; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11973 = 3'h3 == state ? dirty_1_19 : _GEN_10944; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11974 = 3'h3 == state ? dirty_1_20 : _GEN_10945; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11975 = 3'h3 == state ? dirty_1_21 : _GEN_10946; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11976 = 3'h3 == state ? dirty_1_22 : _GEN_10947; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11977 = 3'h3 == state ? dirty_1_23 : _GEN_10948; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11978 = 3'h3 == state ? dirty_1_24 : _GEN_10949; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11979 = 3'h3 == state ? dirty_1_25 : _GEN_10950; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11980 = 3'h3 == state ? dirty_1_26 : _GEN_10951; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11981 = 3'h3 == state ? dirty_1_27 : _GEN_10952; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11982 = 3'h3 == state ? dirty_1_28 : _GEN_10953; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11983 = 3'h3 == state ? dirty_1_29 : _GEN_10954; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11984 = 3'h3 == state ? dirty_1_30 : _GEN_10955; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11985 = 3'h3 == state ? dirty_1_31 : _GEN_10956; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11986 = 3'h3 == state ? dirty_1_32 : _GEN_10957; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11987 = 3'h3 == state ? dirty_1_33 : _GEN_10958; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11988 = 3'h3 == state ? dirty_1_34 : _GEN_10959; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11989 = 3'h3 == state ? dirty_1_35 : _GEN_10960; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11990 = 3'h3 == state ? dirty_1_36 : _GEN_10961; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11991 = 3'h3 == state ? dirty_1_37 : _GEN_10962; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11992 = 3'h3 == state ? dirty_1_38 : _GEN_10963; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11993 = 3'h3 == state ? dirty_1_39 : _GEN_10964; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11994 = 3'h3 == state ? dirty_1_40 : _GEN_10965; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11995 = 3'h3 == state ? dirty_1_41 : _GEN_10966; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11996 = 3'h3 == state ? dirty_1_42 : _GEN_10967; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11997 = 3'h3 == state ? dirty_1_43 : _GEN_10968; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11998 = 3'h3 == state ? dirty_1_44 : _GEN_10969; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_11999 = 3'h3 == state ? dirty_1_45 : _GEN_10970; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12000 = 3'h3 == state ? dirty_1_46 : _GEN_10971; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12001 = 3'h3 == state ? dirty_1_47 : _GEN_10972; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12002 = 3'h3 == state ? dirty_1_48 : _GEN_10973; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12003 = 3'h3 == state ? dirty_1_49 : _GEN_10974; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12004 = 3'h3 == state ? dirty_1_50 : _GEN_10975; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12005 = 3'h3 == state ? dirty_1_51 : _GEN_10976; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12006 = 3'h3 == state ? dirty_1_52 : _GEN_10977; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12007 = 3'h3 == state ? dirty_1_53 : _GEN_10978; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12008 = 3'h3 == state ? dirty_1_54 : _GEN_10979; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12009 = 3'h3 == state ? dirty_1_55 : _GEN_10980; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12010 = 3'h3 == state ? dirty_1_56 : _GEN_10981; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12011 = 3'h3 == state ? dirty_1_57 : _GEN_10982; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12012 = 3'h3 == state ? dirty_1_58 : _GEN_10983; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12013 = 3'h3 == state ? dirty_1_59 : _GEN_10984; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12014 = 3'h3 == state ? dirty_1_60 : _GEN_10985; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12015 = 3'h3 == state ? dirty_1_61 : _GEN_10986; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12016 = 3'h3 == state ? dirty_1_62 : _GEN_10987; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12017 = 3'h3 == state ? dirty_1_63 : _GEN_10988; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12018 = 3'h3 == state ? dirty_1_64 : _GEN_10989; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12019 = 3'h3 == state ? dirty_1_65 : _GEN_10990; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12020 = 3'h3 == state ? dirty_1_66 : _GEN_10991; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12021 = 3'h3 == state ? dirty_1_67 : _GEN_10992; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12022 = 3'h3 == state ? dirty_1_68 : _GEN_10993; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12023 = 3'h3 == state ? dirty_1_69 : _GEN_10994; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12024 = 3'h3 == state ? dirty_1_70 : _GEN_10995; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12025 = 3'h3 == state ? dirty_1_71 : _GEN_10996; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12026 = 3'h3 == state ? dirty_1_72 : _GEN_10997; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12027 = 3'h3 == state ? dirty_1_73 : _GEN_10998; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12028 = 3'h3 == state ? dirty_1_74 : _GEN_10999; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12029 = 3'h3 == state ? dirty_1_75 : _GEN_11000; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12030 = 3'h3 == state ? dirty_1_76 : _GEN_11001; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12031 = 3'h3 == state ? dirty_1_77 : _GEN_11002; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12032 = 3'h3 == state ? dirty_1_78 : _GEN_11003; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12033 = 3'h3 == state ? dirty_1_79 : _GEN_11004; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12034 = 3'h3 == state ? dirty_1_80 : _GEN_11005; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12035 = 3'h3 == state ? dirty_1_81 : _GEN_11006; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12036 = 3'h3 == state ? dirty_1_82 : _GEN_11007; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12037 = 3'h3 == state ? dirty_1_83 : _GEN_11008; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12038 = 3'h3 == state ? dirty_1_84 : _GEN_11009; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12039 = 3'h3 == state ? dirty_1_85 : _GEN_11010; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12040 = 3'h3 == state ? dirty_1_86 : _GEN_11011; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12041 = 3'h3 == state ? dirty_1_87 : _GEN_11012; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12042 = 3'h3 == state ? dirty_1_88 : _GEN_11013; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12043 = 3'h3 == state ? dirty_1_89 : _GEN_11014; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12044 = 3'h3 == state ? dirty_1_90 : _GEN_11015; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12045 = 3'h3 == state ? dirty_1_91 : _GEN_11016; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12046 = 3'h3 == state ? dirty_1_92 : _GEN_11017; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12047 = 3'h3 == state ? dirty_1_93 : _GEN_11018; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12048 = 3'h3 == state ? dirty_1_94 : _GEN_11019; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12049 = 3'h3 == state ? dirty_1_95 : _GEN_11020; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12050 = 3'h3 == state ? dirty_1_96 : _GEN_11021; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12051 = 3'h3 == state ? dirty_1_97 : _GEN_11022; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12052 = 3'h3 == state ? dirty_1_98 : _GEN_11023; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12053 = 3'h3 == state ? dirty_1_99 : _GEN_11024; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12054 = 3'h3 == state ? dirty_1_100 : _GEN_11025; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12055 = 3'h3 == state ? dirty_1_101 : _GEN_11026; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12056 = 3'h3 == state ? dirty_1_102 : _GEN_11027; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12057 = 3'h3 == state ? dirty_1_103 : _GEN_11028; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12058 = 3'h3 == state ? dirty_1_104 : _GEN_11029; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12059 = 3'h3 == state ? dirty_1_105 : _GEN_11030; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12060 = 3'h3 == state ? dirty_1_106 : _GEN_11031; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12061 = 3'h3 == state ? dirty_1_107 : _GEN_11032; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12062 = 3'h3 == state ? dirty_1_108 : _GEN_11033; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12063 = 3'h3 == state ? dirty_1_109 : _GEN_11034; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12064 = 3'h3 == state ? dirty_1_110 : _GEN_11035; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12065 = 3'h3 == state ? dirty_1_111 : _GEN_11036; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12066 = 3'h3 == state ? dirty_1_112 : _GEN_11037; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12067 = 3'h3 == state ? dirty_1_113 : _GEN_11038; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12068 = 3'h3 == state ? dirty_1_114 : _GEN_11039; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12069 = 3'h3 == state ? dirty_1_115 : _GEN_11040; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12070 = 3'h3 == state ? dirty_1_116 : _GEN_11041; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12071 = 3'h3 == state ? dirty_1_117 : _GEN_11042; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12072 = 3'h3 == state ? dirty_1_118 : _GEN_11043; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12073 = 3'h3 == state ? dirty_1_119 : _GEN_11044; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12074 = 3'h3 == state ? dirty_1_120 : _GEN_11045; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12075 = 3'h3 == state ? dirty_1_121 : _GEN_11046; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12076 = 3'h3 == state ? dirty_1_122 : _GEN_11047; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12077 = 3'h3 == state ? dirty_1_123 : _GEN_11048; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12078 = 3'h3 == state ? dirty_1_124 : _GEN_11049; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12079 = 3'h3 == state ? dirty_1_125 : _GEN_11050; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12080 = 3'h3 == state ? dirty_1_126 : _GEN_11051; // @[d_cache.scala 64:18 25:26]
  wire  _GEN_12081 = 3'h3 == state ? dirty_1_127 : _GEN_11052; // @[d_cache.scala 64:18 25:26]
  wire [38:0] _GEN_13110 = 3'h2 == state ? {{7'd0}, write_back_addr} : _GEN_11825; // @[d_cache.scala 64:18 30:34]
  wire [38:0] _GEN_14139 = 3'h1 == state ? {{7'd0}, write_back_addr} : _GEN_13110; // @[d_cache.scala 64:18 30:34]
  wire [38:0] _GEN_15168 = 3'h0 == state ? {{7'd0}, write_back_addr} : _GEN_14139; // @[d_cache.scala 64:18 30:34]
  wire [63:0] _GEN_15169 = way1_hit ? _GEN_4497 : 64'h0; // @[d_cache.scala 212:33 213:33 220:33]
  wire [63:0] _GEN_15173 = way0_hit ? _GEN_2957 : _GEN_15169; // @[d_cache.scala 205:23 206:33]
  wire  _GEN_15175 = way0_hit | way1_hit; // @[d_cache.scala 205:23 208:34]
  wire  _GEN_15177 = way1_hit ? 1'h0 : 1'h1; // @[d_cache.scala 244:33 246:35 253:35]
  wire  _GEN_15178 = way0_hit ? 1'h0 : _GEN_15177; // @[d_cache.scala 237:23 239:35]
  wire  _T_36 = state == 3'h3; // @[d_cache.scala 259:21]
  wire  _T_39 = state == 3'h6; // @[d_cache.scala 308:21]
  wire [31:0] _GEN_15181 = state == 3'h6 ? 32'h0 : io_from_lsu_araddr; // @[d_cache.scala 308:35 316:26 332:26]
  wire  _GEN_15182 = state == 3'h6 ? 1'h0 : io_from_lsu_rready; // @[d_cache.scala 308:35 317:26 333:26]
  wire [31:0] _GEN_15183 = state == 3'h6 ? write_back_addr : 32'h0; // @[d_cache.scala 308:35 318:26 334:26]
  wire [63:0] _GEN_15184 = state == 3'h6 ? write_back_data : 64'h0; // @[d_cache.scala 308:35 320:25 336:25]
  wire [31:0] _GEN_15185 = state == 3'h6 ? 32'hffffffff : 32'h0; // @[d_cache.scala 308:35 321:25 337:25]
  wire  _GEN_15187 = state == 3'h5 | _T_39; // @[d_cache.scala 292:31 294:27]
  wire [31:0] _GEN_15188 = state == 3'h5 ? io_from_lsu_araddr : _GEN_15181; // @[d_cache.scala 292:31 300:26]
  wire  _GEN_15189 = state == 3'h5 ? io_from_lsu_rready : _GEN_15182; // @[d_cache.scala 292:31 301:26]
  wire [31:0] _GEN_15190 = state == 3'h5 ? 32'h0 : _GEN_15183; // @[d_cache.scala 292:31 302:26]
  wire  _GEN_15191 = state == 3'h5 ? 1'h0 : _T_39; // @[d_cache.scala 292:31 303:27]
  wire [63:0] _GEN_15192 = state == 3'h5 ? 64'h0 : _GEN_15184; // @[d_cache.scala 292:31 304:25]
  wire [31:0] _GEN_15193 = state == 3'h5 ? 32'h0 : _GEN_15185; // @[d_cache.scala 292:31 305:25]
  wire  _GEN_15195 = state == 3'h4 | _GEN_15187; // @[d_cache.scala 275:31 277:27]
  wire  _GEN_15196 = state == 3'h4 & io_from_axi_wready; // @[d_cache.scala 275:31 279:26]
  wire  _GEN_15197 = state == 3'h4 & io_from_axi_bvalid; // @[d_cache.scala 275:31 280:26]
  wire  _GEN_15198 = state == 3'h4 & io_from_axi_awready; // @[d_cache.scala 275:31 281:27]
  wire [31:0] _GEN_15199 = state == 3'h4 ? 32'h0 : _GEN_15188; // @[d_cache.scala 275:31 283:26]
  wire  _GEN_15200 = state == 3'h4 ? io_from_lsu_rready : _GEN_15189; // @[d_cache.scala 275:31 284:26]
  wire [31:0] _GEN_15201 = state == 3'h4 ? io_from_lsu_awaddr : _GEN_15190; // @[d_cache.scala 275:31 285:26]
  wire  _GEN_15202 = state == 3'h4 ? io_from_lsu_awvalid : _GEN_15191; // @[d_cache.scala 275:31 286:27]
  wire [63:0] _GEN_15203 = state == 3'h4 ? {{32'd0}, io_from_lsu_wdata} : _GEN_15192; // @[d_cache.scala 275:31 287:25]
  wire [31:0] _GEN_15204 = state == 3'h4 ? {{24'd0}, io_from_lsu_wstrb} : _GEN_15193; // @[d_cache.scala 275:31 288:25]
  wire  _GEN_15205 = state == 3'h4 ? io_from_lsu_wvalid : _GEN_15191; // @[d_cache.scala 275:31 289:26]
  wire  _GEN_15206 = state == 3'h4 ? io_from_lsu_bready : _GEN_15191; // @[d_cache.scala 275:31 290:26]
  wire  _GEN_15208 = state == 3'h3 | _GEN_15195; // @[d_cache.scala 259:31 261:27]
  wire  _GEN_15209 = state == 3'h3 ? 1'h0 : _GEN_15196; // @[d_cache.scala 259:31 263:26]
  wire  _GEN_15210 = state == 3'h3 ? 1'h0 : _GEN_15197; // @[d_cache.scala 259:31 264:26]
  wire  _GEN_15211 = state == 3'h3 ? 1'h0 : _GEN_15198; // @[d_cache.scala 259:31 265:27]
  wire [31:0] _GEN_15213 = state == 3'h3 ? io_from_lsu_araddr : _GEN_15199; // @[d_cache.scala 259:31 267:26]
  wire  _GEN_15214 = state == 3'h3 ? io_from_lsu_rready : _GEN_15200; // @[d_cache.scala 259:31 268:26]
  wire [31:0] _GEN_15215 = state == 3'h3 ? 32'h0 : _GEN_15201; // @[d_cache.scala 259:31 269:26]
  wire  _GEN_15216 = state == 3'h3 ? 1'h0 : _GEN_15202; // @[d_cache.scala 259:31 270:27]
  wire [63:0] _GEN_15217 = state == 3'h3 ? 64'h0 : _GEN_15203; // @[d_cache.scala 259:31 271:25]
  wire [31:0] _GEN_15218 = state == 3'h3 ? 32'h0 : _GEN_15204; // @[d_cache.scala 259:31 272:25]
  wire  _GEN_15219 = state == 3'h3 ? 1'h0 : _GEN_15205; // @[d_cache.scala 259:31 273:26]
  wire  _GEN_15220 = state == 3'h3 ? 1'h0 : _GEN_15206; // @[d_cache.scala 259:31 274:26]
  wire  _GEN_15221 = state == 3'h2 ? 1'h0 : _T_36; // @[d_cache.scala 227:33 228:27]
  wire [31:0] _GEN_15222 = state == 3'h2 ? io_from_lsu_araddr : _GEN_15213; // @[d_cache.scala 227:33 229:26]
  wire  _GEN_15223 = state == 3'h2 ? 1'h0 : _GEN_15214; // @[d_cache.scala 227:33 230:26]
  wire [31:0] _GEN_15224 = state == 3'h2 ? 32'h0 : _GEN_15215; // @[d_cache.scala 227:33 231:26]
  wire  _GEN_15225 = state == 3'h2 ? 1'h0 : _GEN_15216; // @[d_cache.scala 227:33 232:27]
  wire [63:0] _GEN_15226 = state == 3'h2 ? 64'h0 : _GEN_15217; // @[d_cache.scala 227:33 233:25]
  wire [31:0] _GEN_15227 = state == 3'h2 ? 32'h0 : _GEN_15218; // @[d_cache.scala 227:33 234:25]
  wire  _GEN_15228 = state == 3'h2 ? 1'h0 : _GEN_15219; // @[d_cache.scala 227:33 235:26]
  wire  _GEN_15229 = state == 3'h2 ? 1'h0 : _GEN_15220; // @[d_cache.scala 227:33 236:26]
  wire  _GEN_15231 = state == 3'h2 ? _GEN_15178 : _GEN_15208; // @[d_cache.scala 227:33]
  wire  _GEN_15232 = state == 3'h2 ? _GEN_15175 : _GEN_15209; // @[d_cache.scala 227:33]
  wire  _GEN_15233 = state == 3'h2 ? _GEN_15175 : _GEN_15211; // @[d_cache.scala 227:33]
  wire  _GEN_15234 = state == 3'h2 ? _GEN_15175 : _GEN_15210; // @[d_cache.scala 227:33]
  wire  _GEN_15235 = state == 3'h1 ? 1'h0 : _GEN_15221; // @[d_cache.scala 195:33 196:27]
  wire [31:0] _GEN_15236 = state == 3'h1 ? io_from_lsu_araddr : _GEN_15222; // @[d_cache.scala 195:33 197:26]
  wire  _GEN_15237 = state == 3'h1 ? io_from_lsu_rready : _GEN_15223; // @[d_cache.scala 195:33 198:26]
  wire [31:0] _GEN_15238 = state == 3'h1 ? 32'h0 : _GEN_15224; // @[d_cache.scala 195:33 199:26]
  wire  _GEN_15239 = state == 3'h1 ? 1'h0 : _GEN_15225; // @[d_cache.scala 195:33 200:27]
  wire [63:0] _GEN_15240 = state == 3'h1 ? 64'h0 : _GEN_15226; // @[d_cache.scala 195:33 201:25]
  wire [31:0] _GEN_15241 = state == 3'h1 ? 32'h0 : _GEN_15227; // @[d_cache.scala 195:33 202:25]
  wire  _GEN_15242 = state == 3'h1 ? 1'h0 : _GEN_15228; // @[d_cache.scala 195:33 203:26]
  wire  _GEN_15243 = state == 3'h1 ? io_from_lsu_bready : _GEN_15229; // @[d_cache.scala 195:33 204:26]
  wire [63:0] _GEN_15244 = state == 3'h1 ? _GEN_15173 : 64'h0; // @[d_cache.scala 195:33]
  wire  _GEN_15245 = state == 3'h1 | _GEN_15231; // @[d_cache.scala 195:33]
  wire  _GEN_15246 = state == 3'h1 & _GEN_15175; // @[d_cache.scala 195:33]
  wire  _GEN_15247 = state == 3'h1 ? 1'h0 : _GEN_15232; // @[d_cache.scala 195:33]
  wire  _GEN_15248 = state == 3'h1 ? 1'h0 : _GEN_15233; // @[d_cache.scala 195:33]
  wire  _GEN_15249 = state == 3'h1 ? 1'h0 : _GEN_15234; // @[d_cache.scala 195:33]
  wire [63:0] _GEN_15261 = state == 3'h0 ? 64'h0 : _GEN_15240; // @[d_cache.scala 179:23 191:25]
  wire [31:0] _GEN_15262 = state == 3'h0 ? 32'h0 : _GEN_15241; // @[d_cache.scala 179:23 192:25]
  wire [38:0] _GEN_16293 = reset ? 39'h0 : _GEN_15168; // @[d_cache.scala 30:{34,34}]
  wire  _GEN_16295 = ~_T_16 & _T_17; // @[d_cache.scala 76:27]
  assign io_to_lsu_arready = state == 3'h0 ? io_from_axi_arready : _GEN_15245; // @[d_cache.scala 179:23 181:27]
  assign io_to_lsu_rdata = state == 3'h0 ? 64'h0 : _GEN_15244; // @[d_cache.scala 179:23 180:25]
  assign io_to_lsu_rvalid = state == 3'h0 ? 1'h0 : _GEN_15246; // @[d_cache.scala 179:23 182:26]
  assign io_to_lsu_awready = state == 3'h0 ? io_from_axi_awready : _GEN_15248; // @[d_cache.scala 179:23 185:27]
  assign io_to_lsu_wready = state == 3'h0 ? 1'h0 : _GEN_15247; // @[d_cache.scala 179:23 183:26]
  assign io_to_lsu_bvalid = state == 3'h0 ? 1'h0 : _GEN_15249; // @[d_cache.scala 179:23 184:26]
  assign io_to_axi_araddr = state == 3'h0 ? io_from_lsu_araddr : _GEN_15236; // @[d_cache.scala 179:23 187:26]
  assign io_to_axi_arvalid = state == 3'h0 ? 1'h0 : _GEN_15235; // @[d_cache.scala 179:23 186:27]
  assign io_to_axi_rready = state == 3'h0 ? io_from_lsu_rready : _GEN_15237; // @[d_cache.scala 179:23 188:26]
  assign io_to_axi_awaddr = state == 3'h0 ? 32'h0 : _GEN_15238; // @[d_cache.scala 179:23 189:26]
  assign io_to_axi_awvalid = state == 3'h0 ? 1'h0 : _GEN_15239; // @[d_cache.scala 179:23 190:27]
  assign io_to_axi_wdata = _GEN_15261[31:0];
  assign io_to_axi_wstrb = _GEN_15262[7:0];
  assign io_to_axi_wvalid = state == 3'h0 ? 1'h0 : _GEN_15242; // @[d_cache.scala 179:23 193:26]
  assign io_to_axi_bready = state == 3'h0 ? io_from_lsu_bready : _GEN_15243; // @[d_cache.scala 179:23 194:26]
  always @(posedge clock) begin
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_0 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_0 <= _GEN_1547;
        end else begin
          ram_0_0 <= _GEN_11055;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_1 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_1 <= _GEN_1548;
        end else begin
          ram_0_1 <= _GEN_11056;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_2 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_2 <= _GEN_1549;
        end else begin
          ram_0_2 <= _GEN_11057;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_3 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_3 <= _GEN_1550;
        end else begin
          ram_0_3 <= _GEN_11058;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_4 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_4 <= _GEN_1551;
        end else begin
          ram_0_4 <= _GEN_11059;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_5 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_5 <= _GEN_1552;
        end else begin
          ram_0_5 <= _GEN_11060;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_6 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_6 <= _GEN_1553;
        end else begin
          ram_0_6 <= _GEN_11061;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_7 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_7 <= _GEN_1554;
        end else begin
          ram_0_7 <= _GEN_11062;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_8 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_8 <= _GEN_1555;
        end else begin
          ram_0_8 <= _GEN_11063;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_9 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_9 <= _GEN_1556;
        end else begin
          ram_0_9 <= _GEN_11064;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_10 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_10 <= _GEN_1557;
        end else begin
          ram_0_10 <= _GEN_11065;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_11 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_11 <= _GEN_1558;
        end else begin
          ram_0_11 <= _GEN_11066;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_12 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_12 <= _GEN_1559;
        end else begin
          ram_0_12 <= _GEN_11067;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_13 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_13 <= _GEN_1560;
        end else begin
          ram_0_13 <= _GEN_11068;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_14 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_14 <= _GEN_1561;
        end else begin
          ram_0_14 <= _GEN_11069;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_15 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_15 <= _GEN_1562;
        end else begin
          ram_0_15 <= _GEN_11070;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_16 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_16 <= _GEN_1563;
        end else begin
          ram_0_16 <= _GEN_11071;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_17 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_17 <= _GEN_1564;
        end else begin
          ram_0_17 <= _GEN_11072;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_18 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_18 <= _GEN_1565;
        end else begin
          ram_0_18 <= _GEN_11073;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_19 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_19 <= _GEN_1566;
        end else begin
          ram_0_19 <= _GEN_11074;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_20 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_20 <= _GEN_1567;
        end else begin
          ram_0_20 <= _GEN_11075;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_21 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_21 <= _GEN_1568;
        end else begin
          ram_0_21 <= _GEN_11076;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_22 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_22 <= _GEN_1569;
        end else begin
          ram_0_22 <= _GEN_11077;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_23 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_23 <= _GEN_1570;
        end else begin
          ram_0_23 <= _GEN_11078;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_24 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_24 <= _GEN_1571;
        end else begin
          ram_0_24 <= _GEN_11079;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_25 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_25 <= _GEN_1572;
        end else begin
          ram_0_25 <= _GEN_11080;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_26 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_26 <= _GEN_1573;
        end else begin
          ram_0_26 <= _GEN_11081;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_27 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_27 <= _GEN_1574;
        end else begin
          ram_0_27 <= _GEN_11082;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_28 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_28 <= _GEN_1575;
        end else begin
          ram_0_28 <= _GEN_11083;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_29 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_29 <= _GEN_1576;
        end else begin
          ram_0_29 <= _GEN_11084;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_30 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_30 <= _GEN_1577;
        end else begin
          ram_0_30 <= _GEN_11085;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_31 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_31 <= _GEN_1578;
        end else begin
          ram_0_31 <= _GEN_11086;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_32 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_32 <= _GEN_1579;
        end else begin
          ram_0_32 <= _GEN_11087;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_33 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_33 <= _GEN_1580;
        end else begin
          ram_0_33 <= _GEN_11088;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_34 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_34 <= _GEN_1581;
        end else begin
          ram_0_34 <= _GEN_11089;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_35 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_35 <= _GEN_1582;
        end else begin
          ram_0_35 <= _GEN_11090;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_36 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_36 <= _GEN_1583;
        end else begin
          ram_0_36 <= _GEN_11091;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_37 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_37 <= _GEN_1584;
        end else begin
          ram_0_37 <= _GEN_11092;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_38 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_38 <= _GEN_1585;
        end else begin
          ram_0_38 <= _GEN_11093;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_39 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_39 <= _GEN_1586;
        end else begin
          ram_0_39 <= _GEN_11094;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_40 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_40 <= _GEN_1587;
        end else begin
          ram_0_40 <= _GEN_11095;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_41 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_41 <= _GEN_1588;
        end else begin
          ram_0_41 <= _GEN_11096;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_42 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_42 <= _GEN_1589;
        end else begin
          ram_0_42 <= _GEN_11097;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_43 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_43 <= _GEN_1590;
        end else begin
          ram_0_43 <= _GEN_11098;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_44 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_44 <= _GEN_1591;
        end else begin
          ram_0_44 <= _GEN_11099;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_45 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_45 <= _GEN_1592;
        end else begin
          ram_0_45 <= _GEN_11100;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_46 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_46 <= _GEN_1593;
        end else begin
          ram_0_46 <= _GEN_11101;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_47 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_47 <= _GEN_1594;
        end else begin
          ram_0_47 <= _GEN_11102;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_48 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_48 <= _GEN_1595;
        end else begin
          ram_0_48 <= _GEN_11103;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_49 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_49 <= _GEN_1596;
        end else begin
          ram_0_49 <= _GEN_11104;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_50 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_50 <= _GEN_1597;
        end else begin
          ram_0_50 <= _GEN_11105;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_51 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_51 <= _GEN_1598;
        end else begin
          ram_0_51 <= _GEN_11106;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_52 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_52 <= _GEN_1599;
        end else begin
          ram_0_52 <= _GEN_11107;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_53 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_53 <= _GEN_1600;
        end else begin
          ram_0_53 <= _GEN_11108;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_54 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_54 <= _GEN_1601;
        end else begin
          ram_0_54 <= _GEN_11109;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_55 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_55 <= _GEN_1602;
        end else begin
          ram_0_55 <= _GEN_11110;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_56 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_56 <= _GEN_1603;
        end else begin
          ram_0_56 <= _GEN_11111;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_57 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_57 <= _GEN_1604;
        end else begin
          ram_0_57 <= _GEN_11112;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_58 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_58 <= _GEN_1605;
        end else begin
          ram_0_58 <= _GEN_11113;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_59 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_59 <= _GEN_1606;
        end else begin
          ram_0_59 <= _GEN_11114;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_60 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_60 <= _GEN_1607;
        end else begin
          ram_0_60 <= _GEN_11115;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_61 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_61 <= _GEN_1608;
        end else begin
          ram_0_61 <= _GEN_11116;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_62 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_62 <= _GEN_1609;
        end else begin
          ram_0_62 <= _GEN_11117;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_63 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_63 <= _GEN_1610;
        end else begin
          ram_0_63 <= _GEN_11118;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_64 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_64 <= _GEN_1611;
        end else begin
          ram_0_64 <= _GEN_11119;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_65 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_65 <= _GEN_1612;
        end else begin
          ram_0_65 <= _GEN_11120;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_66 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_66 <= _GEN_1613;
        end else begin
          ram_0_66 <= _GEN_11121;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_67 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_67 <= _GEN_1614;
        end else begin
          ram_0_67 <= _GEN_11122;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_68 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_68 <= _GEN_1615;
        end else begin
          ram_0_68 <= _GEN_11123;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_69 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_69 <= _GEN_1616;
        end else begin
          ram_0_69 <= _GEN_11124;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_70 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_70 <= _GEN_1617;
        end else begin
          ram_0_70 <= _GEN_11125;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_71 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_71 <= _GEN_1618;
        end else begin
          ram_0_71 <= _GEN_11126;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_72 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_72 <= _GEN_1619;
        end else begin
          ram_0_72 <= _GEN_11127;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_73 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_73 <= _GEN_1620;
        end else begin
          ram_0_73 <= _GEN_11128;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_74 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_74 <= _GEN_1621;
        end else begin
          ram_0_74 <= _GEN_11129;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_75 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_75 <= _GEN_1622;
        end else begin
          ram_0_75 <= _GEN_11130;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_76 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_76 <= _GEN_1623;
        end else begin
          ram_0_76 <= _GEN_11131;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_77 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_77 <= _GEN_1624;
        end else begin
          ram_0_77 <= _GEN_11132;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_78 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_78 <= _GEN_1625;
        end else begin
          ram_0_78 <= _GEN_11133;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_79 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_79 <= _GEN_1626;
        end else begin
          ram_0_79 <= _GEN_11134;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_80 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_80 <= _GEN_1627;
        end else begin
          ram_0_80 <= _GEN_11135;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_81 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_81 <= _GEN_1628;
        end else begin
          ram_0_81 <= _GEN_11136;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_82 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_82 <= _GEN_1629;
        end else begin
          ram_0_82 <= _GEN_11137;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_83 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_83 <= _GEN_1630;
        end else begin
          ram_0_83 <= _GEN_11138;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_84 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_84 <= _GEN_1631;
        end else begin
          ram_0_84 <= _GEN_11139;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_85 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_85 <= _GEN_1632;
        end else begin
          ram_0_85 <= _GEN_11140;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_86 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_86 <= _GEN_1633;
        end else begin
          ram_0_86 <= _GEN_11141;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_87 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_87 <= _GEN_1634;
        end else begin
          ram_0_87 <= _GEN_11142;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_88 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_88 <= _GEN_1635;
        end else begin
          ram_0_88 <= _GEN_11143;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_89 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_89 <= _GEN_1636;
        end else begin
          ram_0_89 <= _GEN_11144;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_90 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_90 <= _GEN_1637;
        end else begin
          ram_0_90 <= _GEN_11145;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_91 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_91 <= _GEN_1638;
        end else begin
          ram_0_91 <= _GEN_11146;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_92 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_92 <= _GEN_1639;
        end else begin
          ram_0_92 <= _GEN_11147;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_93 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_93 <= _GEN_1640;
        end else begin
          ram_0_93 <= _GEN_11148;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_94 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_94 <= _GEN_1641;
        end else begin
          ram_0_94 <= _GEN_11149;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_95 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_95 <= _GEN_1642;
        end else begin
          ram_0_95 <= _GEN_11150;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_96 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_96 <= _GEN_1643;
        end else begin
          ram_0_96 <= _GEN_11151;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_97 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_97 <= _GEN_1644;
        end else begin
          ram_0_97 <= _GEN_11152;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_98 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_98 <= _GEN_1645;
        end else begin
          ram_0_98 <= _GEN_11153;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_99 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_99 <= _GEN_1646;
        end else begin
          ram_0_99 <= _GEN_11154;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_100 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_100 <= _GEN_1647;
        end else begin
          ram_0_100 <= _GEN_11155;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_101 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_101 <= _GEN_1648;
        end else begin
          ram_0_101 <= _GEN_11156;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_102 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_102 <= _GEN_1649;
        end else begin
          ram_0_102 <= _GEN_11157;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_103 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_103 <= _GEN_1650;
        end else begin
          ram_0_103 <= _GEN_11158;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_104 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_104 <= _GEN_1651;
        end else begin
          ram_0_104 <= _GEN_11159;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_105 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_105 <= _GEN_1652;
        end else begin
          ram_0_105 <= _GEN_11160;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_106 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_106 <= _GEN_1653;
        end else begin
          ram_0_106 <= _GEN_11161;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_107 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_107 <= _GEN_1654;
        end else begin
          ram_0_107 <= _GEN_11162;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_108 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_108 <= _GEN_1655;
        end else begin
          ram_0_108 <= _GEN_11163;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_109 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_109 <= _GEN_1656;
        end else begin
          ram_0_109 <= _GEN_11164;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_110 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_110 <= _GEN_1657;
        end else begin
          ram_0_110 <= _GEN_11165;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_111 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_111 <= _GEN_1658;
        end else begin
          ram_0_111 <= _GEN_11166;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_112 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_112 <= _GEN_1659;
        end else begin
          ram_0_112 <= _GEN_11167;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_113 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_113 <= _GEN_1660;
        end else begin
          ram_0_113 <= _GEN_11168;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_114 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_114 <= _GEN_1661;
        end else begin
          ram_0_114 <= _GEN_11169;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_115 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_115 <= _GEN_1662;
        end else begin
          ram_0_115 <= _GEN_11170;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_116 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_116 <= _GEN_1663;
        end else begin
          ram_0_116 <= _GEN_11171;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_117 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_117 <= _GEN_1664;
        end else begin
          ram_0_117 <= _GEN_11172;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_118 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_118 <= _GEN_1665;
        end else begin
          ram_0_118 <= _GEN_11173;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_119 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_119 <= _GEN_1666;
        end else begin
          ram_0_119 <= _GEN_11174;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_120 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_120 <= _GEN_1667;
        end else begin
          ram_0_120 <= _GEN_11175;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_121 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_121 <= _GEN_1668;
        end else begin
          ram_0_121 <= _GEN_11176;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_122 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_122 <= _GEN_1669;
        end else begin
          ram_0_122 <= _GEN_11177;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_123 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_123 <= _GEN_1670;
        end else begin
          ram_0_123 <= _GEN_11178;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_124 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_124 <= _GEN_1671;
        end else begin
          ram_0_124 <= _GEN_11179;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_125 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_125 <= _GEN_1672;
        end else begin
          ram_0_125 <= _GEN_11180;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_126 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_126 <= _GEN_1673;
        end else begin
          ram_0_126 <= _GEN_11181;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_127 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_0_127 <= _GEN_1674;
        end else begin
          ram_0_127 <= _GEN_11182;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_0 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_0 <= _GEN_1803;
        end else begin
          ram_1_0 <= _GEN_11440;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_1 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_1 <= _GEN_1804;
        end else begin
          ram_1_1 <= _GEN_11441;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_2 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_2 <= _GEN_1805;
        end else begin
          ram_1_2 <= _GEN_11442;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_3 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_3 <= _GEN_1806;
        end else begin
          ram_1_3 <= _GEN_11443;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_4 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_4 <= _GEN_1807;
        end else begin
          ram_1_4 <= _GEN_11444;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_5 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_5 <= _GEN_1808;
        end else begin
          ram_1_5 <= _GEN_11445;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_6 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_6 <= _GEN_1809;
        end else begin
          ram_1_6 <= _GEN_11446;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_7 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_7 <= _GEN_1810;
        end else begin
          ram_1_7 <= _GEN_11447;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_8 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_8 <= _GEN_1811;
        end else begin
          ram_1_8 <= _GEN_11448;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_9 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_9 <= _GEN_1812;
        end else begin
          ram_1_9 <= _GEN_11449;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_10 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_10 <= _GEN_1813;
        end else begin
          ram_1_10 <= _GEN_11450;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_11 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_11 <= _GEN_1814;
        end else begin
          ram_1_11 <= _GEN_11451;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_12 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_12 <= _GEN_1815;
        end else begin
          ram_1_12 <= _GEN_11452;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_13 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_13 <= _GEN_1816;
        end else begin
          ram_1_13 <= _GEN_11453;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_14 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_14 <= _GEN_1817;
        end else begin
          ram_1_14 <= _GEN_11454;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_15 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_15 <= _GEN_1818;
        end else begin
          ram_1_15 <= _GEN_11455;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_16 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_16 <= _GEN_1819;
        end else begin
          ram_1_16 <= _GEN_11456;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_17 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_17 <= _GEN_1820;
        end else begin
          ram_1_17 <= _GEN_11457;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_18 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_18 <= _GEN_1821;
        end else begin
          ram_1_18 <= _GEN_11458;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_19 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_19 <= _GEN_1822;
        end else begin
          ram_1_19 <= _GEN_11459;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_20 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_20 <= _GEN_1823;
        end else begin
          ram_1_20 <= _GEN_11460;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_21 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_21 <= _GEN_1824;
        end else begin
          ram_1_21 <= _GEN_11461;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_22 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_22 <= _GEN_1825;
        end else begin
          ram_1_22 <= _GEN_11462;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_23 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_23 <= _GEN_1826;
        end else begin
          ram_1_23 <= _GEN_11463;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_24 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_24 <= _GEN_1827;
        end else begin
          ram_1_24 <= _GEN_11464;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_25 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_25 <= _GEN_1828;
        end else begin
          ram_1_25 <= _GEN_11465;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_26 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_26 <= _GEN_1829;
        end else begin
          ram_1_26 <= _GEN_11466;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_27 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_27 <= _GEN_1830;
        end else begin
          ram_1_27 <= _GEN_11467;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_28 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_28 <= _GEN_1831;
        end else begin
          ram_1_28 <= _GEN_11468;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_29 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_29 <= _GEN_1832;
        end else begin
          ram_1_29 <= _GEN_11469;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_30 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_30 <= _GEN_1833;
        end else begin
          ram_1_30 <= _GEN_11470;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_31 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_31 <= _GEN_1834;
        end else begin
          ram_1_31 <= _GEN_11471;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_32 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_32 <= _GEN_1835;
        end else begin
          ram_1_32 <= _GEN_11472;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_33 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_33 <= _GEN_1836;
        end else begin
          ram_1_33 <= _GEN_11473;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_34 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_34 <= _GEN_1837;
        end else begin
          ram_1_34 <= _GEN_11474;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_35 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_35 <= _GEN_1838;
        end else begin
          ram_1_35 <= _GEN_11475;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_36 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_36 <= _GEN_1839;
        end else begin
          ram_1_36 <= _GEN_11476;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_37 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_37 <= _GEN_1840;
        end else begin
          ram_1_37 <= _GEN_11477;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_38 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_38 <= _GEN_1841;
        end else begin
          ram_1_38 <= _GEN_11478;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_39 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_39 <= _GEN_1842;
        end else begin
          ram_1_39 <= _GEN_11479;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_40 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_40 <= _GEN_1843;
        end else begin
          ram_1_40 <= _GEN_11480;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_41 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_41 <= _GEN_1844;
        end else begin
          ram_1_41 <= _GEN_11481;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_42 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_42 <= _GEN_1845;
        end else begin
          ram_1_42 <= _GEN_11482;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_43 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_43 <= _GEN_1846;
        end else begin
          ram_1_43 <= _GEN_11483;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_44 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_44 <= _GEN_1847;
        end else begin
          ram_1_44 <= _GEN_11484;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_45 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_45 <= _GEN_1848;
        end else begin
          ram_1_45 <= _GEN_11485;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_46 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_46 <= _GEN_1849;
        end else begin
          ram_1_46 <= _GEN_11486;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_47 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_47 <= _GEN_1850;
        end else begin
          ram_1_47 <= _GEN_11487;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_48 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_48 <= _GEN_1851;
        end else begin
          ram_1_48 <= _GEN_11488;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_49 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_49 <= _GEN_1852;
        end else begin
          ram_1_49 <= _GEN_11489;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_50 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_50 <= _GEN_1853;
        end else begin
          ram_1_50 <= _GEN_11490;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_51 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_51 <= _GEN_1854;
        end else begin
          ram_1_51 <= _GEN_11491;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_52 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_52 <= _GEN_1855;
        end else begin
          ram_1_52 <= _GEN_11492;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_53 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_53 <= _GEN_1856;
        end else begin
          ram_1_53 <= _GEN_11493;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_54 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_54 <= _GEN_1857;
        end else begin
          ram_1_54 <= _GEN_11494;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_55 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_55 <= _GEN_1858;
        end else begin
          ram_1_55 <= _GEN_11495;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_56 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_56 <= _GEN_1859;
        end else begin
          ram_1_56 <= _GEN_11496;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_57 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_57 <= _GEN_1860;
        end else begin
          ram_1_57 <= _GEN_11497;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_58 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_58 <= _GEN_1861;
        end else begin
          ram_1_58 <= _GEN_11498;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_59 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_59 <= _GEN_1862;
        end else begin
          ram_1_59 <= _GEN_11499;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_60 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_60 <= _GEN_1863;
        end else begin
          ram_1_60 <= _GEN_11500;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_61 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_61 <= _GEN_1864;
        end else begin
          ram_1_61 <= _GEN_11501;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_62 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_62 <= _GEN_1865;
        end else begin
          ram_1_62 <= _GEN_11502;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_63 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_63 <= _GEN_1866;
        end else begin
          ram_1_63 <= _GEN_11503;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_64 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_64 <= _GEN_1867;
        end else begin
          ram_1_64 <= _GEN_11504;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_65 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_65 <= _GEN_1868;
        end else begin
          ram_1_65 <= _GEN_11505;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_66 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_66 <= _GEN_1869;
        end else begin
          ram_1_66 <= _GEN_11506;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_67 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_67 <= _GEN_1870;
        end else begin
          ram_1_67 <= _GEN_11507;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_68 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_68 <= _GEN_1871;
        end else begin
          ram_1_68 <= _GEN_11508;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_69 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_69 <= _GEN_1872;
        end else begin
          ram_1_69 <= _GEN_11509;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_70 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_70 <= _GEN_1873;
        end else begin
          ram_1_70 <= _GEN_11510;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_71 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_71 <= _GEN_1874;
        end else begin
          ram_1_71 <= _GEN_11511;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_72 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_72 <= _GEN_1875;
        end else begin
          ram_1_72 <= _GEN_11512;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_73 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_73 <= _GEN_1876;
        end else begin
          ram_1_73 <= _GEN_11513;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_74 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_74 <= _GEN_1877;
        end else begin
          ram_1_74 <= _GEN_11514;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_75 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_75 <= _GEN_1878;
        end else begin
          ram_1_75 <= _GEN_11515;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_76 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_76 <= _GEN_1879;
        end else begin
          ram_1_76 <= _GEN_11516;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_77 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_77 <= _GEN_1880;
        end else begin
          ram_1_77 <= _GEN_11517;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_78 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_78 <= _GEN_1881;
        end else begin
          ram_1_78 <= _GEN_11518;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_79 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_79 <= _GEN_1882;
        end else begin
          ram_1_79 <= _GEN_11519;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_80 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_80 <= _GEN_1883;
        end else begin
          ram_1_80 <= _GEN_11520;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_81 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_81 <= _GEN_1884;
        end else begin
          ram_1_81 <= _GEN_11521;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_82 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_82 <= _GEN_1885;
        end else begin
          ram_1_82 <= _GEN_11522;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_83 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_83 <= _GEN_1886;
        end else begin
          ram_1_83 <= _GEN_11523;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_84 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_84 <= _GEN_1887;
        end else begin
          ram_1_84 <= _GEN_11524;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_85 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_85 <= _GEN_1888;
        end else begin
          ram_1_85 <= _GEN_11525;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_86 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_86 <= _GEN_1889;
        end else begin
          ram_1_86 <= _GEN_11526;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_87 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_87 <= _GEN_1890;
        end else begin
          ram_1_87 <= _GEN_11527;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_88 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_88 <= _GEN_1891;
        end else begin
          ram_1_88 <= _GEN_11528;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_89 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_89 <= _GEN_1892;
        end else begin
          ram_1_89 <= _GEN_11529;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_90 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_90 <= _GEN_1893;
        end else begin
          ram_1_90 <= _GEN_11530;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_91 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_91 <= _GEN_1894;
        end else begin
          ram_1_91 <= _GEN_11531;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_92 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_92 <= _GEN_1895;
        end else begin
          ram_1_92 <= _GEN_11532;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_93 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_93 <= _GEN_1896;
        end else begin
          ram_1_93 <= _GEN_11533;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_94 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_94 <= _GEN_1897;
        end else begin
          ram_1_94 <= _GEN_11534;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_95 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_95 <= _GEN_1898;
        end else begin
          ram_1_95 <= _GEN_11535;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_96 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_96 <= _GEN_1899;
        end else begin
          ram_1_96 <= _GEN_11536;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_97 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_97 <= _GEN_1900;
        end else begin
          ram_1_97 <= _GEN_11537;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_98 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_98 <= _GEN_1901;
        end else begin
          ram_1_98 <= _GEN_11538;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_99 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_99 <= _GEN_1902;
        end else begin
          ram_1_99 <= _GEN_11539;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_100 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_100 <= _GEN_1903;
        end else begin
          ram_1_100 <= _GEN_11540;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_101 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_101 <= _GEN_1904;
        end else begin
          ram_1_101 <= _GEN_11541;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_102 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_102 <= _GEN_1905;
        end else begin
          ram_1_102 <= _GEN_11542;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_103 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_103 <= _GEN_1906;
        end else begin
          ram_1_103 <= _GEN_11543;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_104 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_104 <= _GEN_1907;
        end else begin
          ram_1_104 <= _GEN_11544;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_105 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_105 <= _GEN_1908;
        end else begin
          ram_1_105 <= _GEN_11545;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_106 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_106 <= _GEN_1909;
        end else begin
          ram_1_106 <= _GEN_11546;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_107 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_107 <= _GEN_1910;
        end else begin
          ram_1_107 <= _GEN_11547;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_108 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_108 <= _GEN_1911;
        end else begin
          ram_1_108 <= _GEN_11548;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_109 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_109 <= _GEN_1912;
        end else begin
          ram_1_109 <= _GEN_11549;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_110 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_110 <= _GEN_1913;
        end else begin
          ram_1_110 <= _GEN_11550;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_111 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_111 <= _GEN_1914;
        end else begin
          ram_1_111 <= _GEN_11551;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_112 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_112 <= _GEN_1915;
        end else begin
          ram_1_112 <= _GEN_11552;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_113 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_113 <= _GEN_1916;
        end else begin
          ram_1_113 <= _GEN_11553;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_114 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_114 <= _GEN_1917;
        end else begin
          ram_1_114 <= _GEN_11554;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_115 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_115 <= _GEN_1918;
        end else begin
          ram_1_115 <= _GEN_11555;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_116 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_116 <= _GEN_1919;
        end else begin
          ram_1_116 <= _GEN_11556;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_117 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_117 <= _GEN_1920;
        end else begin
          ram_1_117 <= _GEN_11557;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_118 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_118 <= _GEN_1921;
        end else begin
          ram_1_118 <= _GEN_11558;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_119 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_119 <= _GEN_1922;
        end else begin
          ram_1_119 <= _GEN_11559;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_120 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_120 <= _GEN_1923;
        end else begin
          ram_1_120 <= _GEN_11560;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_121 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_121 <= _GEN_1924;
        end else begin
          ram_1_121 <= _GEN_11561;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_122 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_122 <= _GEN_1925;
        end else begin
          ram_1_122 <= _GEN_11562;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_123 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_123 <= _GEN_1926;
        end else begin
          ram_1_123 <= _GEN_11563;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_124 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_124 <= _GEN_1927;
        end else begin
          ram_1_124 <= _GEN_11564;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_125 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_125 <= _GEN_1928;
        end else begin
          ram_1_125 <= _GEN_11565;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_126 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_126 <= _GEN_1929;
        end else begin
          ram_1_126 <= _GEN_11566;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_127 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          ram_1_127 <= _GEN_1930;
        end else begin
          ram_1_127 <= _GEN_11567;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_0 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_0 <= _GEN_11183;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_1 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_1 <= _GEN_11184;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_2 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_2 <= _GEN_11185;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_3 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_3 <= _GEN_11186;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_4 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_4 <= _GEN_11187;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_5 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_5 <= _GEN_11188;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_6 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_6 <= _GEN_11189;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_7 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_7 <= _GEN_11190;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_8 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_8 <= _GEN_11191;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_9 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_9 <= _GEN_11192;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_10 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_10 <= _GEN_11193;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_11 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_11 <= _GEN_11194;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_12 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_12 <= _GEN_11195;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_13 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_13 <= _GEN_11196;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_14 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_14 <= _GEN_11197;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_15 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_15 <= _GEN_11198;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_16 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_16 <= _GEN_11199;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_17 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_17 <= _GEN_11200;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_18 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_18 <= _GEN_11201;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_19 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_19 <= _GEN_11202;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_20 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_20 <= _GEN_11203;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_21 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_21 <= _GEN_11204;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_22 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_22 <= _GEN_11205;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_23 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_23 <= _GEN_11206;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_24 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_24 <= _GEN_11207;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_25 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_25 <= _GEN_11208;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_26 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_26 <= _GEN_11209;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_27 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_27 <= _GEN_11210;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_28 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_28 <= _GEN_11211;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_29 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_29 <= _GEN_11212;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_30 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_30 <= _GEN_11213;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_31 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_31 <= _GEN_11214;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_32 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_32 <= _GEN_11215;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_33 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_33 <= _GEN_11216;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_34 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_34 <= _GEN_11217;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_35 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_35 <= _GEN_11218;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_36 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_36 <= _GEN_11219;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_37 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_37 <= _GEN_11220;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_38 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_38 <= _GEN_11221;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_39 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_39 <= _GEN_11222;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_40 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_40 <= _GEN_11223;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_41 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_41 <= _GEN_11224;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_42 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_42 <= _GEN_11225;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_43 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_43 <= _GEN_11226;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_44 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_44 <= _GEN_11227;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_45 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_45 <= _GEN_11228;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_46 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_46 <= _GEN_11229;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_47 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_47 <= _GEN_11230;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_48 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_48 <= _GEN_11231;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_49 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_49 <= _GEN_11232;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_50 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_50 <= _GEN_11233;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_51 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_51 <= _GEN_11234;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_52 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_52 <= _GEN_11235;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_53 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_53 <= _GEN_11236;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_54 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_54 <= _GEN_11237;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_55 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_55 <= _GEN_11238;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_56 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_56 <= _GEN_11239;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_57 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_57 <= _GEN_11240;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_58 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_58 <= _GEN_11241;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_59 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_59 <= _GEN_11242;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_60 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_60 <= _GEN_11243;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_61 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_61 <= _GEN_11244;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_62 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_62 <= _GEN_11245;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_63 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_63 <= _GEN_11246;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_64 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_64 <= _GEN_11247;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_65 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_65 <= _GEN_11248;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_66 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_66 <= _GEN_11249;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_67 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_67 <= _GEN_11250;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_68 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_68 <= _GEN_11251;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_69 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_69 <= _GEN_11252;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_70 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_70 <= _GEN_11253;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_71 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_71 <= _GEN_11254;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_72 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_72 <= _GEN_11255;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_73 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_73 <= _GEN_11256;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_74 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_74 <= _GEN_11257;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_75 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_75 <= _GEN_11258;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_76 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_76 <= _GEN_11259;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_77 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_77 <= _GEN_11260;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_78 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_78 <= _GEN_11261;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_79 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_79 <= _GEN_11262;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_80 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_80 <= _GEN_11263;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_81 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_81 <= _GEN_11264;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_82 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_82 <= _GEN_11265;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_83 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_83 <= _GEN_11266;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_84 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_84 <= _GEN_11267;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_85 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_85 <= _GEN_11268;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_86 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_86 <= _GEN_11269;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_87 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_87 <= _GEN_11270;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_88 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_88 <= _GEN_11271;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_89 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_89 <= _GEN_11272;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_90 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_90 <= _GEN_11273;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_91 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_91 <= _GEN_11274;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_92 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_92 <= _GEN_11275;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_93 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_93 <= _GEN_11276;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_94 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_94 <= _GEN_11277;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_95 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_95 <= _GEN_11278;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_96 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_96 <= _GEN_11279;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_97 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_97 <= _GEN_11280;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_98 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_98 <= _GEN_11281;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_99 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_99 <= _GEN_11282;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_100 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_100 <= _GEN_11283;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_101 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_101 <= _GEN_11284;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_102 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_102 <= _GEN_11285;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_103 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_103 <= _GEN_11286;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_104 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_104 <= _GEN_11287;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_105 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_105 <= _GEN_11288;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_106 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_106 <= _GEN_11289;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_107 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_107 <= _GEN_11290;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_108 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_108 <= _GEN_11291;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_109 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_109 <= _GEN_11292;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_110 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_110 <= _GEN_11293;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_111 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_111 <= _GEN_11294;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_112 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_112 <= _GEN_11295;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_113 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_113 <= _GEN_11296;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_114 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_114 <= _GEN_11297;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_115 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_115 <= _GEN_11298;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_116 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_116 <= _GEN_11299;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_117 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_117 <= _GEN_11300;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_118 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_118 <= _GEN_11301;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_119 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_119 <= _GEN_11302;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_120 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_120 <= _GEN_11303;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_121 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_121 <= _GEN_11304;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_122 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_122 <= _GEN_11305;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_123 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_123 <= _GEN_11306;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_124 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_124 <= _GEN_11307;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_125 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_125 <= _GEN_11308;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_126 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_126 <= _GEN_11309;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_127 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_0_127 <= _GEN_11310;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_0 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_0 <= _GEN_11568;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_1 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_1 <= _GEN_11569;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_2 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_2 <= _GEN_11570;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_3 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_3 <= _GEN_11571;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_4 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_4 <= _GEN_11572;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_5 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_5 <= _GEN_11573;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_6 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_6 <= _GEN_11574;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_7 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_7 <= _GEN_11575;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_8 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_8 <= _GEN_11576;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_9 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_9 <= _GEN_11577;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_10 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_10 <= _GEN_11578;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_11 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_11 <= _GEN_11579;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_12 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_12 <= _GEN_11580;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_13 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_13 <= _GEN_11581;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_14 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_14 <= _GEN_11582;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_15 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_15 <= _GEN_11583;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_16 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_16 <= _GEN_11584;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_17 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_17 <= _GEN_11585;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_18 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_18 <= _GEN_11586;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_19 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_19 <= _GEN_11587;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_20 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_20 <= _GEN_11588;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_21 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_21 <= _GEN_11589;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_22 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_22 <= _GEN_11590;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_23 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_23 <= _GEN_11591;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_24 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_24 <= _GEN_11592;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_25 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_25 <= _GEN_11593;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_26 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_26 <= _GEN_11594;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_27 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_27 <= _GEN_11595;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_28 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_28 <= _GEN_11596;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_29 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_29 <= _GEN_11597;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_30 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_30 <= _GEN_11598;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_31 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_31 <= _GEN_11599;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_32 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_32 <= _GEN_11600;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_33 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_33 <= _GEN_11601;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_34 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_34 <= _GEN_11602;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_35 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_35 <= _GEN_11603;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_36 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_36 <= _GEN_11604;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_37 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_37 <= _GEN_11605;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_38 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_38 <= _GEN_11606;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_39 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_39 <= _GEN_11607;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_40 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_40 <= _GEN_11608;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_41 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_41 <= _GEN_11609;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_42 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_42 <= _GEN_11610;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_43 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_43 <= _GEN_11611;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_44 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_44 <= _GEN_11612;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_45 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_45 <= _GEN_11613;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_46 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_46 <= _GEN_11614;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_47 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_47 <= _GEN_11615;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_48 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_48 <= _GEN_11616;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_49 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_49 <= _GEN_11617;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_50 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_50 <= _GEN_11618;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_51 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_51 <= _GEN_11619;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_52 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_52 <= _GEN_11620;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_53 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_53 <= _GEN_11621;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_54 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_54 <= _GEN_11622;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_55 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_55 <= _GEN_11623;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_56 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_56 <= _GEN_11624;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_57 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_57 <= _GEN_11625;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_58 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_58 <= _GEN_11626;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_59 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_59 <= _GEN_11627;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_60 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_60 <= _GEN_11628;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_61 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_61 <= _GEN_11629;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_62 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_62 <= _GEN_11630;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_63 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_63 <= _GEN_11631;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_64 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_64 <= _GEN_11632;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_65 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_65 <= _GEN_11633;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_66 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_66 <= _GEN_11634;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_67 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_67 <= _GEN_11635;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_68 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_68 <= _GEN_11636;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_69 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_69 <= _GEN_11637;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_70 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_70 <= _GEN_11638;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_71 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_71 <= _GEN_11639;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_72 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_72 <= _GEN_11640;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_73 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_73 <= _GEN_11641;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_74 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_74 <= _GEN_11642;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_75 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_75 <= _GEN_11643;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_76 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_76 <= _GEN_11644;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_77 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_77 <= _GEN_11645;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_78 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_78 <= _GEN_11646;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_79 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_79 <= _GEN_11647;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_80 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_80 <= _GEN_11648;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_81 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_81 <= _GEN_11649;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_82 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_82 <= _GEN_11650;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_83 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_83 <= _GEN_11651;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_84 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_84 <= _GEN_11652;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_85 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_85 <= _GEN_11653;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_86 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_86 <= _GEN_11654;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_87 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_87 <= _GEN_11655;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_88 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_88 <= _GEN_11656;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_89 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_89 <= _GEN_11657;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_90 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_90 <= _GEN_11658;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_91 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_91 <= _GEN_11659;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_92 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_92 <= _GEN_11660;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_93 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_93 <= _GEN_11661;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_94 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_94 <= _GEN_11662;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_95 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_95 <= _GEN_11663;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_96 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_96 <= _GEN_11664;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_97 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_97 <= _GEN_11665;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_98 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_98 <= _GEN_11666;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_99 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_99 <= _GEN_11667;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_100 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_100 <= _GEN_11668;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_101 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_101 <= _GEN_11669;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_102 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_102 <= _GEN_11670;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_103 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_103 <= _GEN_11671;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_104 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_104 <= _GEN_11672;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_105 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_105 <= _GEN_11673;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_106 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_106 <= _GEN_11674;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_107 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_107 <= _GEN_11675;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_108 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_108 <= _GEN_11676;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_109 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_109 <= _GEN_11677;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_110 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_110 <= _GEN_11678;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_111 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_111 <= _GEN_11679;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_112 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_112 <= _GEN_11680;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_113 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_113 <= _GEN_11681;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_114 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_114 <= _GEN_11682;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_115 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_115 <= _GEN_11683;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_116 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_116 <= _GEN_11684;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_117 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_117 <= _GEN_11685;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_118 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_118 <= _GEN_11686;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_119 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_119 <= _GEN_11687;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_120 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_120 <= _GEN_11688;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_121 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_121 <= _GEN_11689;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_122 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_122 <= _GEN_11690;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_123 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_123 <= _GEN_11691;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_124 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_124 <= _GEN_11692;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_125 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_125 <= _GEN_11693;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_126 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_126 <= _GEN_11694;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_127 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          tag_1_127 <= _GEN_11695;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_0 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_0 <= _GEN_11311;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_1 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_1 <= _GEN_11312;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_2 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_2 <= _GEN_11313;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_3 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_3 <= _GEN_11314;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_4 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_4 <= _GEN_11315;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_5 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_5 <= _GEN_11316;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_6 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_6 <= _GEN_11317;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_7 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_7 <= _GEN_11318;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_8 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_8 <= _GEN_11319;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_9 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_9 <= _GEN_11320;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_10 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_10 <= _GEN_11321;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_11 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_11 <= _GEN_11322;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_12 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_12 <= _GEN_11323;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_13 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_13 <= _GEN_11324;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_14 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_14 <= _GEN_11325;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_15 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_15 <= _GEN_11326;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_16 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_16 <= _GEN_11327;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_17 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_17 <= _GEN_11328;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_18 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_18 <= _GEN_11329;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_19 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_19 <= _GEN_11330;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_20 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_20 <= _GEN_11331;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_21 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_21 <= _GEN_11332;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_22 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_22 <= _GEN_11333;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_23 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_23 <= _GEN_11334;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_24 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_24 <= _GEN_11335;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_25 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_25 <= _GEN_11336;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_26 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_26 <= _GEN_11337;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_27 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_27 <= _GEN_11338;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_28 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_28 <= _GEN_11339;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_29 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_29 <= _GEN_11340;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_30 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_30 <= _GEN_11341;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_31 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_31 <= _GEN_11342;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_32 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_32 <= _GEN_11343;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_33 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_33 <= _GEN_11344;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_34 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_34 <= _GEN_11345;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_35 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_35 <= _GEN_11346;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_36 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_36 <= _GEN_11347;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_37 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_37 <= _GEN_11348;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_38 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_38 <= _GEN_11349;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_39 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_39 <= _GEN_11350;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_40 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_40 <= _GEN_11351;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_41 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_41 <= _GEN_11352;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_42 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_42 <= _GEN_11353;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_43 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_43 <= _GEN_11354;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_44 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_44 <= _GEN_11355;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_45 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_45 <= _GEN_11356;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_46 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_46 <= _GEN_11357;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_47 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_47 <= _GEN_11358;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_48 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_48 <= _GEN_11359;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_49 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_49 <= _GEN_11360;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_50 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_50 <= _GEN_11361;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_51 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_51 <= _GEN_11362;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_52 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_52 <= _GEN_11363;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_53 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_53 <= _GEN_11364;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_54 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_54 <= _GEN_11365;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_55 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_55 <= _GEN_11366;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_56 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_56 <= _GEN_11367;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_57 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_57 <= _GEN_11368;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_58 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_58 <= _GEN_11369;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_59 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_59 <= _GEN_11370;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_60 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_60 <= _GEN_11371;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_61 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_61 <= _GEN_11372;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_62 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_62 <= _GEN_11373;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_63 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_63 <= _GEN_11374;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_64 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_64 <= _GEN_11375;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_65 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_65 <= _GEN_11376;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_66 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_66 <= _GEN_11377;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_67 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_67 <= _GEN_11378;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_68 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_68 <= _GEN_11379;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_69 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_69 <= _GEN_11380;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_70 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_70 <= _GEN_11381;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_71 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_71 <= _GEN_11382;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_72 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_72 <= _GEN_11383;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_73 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_73 <= _GEN_11384;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_74 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_74 <= _GEN_11385;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_75 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_75 <= _GEN_11386;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_76 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_76 <= _GEN_11387;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_77 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_77 <= _GEN_11388;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_78 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_78 <= _GEN_11389;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_79 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_79 <= _GEN_11390;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_80 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_80 <= _GEN_11391;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_81 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_81 <= _GEN_11392;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_82 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_82 <= _GEN_11393;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_83 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_83 <= _GEN_11394;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_84 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_84 <= _GEN_11395;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_85 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_85 <= _GEN_11396;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_86 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_86 <= _GEN_11397;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_87 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_87 <= _GEN_11398;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_88 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_88 <= _GEN_11399;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_89 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_89 <= _GEN_11400;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_90 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_90 <= _GEN_11401;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_91 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_91 <= _GEN_11402;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_92 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_92 <= _GEN_11403;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_93 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_93 <= _GEN_11404;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_94 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_94 <= _GEN_11405;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_95 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_95 <= _GEN_11406;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_96 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_96 <= _GEN_11407;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_97 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_97 <= _GEN_11408;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_98 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_98 <= _GEN_11409;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_99 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_99 <= _GEN_11410;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_100 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_100 <= _GEN_11411;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_101 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_101 <= _GEN_11412;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_102 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_102 <= _GEN_11413;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_103 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_103 <= _GEN_11414;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_104 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_104 <= _GEN_11415;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_105 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_105 <= _GEN_11416;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_106 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_106 <= _GEN_11417;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_107 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_107 <= _GEN_11418;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_108 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_108 <= _GEN_11419;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_109 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_109 <= _GEN_11420;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_110 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_110 <= _GEN_11421;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_111 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_111 <= _GEN_11422;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_112 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_112 <= _GEN_11423;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_113 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_113 <= _GEN_11424;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_114 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_114 <= _GEN_11425;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_115 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_115 <= _GEN_11426;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_116 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_116 <= _GEN_11427;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_117 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_117 <= _GEN_11428;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_118 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_118 <= _GEN_11429;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_119 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_119 <= _GEN_11430;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_120 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_120 <= _GEN_11431;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_121 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_121 <= _GEN_11432;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_122 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_122 <= _GEN_11433;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_123 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_123 <= _GEN_11434;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_124 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_124 <= _GEN_11435;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_125 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_125 <= _GEN_11436;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_126 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_126 <= _GEN_11437;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_127 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_0_127 <= _GEN_11438;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_0 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_0 <= _GEN_11696;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_1 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_1 <= _GEN_11697;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_2 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_2 <= _GEN_11698;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_3 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_3 <= _GEN_11699;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_4 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_4 <= _GEN_11700;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_5 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_5 <= _GEN_11701;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_6 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_6 <= _GEN_11702;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_7 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_7 <= _GEN_11703;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_8 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_8 <= _GEN_11704;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_9 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_9 <= _GEN_11705;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_10 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_10 <= _GEN_11706;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_11 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_11 <= _GEN_11707;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_12 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_12 <= _GEN_11708;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_13 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_13 <= _GEN_11709;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_14 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_14 <= _GEN_11710;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_15 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_15 <= _GEN_11711;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_16 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_16 <= _GEN_11712;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_17 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_17 <= _GEN_11713;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_18 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_18 <= _GEN_11714;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_19 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_19 <= _GEN_11715;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_20 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_20 <= _GEN_11716;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_21 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_21 <= _GEN_11717;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_22 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_22 <= _GEN_11718;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_23 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_23 <= _GEN_11719;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_24 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_24 <= _GEN_11720;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_25 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_25 <= _GEN_11721;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_26 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_26 <= _GEN_11722;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_27 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_27 <= _GEN_11723;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_28 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_28 <= _GEN_11724;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_29 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_29 <= _GEN_11725;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_30 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_30 <= _GEN_11726;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_31 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_31 <= _GEN_11727;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_32 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_32 <= _GEN_11728;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_33 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_33 <= _GEN_11729;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_34 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_34 <= _GEN_11730;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_35 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_35 <= _GEN_11731;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_36 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_36 <= _GEN_11732;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_37 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_37 <= _GEN_11733;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_38 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_38 <= _GEN_11734;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_39 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_39 <= _GEN_11735;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_40 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_40 <= _GEN_11736;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_41 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_41 <= _GEN_11737;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_42 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_42 <= _GEN_11738;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_43 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_43 <= _GEN_11739;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_44 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_44 <= _GEN_11740;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_45 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_45 <= _GEN_11741;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_46 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_46 <= _GEN_11742;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_47 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_47 <= _GEN_11743;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_48 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_48 <= _GEN_11744;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_49 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_49 <= _GEN_11745;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_50 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_50 <= _GEN_11746;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_51 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_51 <= _GEN_11747;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_52 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_52 <= _GEN_11748;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_53 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_53 <= _GEN_11749;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_54 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_54 <= _GEN_11750;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_55 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_55 <= _GEN_11751;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_56 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_56 <= _GEN_11752;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_57 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_57 <= _GEN_11753;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_58 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_58 <= _GEN_11754;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_59 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_59 <= _GEN_11755;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_60 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_60 <= _GEN_11756;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_61 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_61 <= _GEN_11757;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_62 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_62 <= _GEN_11758;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_63 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_63 <= _GEN_11759;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_64 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_64 <= _GEN_11760;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_65 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_65 <= _GEN_11761;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_66 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_66 <= _GEN_11762;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_67 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_67 <= _GEN_11763;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_68 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_68 <= _GEN_11764;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_69 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_69 <= _GEN_11765;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_70 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_70 <= _GEN_11766;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_71 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_71 <= _GEN_11767;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_72 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_72 <= _GEN_11768;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_73 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_73 <= _GEN_11769;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_74 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_74 <= _GEN_11770;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_75 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_75 <= _GEN_11771;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_76 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_76 <= _GEN_11772;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_77 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_77 <= _GEN_11773;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_78 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_78 <= _GEN_11774;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_79 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_79 <= _GEN_11775;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_80 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_80 <= _GEN_11776;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_81 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_81 <= _GEN_11777;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_82 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_82 <= _GEN_11778;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_83 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_83 <= _GEN_11779;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_84 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_84 <= _GEN_11780;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_85 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_85 <= _GEN_11781;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_86 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_86 <= _GEN_11782;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_87 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_87 <= _GEN_11783;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_88 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_88 <= _GEN_11784;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_89 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_89 <= _GEN_11785;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_90 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_90 <= _GEN_11786;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_91 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_91 <= _GEN_11787;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_92 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_92 <= _GEN_11788;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_93 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_93 <= _GEN_11789;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_94 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_94 <= _GEN_11790;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_95 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_95 <= _GEN_11791;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_96 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_96 <= _GEN_11792;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_97 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_97 <= _GEN_11793;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_98 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_98 <= _GEN_11794;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_99 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_99 <= _GEN_11795;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_100 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_100 <= _GEN_11796;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_101 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_101 <= _GEN_11797;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_102 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_102 <= _GEN_11798;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_103 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_103 <= _GEN_11799;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_104 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_104 <= _GEN_11800;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_105 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_105 <= _GEN_11801;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_106 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_106 <= _GEN_11802;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_107 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_107 <= _GEN_11803;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_108 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_108 <= _GEN_11804;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_109 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_109 <= _GEN_11805;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_110 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_110 <= _GEN_11806;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_111 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_111 <= _GEN_11807;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_112 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_112 <= _GEN_11808;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_113 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_113 <= _GEN_11809;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_114 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_114 <= _GEN_11810;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_115 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_115 <= _GEN_11811;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_116 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_116 <= _GEN_11812;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_117 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_117 <= _GEN_11813;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_118 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_118 <= _GEN_11814;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_119 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_119 <= _GEN_11815;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_120 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_120 <= _GEN_11816;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_121 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_121 <= _GEN_11817;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_122 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_122 <= _GEN_11818;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_123 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_123 <= _GEN_11819;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_124 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_124 <= _GEN_11820;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_125 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_125 <= _GEN_11821;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_126 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_126 <= _GEN_11822;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_127 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          valid_1_127 <= _GEN_11823;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_0 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_0 <= _GEN_1675;
        end else begin
          dirty_0_0 <= _GEN_11826;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_1 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_1 <= _GEN_1676;
        end else begin
          dirty_0_1 <= _GEN_11827;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_2 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_2 <= _GEN_1677;
        end else begin
          dirty_0_2 <= _GEN_11828;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_3 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_3 <= _GEN_1678;
        end else begin
          dirty_0_3 <= _GEN_11829;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_4 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_4 <= _GEN_1679;
        end else begin
          dirty_0_4 <= _GEN_11830;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_5 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_5 <= _GEN_1680;
        end else begin
          dirty_0_5 <= _GEN_11831;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_6 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_6 <= _GEN_1681;
        end else begin
          dirty_0_6 <= _GEN_11832;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_7 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_7 <= _GEN_1682;
        end else begin
          dirty_0_7 <= _GEN_11833;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_8 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_8 <= _GEN_1683;
        end else begin
          dirty_0_8 <= _GEN_11834;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_9 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_9 <= _GEN_1684;
        end else begin
          dirty_0_9 <= _GEN_11835;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_10 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_10 <= _GEN_1685;
        end else begin
          dirty_0_10 <= _GEN_11836;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_11 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_11 <= _GEN_1686;
        end else begin
          dirty_0_11 <= _GEN_11837;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_12 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_12 <= _GEN_1687;
        end else begin
          dirty_0_12 <= _GEN_11838;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_13 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_13 <= _GEN_1688;
        end else begin
          dirty_0_13 <= _GEN_11839;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_14 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_14 <= _GEN_1689;
        end else begin
          dirty_0_14 <= _GEN_11840;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_15 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_15 <= _GEN_1690;
        end else begin
          dirty_0_15 <= _GEN_11841;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_16 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_16 <= _GEN_1691;
        end else begin
          dirty_0_16 <= _GEN_11842;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_17 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_17 <= _GEN_1692;
        end else begin
          dirty_0_17 <= _GEN_11843;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_18 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_18 <= _GEN_1693;
        end else begin
          dirty_0_18 <= _GEN_11844;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_19 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_19 <= _GEN_1694;
        end else begin
          dirty_0_19 <= _GEN_11845;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_20 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_20 <= _GEN_1695;
        end else begin
          dirty_0_20 <= _GEN_11846;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_21 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_21 <= _GEN_1696;
        end else begin
          dirty_0_21 <= _GEN_11847;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_22 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_22 <= _GEN_1697;
        end else begin
          dirty_0_22 <= _GEN_11848;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_23 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_23 <= _GEN_1698;
        end else begin
          dirty_0_23 <= _GEN_11849;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_24 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_24 <= _GEN_1699;
        end else begin
          dirty_0_24 <= _GEN_11850;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_25 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_25 <= _GEN_1700;
        end else begin
          dirty_0_25 <= _GEN_11851;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_26 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_26 <= _GEN_1701;
        end else begin
          dirty_0_26 <= _GEN_11852;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_27 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_27 <= _GEN_1702;
        end else begin
          dirty_0_27 <= _GEN_11853;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_28 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_28 <= _GEN_1703;
        end else begin
          dirty_0_28 <= _GEN_11854;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_29 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_29 <= _GEN_1704;
        end else begin
          dirty_0_29 <= _GEN_11855;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_30 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_30 <= _GEN_1705;
        end else begin
          dirty_0_30 <= _GEN_11856;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_31 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_31 <= _GEN_1706;
        end else begin
          dirty_0_31 <= _GEN_11857;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_32 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_32 <= _GEN_1707;
        end else begin
          dirty_0_32 <= _GEN_11858;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_33 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_33 <= _GEN_1708;
        end else begin
          dirty_0_33 <= _GEN_11859;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_34 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_34 <= _GEN_1709;
        end else begin
          dirty_0_34 <= _GEN_11860;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_35 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_35 <= _GEN_1710;
        end else begin
          dirty_0_35 <= _GEN_11861;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_36 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_36 <= _GEN_1711;
        end else begin
          dirty_0_36 <= _GEN_11862;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_37 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_37 <= _GEN_1712;
        end else begin
          dirty_0_37 <= _GEN_11863;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_38 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_38 <= _GEN_1713;
        end else begin
          dirty_0_38 <= _GEN_11864;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_39 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_39 <= _GEN_1714;
        end else begin
          dirty_0_39 <= _GEN_11865;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_40 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_40 <= _GEN_1715;
        end else begin
          dirty_0_40 <= _GEN_11866;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_41 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_41 <= _GEN_1716;
        end else begin
          dirty_0_41 <= _GEN_11867;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_42 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_42 <= _GEN_1717;
        end else begin
          dirty_0_42 <= _GEN_11868;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_43 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_43 <= _GEN_1718;
        end else begin
          dirty_0_43 <= _GEN_11869;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_44 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_44 <= _GEN_1719;
        end else begin
          dirty_0_44 <= _GEN_11870;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_45 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_45 <= _GEN_1720;
        end else begin
          dirty_0_45 <= _GEN_11871;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_46 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_46 <= _GEN_1721;
        end else begin
          dirty_0_46 <= _GEN_11872;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_47 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_47 <= _GEN_1722;
        end else begin
          dirty_0_47 <= _GEN_11873;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_48 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_48 <= _GEN_1723;
        end else begin
          dirty_0_48 <= _GEN_11874;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_49 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_49 <= _GEN_1724;
        end else begin
          dirty_0_49 <= _GEN_11875;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_50 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_50 <= _GEN_1725;
        end else begin
          dirty_0_50 <= _GEN_11876;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_51 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_51 <= _GEN_1726;
        end else begin
          dirty_0_51 <= _GEN_11877;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_52 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_52 <= _GEN_1727;
        end else begin
          dirty_0_52 <= _GEN_11878;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_53 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_53 <= _GEN_1728;
        end else begin
          dirty_0_53 <= _GEN_11879;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_54 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_54 <= _GEN_1729;
        end else begin
          dirty_0_54 <= _GEN_11880;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_55 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_55 <= _GEN_1730;
        end else begin
          dirty_0_55 <= _GEN_11881;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_56 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_56 <= _GEN_1731;
        end else begin
          dirty_0_56 <= _GEN_11882;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_57 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_57 <= _GEN_1732;
        end else begin
          dirty_0_57 <= _GEN_11883;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_58 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_58 <= _GEN_1733;
        end else begin
          dirty_0_58 <= _GEN_11884;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_59 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_59 <= _GEN_1734;
        end else begin
          dirty_0_59 <= _GEN_11885;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_60 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_60 <= _GEN_1735;
        end else begin
          dirty_0_60 <= _GEN_11886;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_61 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_61 <= _GEN_1736;
        end else begin
          dirty_0_61 <= _GEN_11887;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_62 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_62 <= _GEN_1737;
        end else begin
          dirty_0_62 <= _GEN_11888;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_63 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_63 <= _GEN_1738;
        end else begin
          dirty_0_63 <= _GEN_11889;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_64 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_64 <= _GEN_1739;
        end else begin
          dirty_0_64 <= _GEN_11890;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_65 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_65 <= _GEN_1740;
        end else begin
          dirty_0_65 <= _GEN_11891;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_66 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_66 <= _GEN_1741;
        end else begin
          dirty_0_66 <= _GEN_11892;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_67 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_67 <= _GEN_1742;
        end else begin
          dirty_0_67 <= _GEN_11893;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_68 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_68 <= _GEN_1743;
        end else begin
          dirty_0_68 <= _GEN_11894;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_69 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_69 <= _GEN_1744;
        end else begin
          dirty_0_69 <= _GEN_11895;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_70 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_70 <= _GEN_1745;
        end else begin
          dirty_0_70 <= _GEN_11896;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_71 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_71 <= _GEN_1746;
        end else begin
          dirty_0_71 <= _GEN_11897;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_72 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_72 <= _GEN_1747;
        end else begin
          dirty_0_72 <= _GEN_11898;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_73 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_73 <= _GEN_1748;
        end else begin
          dirty_0_73 <= _GEN_11899;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_74 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_74 <= _GEN_1749;
        end else begin
          dirty_0_74 <= _GEN_11900;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_75 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_75 <= _GEN_1750;
        end else begin
          dirty_0_75 <= _GEN_11901;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_76 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_76 <= _GEN_1751;
        end else begin
          dirty_0_76 <= _GEN_11902;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_77 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_77 <= _GEN_1752;
        end else begin
          dirty_0_77 <= _GEN_11903;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_78 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_78 <= _GEN_1753;
        end else begin
          dirty_0_78 <= _GEN_11904;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_79 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_79 <= _GEN_1754;
        end else begin
          dirty_0_79 <= _GEN_11905;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_80 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_80 <= _GEN_1755;
        end else begin
          dirty_0_80 <= _GEN_11906;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_81 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_81 <= _GEN_1756;
        end else begin
          dirty_0_81 <= _GEN_11907;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_82 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_82 <= _GEN_1757;
        end else begin
          dirty_0_82 <= _GEN_11908;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_83 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_83 <= _GEN_1758;
        end else begin
          dirty_0_83 <= _GEN_11909;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_84 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_84 <= _GEN_1759;
        end else begin
          dirty_0_84 <= _GEN_11910;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_85 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_85 <= _GEN_1760;
        end else begin
          dirty_0_85 <= _GEN_11911;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_86 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_86 <= _GEN_1761;
        end else begin
          dirty_0_86 <= _GEN_11912;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_87 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_87 <= _GEN_1762;
        end else begin
          dirty_0_87 <= _GEN_11913;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_88 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_88 <= _GEN_1763;
        end else begin
          dirty_0_88 <= _GEN_11914;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_89 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_89 <= _GEN_1764;
        end else begin
          dirty_0_89 <= _GEN_11915;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_90 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_90 <= _GEN_1765;
        end else begin
          dirty_0_90 <= _GEN_11916;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_91 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_91 <= _GEN_1766;
        end else begin
          dirty_0_91 <= _GEN_11917;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_92 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_92 <= _GEN_1767;
        end else begin
          dirty_0_92 <= _GEN_11918;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_93 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_93 <= _GEN_1768;
        end else begin
          dirty_0_93 <= _GEN_11919;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_94 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_94 <= _GEN_1769;
        end else begin
          dirty_0_94 <= _GEN_11920;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_95 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_95 <= _GEN_1770;
        end else begin
          dirty_0_95 <= _GEN_11921;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_96 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_96 <= _GEN_1771;
        end else begin
          dirty_0_96 <= _GEN_11922;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_97 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_97 <= _GEN_1772;
        end else begin
          dirty_0_97 <= _GEN_11923;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_98 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_98 <= _GEN_1773;
        end else begin
          dirty_0_98 <= _GEN_11924;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_99 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_99 <= _GEN_1774;
        end else begin
          dirty_0_99 <= _GEN_11925;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_100 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_100 <= _GEN_1775;
        end else begin
          dirty_0_100 <= _GEN_11926;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_101 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_101 <= _GEN_1776;
        end else begin
          dirty_0_101 <= _GEN_11927;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_102 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_102 <= _GEN_1777;
        end else begin
          dirty_0_102 <= _GEN_11928;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_103 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_103 <= _GEN_1778;
        end else begin
          dirty_0_103 <= _GEN_11929;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_104 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_104 <= _GEN_1779;
        end else begin
          dirty_0_104 <= _GEN_11930;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_105 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_105 <= _GEN_1780;
        end else begin
          dirty_0_105 <= _GEN_11931;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_106 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_106 <= _GEN_1781;
        end else begin
          dirty_0_106 <= _GEN_11932;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_107 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_107 <= _GEN_1782;
        end else begin
          dirty_0_107 <= _GEN_11933;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_108 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_108 <= _GEN_1783;
        end else begin
          dirty_0_108 <= _GEN_11934;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_109 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_109 <= _GEN_1784;
        end else begin
          dirty_0_109 <= _GEN_11935;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_110 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_110 <= _GEN_1785;
        end else begin
          dirty_0_110 <= _GEN_11936;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_111 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_111 <= _GEN_1786;
        end else begin
          dirty_0_111 <= _GEN_11937;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_112 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_112 <= _GEN_1787;
        end else begin
          dirty_0_112 <= _GEN_11938;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_113 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_113 <= _GEN_1788;
        end else begin
          dirty_0_113 <= _GEN_11939;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_114 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_114 <= _GEN_1789;
        end else begin
          dirty_0_114 <= _GEN_11940;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_115 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_115 <= _GEN_1790;
        end else begin
          dirty_0_115 <= _GEN_11941;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_116 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_116 <= _GEN_1791;
        end else begin
          dirty_0_116 <= _GEN_11942;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_117 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_117 <= _GEN_1792;
        end else begin
          dirty_0_117 <= _GEN_11943;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_118 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_118 <= _GEN_1793;
        end else begin
          dirty_0_118 <= _GEN_11944;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_119 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_119 <= _GEN_1794;
        end else begin
          dirty_0_119 <= _GEN_11945;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_120 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_120 <= _GEN_1795;
        end else begin
          dirty_0_120 <= _GEN_11946;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_121 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_121 <= _GEN_1796;
        end else begin
          dirty_0_121 <= _GEN_11947;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_122 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_122 <= _GEN_1797;
        end else begin
          dirty_0_122 <= _GEN_11948;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_123 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_123 <= _GEN_1798;
        end else begin
          dirty_0_123 <= _GEN_11949;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_124 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_124 <= _GEN_1799;
        end else begin
          dirty_0_124 <= _GEN_11950;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_125 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_125 <= _GEN_1800;
        end else begin
          dirty_0_125 <= _GEN_11951;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_126 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_126 <= _GEN_1801;
        end else begin
          dirty_0_126 <= _GEN_11952;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_127 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_0_127 <= _GEN_1802;
        end else begin
          dirty_0_127 <= _GEN_11953;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_0 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_0 <= _GEN_1931;
        end else begin
          dirty_1_0 <= _GEN_11954;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_1 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_1 <= _GEN_1932;
        end else begin
          dirty_1_1 <= _GEN_11955;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_2 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_2 <= _GEN_1933;
        end else begin
          dirty_1_2 <= _GEN_11956;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_3 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_3 <= _GEN_1934;
        end else begin
          dirty_1_3 <= _GEN_11957;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_4 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_4 <= _GEN_1935;
        end else begin
          dirty_1_4 <= _GEN_11958;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_5 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_5 <= _GEN_1936;
        end else begin
          dirty_1_5 <= _GEN_11959;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_6 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_6 <= _GEN_1937;
        end else begin
          dirty_1_6 <= _GEN_11960;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_7 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_7 <= _GEN_1938;
        end else begin
          dirty_1_7 <= _GEN_11961;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_8 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_8 <= _GEN_1939;
        end else begin
          dirty_1_8 <= _GEN_11962;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_9 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_9 <= _GEN_1940;
        end else begin
          dirty_1_9 <= _GEN_11963;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_10 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_10 <= _GEN_1941;
        end else begin
          dirty_1_10 <= _GEN_11964;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_11 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_11 <= _GEN_1942;
        end else begin
          dirty_1_11 <= _GEN_11965;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_12 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_12 <= _GEN_1943;
        end else begin
          dirty_1_12 <= _GEN_11966;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_13 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_13 <= _GEN_1944;
        end else begin
          dirty_1_13 <= _GEN_11967;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_14 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_14 <= _GEN_1945;
        end else begin
          dirty_1_14 <= _GEN_11968;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_15 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_15 <= _GEN_1946;
        end else begin
          dirty_1_15 <= _GEN_11969;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_16 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_16 <= _GEN_1947;
        end else begin
          dirty_1_16 <= _GEN_11970;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_17 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_17 <= _GEN_1948;
        end else begin
          dirty_1_17 <= _GEN_11971;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_18 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_18 <= _GEN_1949;
        end else begin
          dirty_1_18 <= _GEN_11972;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_19 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_19 <= _GEN_1950;
        end else begin
          dirty_1_19 <= _GEN_11973;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_20 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_20 <= _GEN_1951;
        end else begin
          dirty_1_20 <= _GEN_11974;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_21 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_21 <= _GEN_1952;
        end else begin
          dirty_1_21 <= _GEN_11975;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_22 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_22 <= _GEN_1953;
        end else begin
          dirty_1_22 <= _GEN_11976;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_23 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_23 <= _GEN_1954;
        end else begin
          dirty_1_23 <= _GEN_11977;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_24 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_24 <= _GEN_1955;
        end else begin
          dirty_1_24 <= _GEN_11978;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_25 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_25 <= _GEN_1956;
        end else begin
          dirty_1_25 <= _GEN_11979;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_26 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_26 <= _GEN_1957;
        end else begin
          dirty_1_26 <= _GEN_11980;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_27 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_27 <= _GEN_1958;
        end else begin
          dirty_1_27 <= _GEN_11981;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_28 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_28 <= _GEN_1959;
        end else begin
          dirty_1_28 <= _GEN_11982;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_29 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_29 <= _GEN_1960;
        end else begin
          dirty_1_29 <= _GEN_11983;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_30 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_30 <= _GEN_1961;
        end else begin
          dirty_1_30 <= _GEN_11984;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_31 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_31 <= _GEN_1962;
        end else begin
          dirty_1_31 <= _GEN_11985;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_32 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_32 <= _GEN_1963;
        end else begin
          dirty_1_32 <= _GEN_11986;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_33 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_33 <= _GEN_1964;
        end else begin
          dirty_1_33 <= _GEN_11987;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_34 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_34 <= _GEN_1965;
        end else begin
          dirty_1_34 <= _GEN_11988;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_35 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_35 <= _GEN_1966;
        end else begin
          dirty_1_35 <= _GEN_11989;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_36 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_36 <= _GEN_1967;
        end else begin
          dirty_1_36 <= _GEN_11990;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_37 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_37 <= _GEN_1968;
        end else begin
          dirty_1_37 <= _GEN_11991;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_38 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_38 <= _GEN_1969;
        end else begin
          dirty_1_38 <= _GEN_11992;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_39 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_39 <= _GEN_1970;
        end else begin
          dirty_1_39 <= _GEN_11993;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_40 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_40 <= _GEN_1971;
        end else begin
          dirty_1_40 <= _GEN_11994;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_41 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_41 <= _GEN_1972;
        end else begin
          dirty_1_41 <= _GEN_11995;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_42 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_42 <= _GEN_1973;
        end else begin
          dirty_1_42 <= _GEN_11996;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_43 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_43 <= _GEN_1974;
        end else begin
          dirty_1_43 <= _GEN_11997;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_44 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_44 <= _GEN_1975;
        end else begin
          dirty_1_44 <= _GEN_11998;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_45 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_45 <= _GEN_1976;
        end else begin
          dirty_1_45 <= _GEN_11999;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_46 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_46 <= _GEN_1977;
        end else begin
          dirty_1_46 <= _GEN_12000;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_47 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_47 <= _GEN_1978;
        end else begin
          dirty_1_47 <= _GEN_12001;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_48 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_48 <= _GEN_1979;
        end else begin
          dirty_1_48 <= _GEN_12002;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_49 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_49 <= _GEN_1980;
        end else begin
          dirty_1_49 <= _GEN_12003;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_50 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_50 <= _GEN_1981;
        end else begin
          dirty_1_50 <= _GEN_12004;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_51 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_51 <= _GEN_1982;
        end else begin
          dirty_1_51 <= _GEN_12005;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_52 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_52 <= _GEN_1983;
        end else begin
          dirty_1_52 <= _GEN_12006;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_53 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_53 <= _GEN_1984;
        end else begin
          dirty_1_53 <= _GEN_12007;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_54 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_54 <= _GEN_1985;
        end else begin
          dirty_1_54 <= _GEN_12008;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_55 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_55 <= _GEN_1986;
        end else begin
          dirty_1_55 <= _GEN_12009;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_56 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_56 <= _GEN_1987;
        end else begin
          dirty_1_56 <= _GEN_12010;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_57 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_57 <= _GEN_1988;
        end else begin
          dirty_1_57 <= _GEN_12011;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_58 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_58 <= _GEN_1989;
        end else begin
          dirty_1_58 <= _GEN_12012;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_59 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_59 <= _GEN_1990;
        end else begin
          dirty_1_59 <= _GEN_12013;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_60 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_60 <= _GEN_1991;
        end else begin
          dirty_1_60 <= _GEN_12014;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_61 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_61 <= _GEN_1992;
        end else begin
          dirty_1_61 <= _GEN_12015;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_62 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_62 <= _GEN_1993;
        end else begin
          dirty_1_62 <= _GEN_12016;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_63 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_63 <= _GEN_1994;
        end else begin
          dirty_1_63 <= _GEN_12017;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_64 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_64 <= _GEN_1995;
        end else begin
          dirty_1_64 <= _GEN_12018;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_65 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_65 <= _GEN_1996;
        end else begin
          dirty_1_65 <= _GEN_12019;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_66 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_66 <= _GEN_1997;
        end else begin
          dirty_1_66 <= _GEN_12020;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_67 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_67 <= _GEN_1998;
        end else begin
          dirty_1_67 <= _GEN_12021;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_68 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_68 <= _GEN_1999;
        end else begin
          dirty_1_68 <= _GEN_12022;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_69 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_69 <= _GEN_2000;
        end else begin
          dirty_1_69 <= _GEN_12023;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_70 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_70 <= _GEN_2001;
        end else begin
          dirty_1_70 <= _GEN_12024;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_71 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_71 <= _GEN_2002;
        end else begin
          dirty_1_71 <= _GEN_12025;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_72 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_72 <= _GEN_2003;
        end else begin
          dirty_1_72 <= _GEN_12026;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_73 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_73 <= _GEN_2004;
        end else begin
          dirty_1_73 <= _GEN_12027;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_74 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_74 <= _GEN_2005;
        end else begin
          dirty_1_74 <= _GEN_12028;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_75 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_75 <= _GEN_2006;
        end else begin
          dirty_1_75 <= _GEN_12029;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_76 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_76 <= _GEN_2007;
        end else begin
          dirty_1_76 <= _GEN_12030;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_77 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_77 <= _GEN_2008;
        end else begin
          dirty_1_77 <= _GEN_12031;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_78 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_78 <= _GEN_2009;
        end else begin
          dirty_1_78 <= _GEN_12032;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_79 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_79 <= _GEN_2010;
        end else begin
          dirty_1_79 <= _GEN_12033;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_80 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_80 <= _GEN_2011;
        end else begin
          dirty_1_80 <= _GEN_12034;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_81 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_81 <= _GEN_2012;
        end else begin
          dirty_1_81 <= _GEN_12035;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_82 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_82 <= _GEN_2013;
        end else begin
          dirty_1_82 <= _GEN_12036;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_83 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_83 <= _GEN_2014;
        end else begin
          dirty_1_83 <= _GEN_12037;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_84 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_84 <= _GEN_2015;
        end else begin
          dirty_1_84 <= _GEN_12038;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_85 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_85 <= _GEN_2016;
        end else begin
          dirty_1_85 <= _GEN_12039;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_86 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_86 <= _GEN_2017;
        end else begin
          dirty_1_86 <= _GEN_12040;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_87 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_87 <= _GEN_2018;
        end else begin
          dirty_1_87 <= _GEN_12041;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_88 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_88 <= _GEN_2019;
        end else begin
          dirty_1_88 <= _GEN_12042;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_89 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_89 <= _GEN_2020;
        end else begin
          dirty_1_89 <= _GEN_12043;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_90 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_90 <= _GEN_2021;
        end else begin
          dirty_1_90 <= _GEN_12044;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_91 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_91 <= _GEN_2022;
        end else begin
          dirty_1_91 <= _GEN_12045;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_92 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_92 <= _GEN_2023;
        end else begin
          dirty_1_92 <= _GEN_12046;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_93 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_93 <= _GEN_2024;
        end else begin
          dirty_1_93 <= _GEN_12047;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_94 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_94 <= _GEN_2025;
        end else begin
          dirty_1_94 <= _GEN_12048;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_95 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_95 <= _GEN_2026;
        end else begin
          dirty_1_95 <= _GEN_12049;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_96 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_96 <= _GEN_2027;
        end else begin
          dirty_1_96 <= _GEN_12050;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_97 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_97 <= _GEN_2028;
        end else begin
          dirty_1_97 <= _GEN_12051;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_98 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_98 <= _GEN_2029;
        end else begin
          dirty_1_98 <= _GEN_12052;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_99 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_99 <= _GEN_2030;
        end else begin
          dirty_1_99 <= _GEN_12053;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_100 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_100 <= _GEN_2031;
        end else begin
          dirty_1_100 <= _GEN_12054;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_101 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_101 <= _GEN_2032;
        end else begin
          dirty_1_101 <= _GEN_12055;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_102 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_102 <= _GEN_2033;
        end else begin
          dirty_1_102 <= _GEN_12056;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_103 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_103 <= _GEN_2034;
        end else begin
          dirty_1_103 <= _GEN_12057;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_104 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_104 <= _GEN_2035;
        end else begin
          dirty_1_104 <= _GEN_12058;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_105 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_105 <= _GEN_2036;
        end else begin
          dirty_1_105 <= _GEN_12059;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_106 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_106 <= _GEN_2037;
        end else begin
          dirty_1_106 <= _GEN_12060;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_107 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_107 <= _GEN_2038;
        end else begin
          dirty_1_107 <= _GEN_12061;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_108 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_108 <= _GEN_2039;
        end else begin
          dirty_1_108 <= _GEN_12062;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_109 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_109 <= _GEN_2040;
        end else begin
          dirty_1_109 <= _GEN_12063;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_110 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_110 <= _GEN_2041;
        end else begin
          dirty_1_110 <= _GEN_12064;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_111 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_111 <= _GEN_2042;
        end else begin
          dirty_1_111 <= _GEN_12065;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_112 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_112 <= _GEN_2043;
        end else begin
          dirty_1_112 <= _GEN_12066;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_113 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_113 <= _GEN_2044;
        end else begin
          dirty_1_113 <= _GEN_12067;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_114 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_114 <= _GEN_2045;
        end else begin
          dirty_1_114 <= _GEN_12068;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_115 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_115 <= _GEN_2046;
        end else begin
          dirty_1_115 <= _GEN_12069;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_116 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_116 <= _GEN_2047;
        end else begin
          dirty_1_116 <= _GEN_12070;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_117 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_117 <= _GEN_2048;
        end else begin
          dirty_1_117 <= _GEN_12071;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_118 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_118 <= _GEN_2049;
        end else begin
          dirty_1_118 <= _GEN_12072;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_119 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_119 <= _GEN_2050;
        end else begin
          dirty_1_119 <= _GEN_12073;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_120 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_120 <= _GEN_2051;
        end else begin
          dirty_1_120 <= _GEN_12074;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_121 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_121 <= _GEN_2052;
        end else begin
          dirty_1_121 <= _GEN_12075;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_122 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_122 <= _GEN_2053;
        end else begin
          dirty_1_122 <= _GEN_12076;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_123 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_123 <= _GEN_2054;
        end else begin
          dirty_1_123 <= _GEN_12077;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_124 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_124 <= _GEN_2055;
        end else begin
          dirty_1_124 <= _GEN_12078;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_125 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_125 <= _GEN_2056;
        end else begin
          dirty_1_125 <= _GEN_12079;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_126 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_126 <= _GEN_2057;
        end else begin
          dirty_1_126 <= _GEN_12080;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_127 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (3'h2 == state) begin // @[d_cache.scala 64:18]
          dirty_1_127 <= _GEN_2058;
        end else begin
          dirty_1_127 <= _GEN_12081;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:27]
      way0_hit <= 1'h0; // @[d_cache.scala 26:27]
    end else begin
      way0_hit <= _T_4;
    end
    if (reset) begin // @[d_cache.scala 27:27]
      way1_hit <= 1'h0; // @[d_cache.scala 27:27]
    end else begin
      way1_hit <= _T_7;
    end
    if (reset) begin // @[d_cache.scala 29:34]
      write_back_data <= 64'h0; // @[d_cache.scala 29:34]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          write_back_data <= _GEN_11824;
        end
      end
    end
    write_back_addr <= _GEN_16293[31:0]; // @[d_cache.scala 30:{34,34}]
    if (reset) begin // @[d_cache.scala 33:28]
      unuse_way <= 2'h0; // @[d_cache.scala 33:28]
    end else if (~_GEN_255) begin // @[d_cache.scala 52:31]
      unuse_way <= 2'h1; // @[d_cache.scala 53:19]
    end else if (~_GEN_512) begin // @[d_cache.scala 54:37]
      unuse_way <= 2'h2; // @[d_cache.scala 55:19]
    end else begin
      unuse_way <= 2'h0; // @[d_cache.scala 57:19]
    end
    if (reset) begin // @[d_cache.scala 34:31]
      receive_data <= 64'h0; // @[d_cache.scala 34:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          receive_data <= _GEN_11054;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:24]
      quene <= 1'h0; // @[d_cache.scala 35:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 64:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 64:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 64:18]
          quene <= _GEN_11439;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 60:24]
      state <= 3'h0; // @[d_cache.scala 60:24]
    end else if (3'h0 == state) begin // @[d_cache.scala 64:18]
      if (io_from_lsu_arvalid) begin // @[d_cache.scala 66:38]
        state <= 3'h1; // @[d_cache.scala 67:23]
      end else if (io_from_lsu_awvalid) begin // @[d_cache.scala 68:44]
        state <= 3'h2; // @[d_cache.scala 69:23]
      end
    end else if (3'h1 == state) begin // @[d_cache.scala 64:18]
      if (way0_hit) begin // @[d_cache.scala 74:27]
        state <= _GEN_646;
      end else begin
        state <= _GEN_775;
      end
    end else if (3'h2 == state) begin // @[d_cache.scala 64:18]
      state <= _GEN_1546;
    end else begin
      state <= _GEN_11053;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"read addr : %x  write addr : %x\n",io_from_lsu_araddr,io_from_lsu_awaddr); // @[d_cache.scala 15:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"d_cache state:%d\n",state); // @[d_cache.scala 61:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"bvalid:%d\n",io_from_axi_bvalid); // @[d_cache.scala 62:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"receive data:%x\n",receive_data); // @[d_cache.scala 63:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_16 & _T_17 & way0_hit & io_from_lsu_rready & _T_1) begin
          $fwrite(32'h80000002,"dirty_0:%d\n",7'h7f == index ? dirty_0_127 : _GEN_644); // @[d_cache.scala 76:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_16295 & ~way0_hit & way1_hit & io_from_lsu_rready & _T_1) begin
          $fwrite(32'h80000002,"dirty_1:%d\n",7'h7f == index ? dirty_1_127 : _GEN_773); // @[d_cache.scala 82:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"to lsu rdata:%x\n",io_to_lsu_rdata); // @[d_cache.scala 341:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"cacheline0:%x   cacheline1:%x\n",_GEN_2957,_GEN_4497); // @[d_cache.scala 342:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ram_0_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ram_0_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ram_0_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ram_0_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ram_0_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ram_0_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ram_0_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ram_0_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  ram_0_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  ram_0_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  ram_0_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  ram_0_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  ram_0_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  ram_0_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  ram_0_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  ram_0_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  ram_0_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  ram_0_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  ram_0_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  ram_0_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  ram_0_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  ram_0_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  ram_0_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  ram_0_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  ram_0_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  ram_0_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  ram_0_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  ram_0_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  ram_0_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  ram_0_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  ram_0_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  ram_0_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  ram_0_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  ram_0_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  ram_0_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  ram_0_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  ram_0_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  ram_0_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  ram_0_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  ram_0_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  ram_0_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  ram_0_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  ram_0_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  ram_0_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  ram_0_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  ram_0_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  ram_0_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  ram_0_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  ram_0_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  ram_0_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  ram_0_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  ram_0_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  ram_0_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  ram_0_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  ram_0_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  ram_0_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  ram_0_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  ram_0_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  ram_0_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  ram_0_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  ram_0_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  ram_0_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  ram_0_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  ram_0_63 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  ram_0_64 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  ram_0_65 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  ram_0_66 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  ram_0_67 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  ram_0_68 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  ram_0_69 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  ram_0_70 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  ram_0_71 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  ram_0_72 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  ram_0_73 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  ram_0_74 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  ram_0_75 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  ram_0_76 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  ram_0_77 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  ram_0_78 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  ram_0_79 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  ram_0_80 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  ram_0_81 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  ram_0_82 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  ram_0_83 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  ram_0_84 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  ram_0_85 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  ram_0_86 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  ram_0_87 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  ram_0_88 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  ram_0_89 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  ram_0_90 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  ram_0_91 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  ram_0_92 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  ram_0_93 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  ram_0_94 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  ram_0_95 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  ram_0_96 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  ram_0_97 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  ram_0_98 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  ram_0_99 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  ram_0_100 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  ram_0_101 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  ram_0_102 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  ram_0_103 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  ram_0_104 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  ram_0_105 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  ram_0_106 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  ram_0_107 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  ram_0_108 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  ram_0_109 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  ram_0_110 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  ram_0_111 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  ram_0_112 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  ram_0_113 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  ram_0_114 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  ram_0_115 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  ram_0_116 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  ram_0_117 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  ram_0_118 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  ram_0_119 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  ram_0_120 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  ram_0_121 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  ram_0_122 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  ram_0_123 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  ram_0_124 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  ram_0_125 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  ram_0_126 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  ram_0_127 = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  ram_1_0 = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  ram_1_1 = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  ram_1_2 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  ram_1_3 = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  ram_1_4 = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  ram_1_5 = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  ram_1_6 = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  ram_1_7 = _RAND_135[63:0];
  _RAND_136 = {2{`RANDOM}};
  ram_1_8 = _RAND_136[63:0];
  _RAND_137 = {2{`RANDOM}};
  ram_1_9 = _RAND_137[63:0];
  _RAND_138 = {2{`RANDOM}};
  ram_1_10 = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  ram_1_11 = _RAND_139[63:0];
  _RAND_140 = {2{`RANDOM}};
  ram_1_12 = _RAND_140[63:0];
  _RAND_141 = {2{`RANDOM}};
  ram_1_13 = _RAND_141[63:0];
  _RAND_142 = {2{`RANDOM}};
  ram_1_14 = _RAND_142[63:0];
  _RAND_143 = {2{`RANDOM}};
  ram_1_15 = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  ram_1_16 = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  ram_1_17 = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  ram_1_18 = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  ram_1_19 = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  ram_1_20 = _RAND_148[63:0];
  _RAND_149 = {2{`RANDOM}};
  ram_1_21 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  ram_1_22 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  ram_1_23 = _RAND_151[63:0];
  _RAND_152 = {2{`RANDOM}};
  ram_1_24 = _RAND_152[63:0];
  _RAND_153 = {2{`RANDOM}};
  ram_1_25 = _RAND_153[63:0];
  _RAND_154 = {2{`RANDOM}};
  ram_1_26 = _RAND_154[63:0];
  _RAND_155 = {2{`RANDOM}};
  ram_1_27 = _RAND_155[63:0];
  _RAND_156 = {2{`RANDOM}};
  ram_1_28 = _RAND_156[63:0];
  _RAND_157 = {2{`RANDOM}};
  ram_1_29 = _RAND_157[63:0];
  _RAND_158 = {2{`RANDOM}};
  ram_1_30 = _RAND_158[63:0];
  _RAND_159 = {2{`RANDOM}};
  ram_1_31 = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  ram_1_32 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  ram_1_33 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  ram_1_34 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  ram_1_35 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  ram_1_36 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  ram_1_37 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  ram_1_38 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  ram_1_39 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  ram_1_40 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  ram_1_41 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  ram_1_42 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  ram_1_43 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  ram_1_44 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  ram_1_45 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  ram_1_46 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  ram_1_47 = _RAND_175[63:0];
  _RAND_176 = {2{`RANDOM}};
  ram_1_48 = _RAND_176[63:0];
  _RAND_177 = {2{`RANDOM}};
  ram_1_49 = _RAND_177[63:0];
  _RAND_178 = {2{`RANDOM}};
  ram_1_50 = _RAND_178[63:0];
  _RAND_179 = {2{`RANDOM}};
  ram_1_51 = _RAND_179[63:0];
  _RAND_180 = {2{`RANDOM}};
  ram_1_52 = _RAND_180[63:0];
  _RAND_181 = {2{`RANDOM}};
  ram_1_53 = _RAND_181[63:0];
  _RAND_182 = {2{`RANDOM}};
  ram_1_54 = _RAND_182[63:0];
  _RAND_183 = {2{`RANDOM}};
  ram_1_55 = _RAND_183[63:0];
  _RAND_184 = {2{`RANDOM}};
  ram_1_56 = _RAND_184[63:0];
  _RAND_185 = {2{`RANDOM}};
  ram_1_57 = _RAND_185[63:0];
  _RAND_186 = {2{`RANDOM}};
  ram_1_58 = _RAND_186[63:0];
  _RAND_187 = {2{`RANDOM}};
  ram_1_59 = _RAND_187[63:0];
  _RAND_188 = {2{`RANDOM}};
  ram_1_60 = _RAND_188[63:0];
  _RAND_189 = {2{`RANDOM}};
  ram_1_61 = _RAND_189[63:0];
  _RAND_190 = {2{`RANDOM}};
  ram_1_62 = _RAND_190[63:0];
  _RAND_191 = {2{`RANDOM}};
  ram_1_63 = _RAND_191[63:0];
  _RAND_192 = {2{`RANDOM}};
  ram_1_64 = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  ram_1_65 = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  ram_1_66 = _RAND_194[63:0];
  _RAND_195 = {2{`RANDOM}};
  ram_1_67 = _RAND_195[63:0];
  _RAND_196 = {2{`RANDOM}};
  ram_1_68 = _RAND_196[63:0];
  _RAND_197 = {2{`RANDOM}};
  ram_1_69 = _RAND_197[63:0];
  _RAND_198 = {2{`RANDOM}};
  ram_1_70 = _RAND_198[63:0];
  _RAND_199 = {2{`RANDOM}};
  ram_1_71 = _RAND_199[63:0];
  _RAND_200 = {2{`RANDOM}};
  ram_1_72 = _RAND_200[63:0];
  _RAND_201 = {2{`RANDOM}};
  ram_1_73 = _RAND_201[63:0];
  _RAND_202 = {2{`RANDOM}};
  ram_1_74 = _RAND_202[63:0];
  _RAND_203 = {2{`RANDOM}};
  ram_1_75 = _RAND_203[63:0];
  _RAND_204 = {2{`RANDOM}};
  ram_1_76 = _RAND_204[63:0];
  _RAND_205 = {2{`RANDOM}};
  ram_1_77 = _RAND_205[63:0];
  _RAND_206 = {2{`RANDOM}};
  ram_1_78 = _RAND_206[63:0];
  _RAND_207 = {2{`RANDOM}};
  ram_1_79 = _RAND_207[63:0];
  _RAND_208 = {2{`RANDOM}};
  ram_1_80 = _RAND_208[63:0];
  _RAND_209 = {2{`RANDOM}};
  ram_1_81 = _RAND_209[63:0];
  _RAND_210 = {2{`RANDOM}};
  ram_1_82 = _RAND_210[63:0];
  _RAND_211 = {2{`RANDOM}};
  ram_1_83 = _RAND_211[63:0];
  _RAND_212 = {2{`RANDOM}};
  ram_1_84 = _RAND_212[63:0];
  _RAND_213 = {2{`RANDOM}};
  ram_1_85 = _RAND_213[63:0];
  _RAND_214 = {2{`RANDOM}};
  ram_1_86 = _RAND_214[63:0];
  _RAND_215 = {2{`RANDOM}};
  ram_1_87 = _RAND_215[63:0];
  _RAND_216 = {2{`RANDOM}};
  ram_1_88 = _RAND_216[63:0];
  _RAND_217 = {2{`RANDOM}};
  ram_1_89 = _RAND_217[63:0];
  _RAND_218 = {2{`RANDOM}};
  ram_1_90 = _RAND_218[63:0];
  _RAND_219 = {2{`RANDOM}};
  ram_1_91 = _RAND_219[63:0];
  _RAND_220 = {2{`RANDOM}};
  ram_1_92 = _RAND_220[63:0];
  _RAND_221 = {2{`RANDOM}};
  ram_1_93 = _RAND_221[63:0];
  _RAND_222 = {2{`RANDOM}};
  ram_1_94 = _RAND_222[63:0];
  _RAND_223 = {2{`RANDOM}};
  ram_1_95 = _RAND_223[63:0];
  _RAND_224 = {2{`RANDOM}};
  ram_1_96 = _RAND_224[63:0];
  _RAND_225 = {2{`RANDOM}};
  ram_1_97 = _RAND_225[63:0];
  _RAND_226 = {2{`RANDOM}};
  ram_1_98 = _RAND_226[63:0];
  _RAND_227 = {2{`RANDOM}};
  ram_1_99 = _RAND_227[63:0];
  _RAND_228 = {2{`RANDOM}};
  ram_1_100 = _RAND_228[63:0];
  _RAND_229 = {2{`RANDOM}};
  ram_1_101 = _RAND_229[63:0];
  _RAND_230 = {2{`RANDOM}};
  ram_1_102 = _RAND_230[63:0];
  _RAND_231 = {2{`RANDOM}};
  ram_1_103 = _RAND_231[63:0];
  _RAND_232 = {2{`RANDOM}};
  ram_1_104 = _RAND_232[63:0];
  _RAND_233 = {2{`RANDOM}};
  ram_1_105 = _RAND_233[63:0];
  _RAND_234 = {2{`RANDOM}};
  ram_1_106 = _RAND_234[63:0];
  _RAND_235 = {2{`RANDOM}};
  ram_1_107 = _RAND_235[63:0];
  _RAND_236 = {2{`RANDOM}};
  ram_1_108 = _RAND_236[63:0];
  _RAND_237 = {2{`RANDOM}};
  ram_1_109 = _RAND_237[63:0];
  _RAND_238 = {2{`RANDOM}};
  ram_1_110 = _RAND_238[63:0];
  _RAND_239 = {2{`RANDOM}};
  ram_1_111 = _RAND_239[63:0];
  _RAND_240 = {2{`RANDOM}};
  ram_1_112 = _RAND_240[63:0];
  _RAND_241 = {2{`RANDOM}};
  ram_1_113 = _RAND_241[63:0];
  _RAND_242 = {2{`RANDOM}};
  ram_1_114 = _RAND_242[63:0];
  _RAND_243 = {2{`RANDOM}};
  ram_1_115 = _RAND_243[63:0];
  _RAND_244 = {2{`RANDOM}};
  ram_1_116 = _RAND_244[63:0];
  _RAND_245 = {2{`RANDOM}};
  ram_1_117 = _RAND_245[63:0];
  _RAND_246 = {2{`RANDOM}};
  ram_1_118 = _RAND_246[63:0];
  _RAND_247 = {2{`RANDOM}};
  ram_1_119 = _RAND_247[63:0];
  _RAND_248 = {2{`RANDOM}};
  ram_1_120 = _RAND_248[63:0];
  _RAND_249 = {2{`RANDOM}};
  ram_1_121 = _RAND_249[63:0];
  _RAND_250 = {2{`RANDOM}};
  ram_1_122 = _RAND_250[63:0];
  _RAND_251 = {2{`RANDOM}};
  ram_1_123 = _RAND_251[63:0];
  _RAND_252 = {2{`RANDOM}};
  ram_1_124 = _RAND_252[63:0];
  _RAND_253 = {2{`RANDOM}};
  ram_1_125 = _RAND_253[63:0];
  _RAND_254 = {2{`RANDOM}};
  ram_1_126 = _RAND_254[63:0];
  _RAND_255 = {2{`RANDOM}};
  ram_1_127 = _RAND_255[63:0];
  _RAND_256 = {1{`RANDOM}};
  tag_0_0 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  tag_0_1 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  tag_0_2 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  tag_0_3 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  tag_0_4 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  tag_0_5 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  tag_0_6 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  tag_0_7 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  tag_0_8 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  tag_0_9 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  tag_0_10 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  tag_0_11 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  tag_0_12 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  tag_0_13 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  tag_0_14 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  tag_0_15 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  tag_0_16 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  tag_0_17 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  tag_0_18 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  tag_0_19 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  tag_0_20 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  tag_0_21 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  tag_0_22 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  tag_0_23 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  tag_0_24 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  tag_0_25 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  tag_0_26 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  tag_0_27 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  tag_0_28 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  tag_0_29 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  tag_0_30 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  tag_0_31 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  tag_0_32 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  tag_0_33 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  tag_0_34 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  tag_0_35 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  tag_0_36 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  tag_0_37 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  tag_0_38 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  tag_0_39 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  tag_0_40 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  tag_0_41 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  tag_0_42 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  tag_0_43 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  tag_0_44 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  tag_0_45 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  tag_0_46 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  tag_0_47 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  tag_0_48 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  tag_0_49 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  tag_0_50 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  tag_0_51 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  tag_0_52 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  tag_0_53 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  tag_0_54 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  tag_0_55 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  tag_0_56 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  tag_0_57 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  tag_0_58 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  tag_0_59 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  tag_0_60 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  tag_0_61 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  tag_0_62 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  tag_0_63 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  tag_0_64 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  tag_0_65 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  tag_0_66 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  tag_0_67 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  tag_0_68 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  tag_0_69 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  tag_0_70 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  tag_0_71 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  tag_0_72 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  tag_0_73 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  tag_0_74 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  tag_0_75 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  tag_0_76 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  tag_0_77 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  tag_0_78 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  tag_0_79 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  tag_0_80 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  tag_0_81 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  tag_0_82 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  tag_0_83 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  tag_0_84 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  tag_0_85 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  tag_0_86 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  tag_0_87 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  tag_0_88 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  tag_0_89 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  tag_0_90 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  tag_0_91 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  tag_0_92 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  tag_0_93 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  tag_0_94 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  tag_0_95 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  tag_0_96 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  tag_0_97 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  tag_0_98 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  tag_0_99 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  tag_0_100 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  tag_0_101 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  tag_0_102 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  tag_0_103 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  tag_0_104 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  tag_0_105 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  tag_0_106 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  tag_0_107 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  tag_0_108 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  tag_0_109 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  tag_0_110 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  tag_0_111 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  tag_0_112 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  tag_0_113 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  tag_0_114 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  tag_0_115 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  tag_0_116 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  tag_0_117 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  tag_0_118 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  tag_0_119 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  tag_0_120 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  tag_0_121 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  tag_0_122 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  tag_0_123 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  tag_0_124 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  tag_0_125 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  tag_0_126 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  tag_0_127 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  tag_1_0 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  tag_1_1 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  tag_1_2 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  tag_1_3 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  tag_1_4 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  tag_1_5 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  tag_1_6 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  tag_1_7 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  tag_1_8 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  tag_1_9 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  tag_1_10 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  tag_1_11 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  tag_1_12 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  tag_1_13 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  tag_1_14 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  tag_1_15 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  tag_1_16 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  tag_1_17 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  tag_1_18 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  tag_1_19 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  tag_1_20 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  tag_1_21 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  tag_1_22 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  tag_1_23 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  tag_1_24 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  tag_1_25 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  tag_1_26 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  tag_1_27 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  tag_1_28 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  tag_1_29 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  tag_1_30 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  tag_1_31 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  tag_1_32 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  tag_1_33 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  tag_1_34 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  tag_1_35 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  tag_1_36 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  tag_1_37 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  tag_1_38 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  tag_1_39 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  tag_1_40 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  tag_1_41 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  tag_1_42 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  tag_1_43 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  tag_1_44 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  tag_1_45 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  tag_1_46 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  tag_1_47 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  tag_1_48 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  tag_1_49 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  tag_1_50 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  tag_1_51 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  tag_1_52 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  tag_1_53 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  tag_1_54 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  tag_1_55 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  tag_1_56 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  tag_1_57 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  tag_1_58 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  tag_1_59 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  tag_1_60 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  tag_1_61 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  tag_1_62 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  tag_1_63 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  tag_1_64 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  tag_1_65 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  tag_1_66 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  tag_1_67 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  tag_1_68 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  tag_1_69 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  tag_1_70 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  tag_1_71 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  tag_1_72 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  tag_1_73 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  tag_1_74 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  tag_1_75 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  tag_1_76 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  tag_1_77 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  tag_1_78 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  tag_1_79 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  tag_1_80 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  tag_1_81 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  tag_1_82 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  tag_1_83 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  tag_1_84 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  tag_1_85 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  tag_1_86 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  tag_1_87 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  tag_1_88 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  tag_1_89 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  tag_1_90 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  tag_1_91 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  tag_1_92 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  tag_1_93 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  tag_1_94 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  tag_1_95 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  tag_1_96 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  tag_1_97 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  tag_1_98 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  tag_1_99 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  tag_1_100 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  tag_1_101 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  tag_1_102 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  tag_1_103 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  tag_1_104 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  tag_1_105 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  tag_1_106 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  tag_1_107 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  tag_1_108 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  tag_1_109 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  tag_1_110 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  tag_1_111 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  tag_1_112 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  tag_1_113 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  tag_1_114 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  tag_1_115 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  tag_1_116 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  tag_1_117 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  tag_1_118 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  tag_1_119 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  tag_1_120 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  tag_1_121 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  tag_1_122 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  tag_1_123 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  tag_1_124 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  tag_1_125 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  tag_1_126 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  tag_1_127 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  valid_0_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid_0_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  valid_0_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  valid_0_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  valid_0_4 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  valid_0_5 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  valid_0_6 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  valid_0_7 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  valid_0_8 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  valid_0_9 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  valid_0_10 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  valid_0_11 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  valid_0_12 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  valid_0_13 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  valid_0_14 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  valid_0_15 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  valid_0_16 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  valid_0_17 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  valid_0_18 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  valid_0_19 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  valid_0_20 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  valid_0_21 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  valid_0_22 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  valid_0_23 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  valid_0_24 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  valid_0_25 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  valid_0_26 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  valid_0_27 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  valid_0_28 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  valid_0_29 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  valid_0_30 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  valid_0_31 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  valid_0_32 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  valid_0_33 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  valid_0_34 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  valid_0_35 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  valid_0_36 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  valid_0_37 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  valid_0_38 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  valid_0_39 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  valid_0_40 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  valid_0_41 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  valid_0_42 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  valid_0_43 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  valid_0_44 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  valid_0_45 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  valid_0_46 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  valid_0_47 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  valid_0_48 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  valid_0_49 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  valid_0_50 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  valid_0_51 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  valid_0_52 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  valid_0_53 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  valid_0_54 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  valid_0_55 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  valid_0_56 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  valid_0_57 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  valid_0_58 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  valid_0_59 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  valid_0_60 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  valid_0_61 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  valid_0_62 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  valid_0_63 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  valid_0_64 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  valid_0_65 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  valid_0_66 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  valid_0_67 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  valid_0_68 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  valid_0_69 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  valid_0_70 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  valid_0_71 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  valid_0_72 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  valid_0_73 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  valid_0_74 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  valid_0_75 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  valid_0_76 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  valid_0_77 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  valid_0_78 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  valid_0_79 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  valid_0_80 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  valid_0_81 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  valid_0_82 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  valid_0_83 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  valid_0_84 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  valid_0_85 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  valid_0_86 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  valid_0_87 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  valid_0_88 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  valid_0_89 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  valid_0_90 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  valid_0_91 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  valid_0_92 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  valid_0_93 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  valid_0_94 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  valid_0_95 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  valid_0_96 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  valid_0_97 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  valid_0_98 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  valid_0_99 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  valid_0_100 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  valid_0_101 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  valid_0_102 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  valid_0_103 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  valid_0_104 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  valid_0_105 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  valid_0_106 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  valid_0_107 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  valid_0_108 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  valid_0_109 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  valid_0_110 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  valid_0_111 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  valid_0_112 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  valid_0_113 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  valid_0_114 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  valid_0_115 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  valid_0_116 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  valid_0_117 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  valid_0_118 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  valid_0_119 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  valid_0_120 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  valid_0_121 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  valid_0_122 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  valid_0_123 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  valid_0_124 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  valid_0_125 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  valid_0_126 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  valid_0_127 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  valid_1_0 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  valid_1_1 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  valid_1_2 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  valid_1_3 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  valid_1_4 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  valid_1_5 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  valid_1_6 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  valid_1_7 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  valid_1_8 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  valid_1_9 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  valid_1_10 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  valid_1_11 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  valid_1_12 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  valid_1_13 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  valid_1_14 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  valid_1_15 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  valid_1_16 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  valid_1_17 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  valid_1_18 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  valid_1_19 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  valid_1_20 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  valid_1_21 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  valid_1_22 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  valid_1_23 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  valid_1_24 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  valid_1_25 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  valid_1_26 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  valid_1_27 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  valid_1_28 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  valid_1_29 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  valid_1_30 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  valid_1_31 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  valid_1_32 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  valid_1_33 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  valid_1_34 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  valid_1_35 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  valid_1_36 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  valid_1_37 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  valid_1_38 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  valid_1_39 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  valid_1_40 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  valid_1_41 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  valid_1_42 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  valid_1_43 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  valid_1_44 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  valid_1_45 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  valid_1_46 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  valid_1_47 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  valid_1_48 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  valid_1_49 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  valid_1_50 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  valid_1_51 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  valid_1_52 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  valid_1_53 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  valid_1_54 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  valid_1_55 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  valid_1_56 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  valid_1_57 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  valid_1_58 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  valid_1_59 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  valid_1_60 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  valid_1_61 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  valid_1_62 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  valid_1_63 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  valid_1_64 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  valid_1_65 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  valid_1_66 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  valid_1_67 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  valid_1_68 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  valid_1_69 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  valid_1_70 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  valid_1_71 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  valid_1_72 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  valid_1_73 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  valid_1_74 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  valid_1_75 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  valid_1_76 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  valid_1_77 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  valid_1_78 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  valid_1_79 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  valid_1_80 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  valid_1_81 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  valid_1_82 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  valid_1_83 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  valid_1_84 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  valid_1_85 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  valid_1_86 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  valid_1_87 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  valid_1_88 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  valid_1_89 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  valid_1_90 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  valid_1_91 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  valid_1_92 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  valid_1_93 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  valid_1_94 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  valid_1_95 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  valid_1_96 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  valid_1_97 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  valid_1_98 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  valid_1_99 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  valid_1_100 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  valid_1_101 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  valid_1_102 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  valid_1_103 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  valid_1_104 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  valid_1_105 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  valid_1_106 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  valid_1_107 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  valid_1_108 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  valid_1_109 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  valid_1_110 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  valid_1_111 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  valid_1_112 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  valid_1_113 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  valid_1_114 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  valid_1_115 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  valid_1_116 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  valid_1_117 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  valid_1_118 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  valid_1_119 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  valid_1_120 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  valid_1_121 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  valid_1_122 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  valid_1_123 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  valid_1_124 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  valid_1_125 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  valid_1_126 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  valid_1_127 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  dirty_0_0 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  dirty_0_1 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  dirty_0_2 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  dirty_0_3 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  dirty_0_4 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  dirty_0_5 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  dirty_0_6 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  dirty_0_7 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  dirty_0_8 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  dirty_0_9 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  dirty_0_10 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  dirty_0_11 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  dirty_0_12 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  dirty_0_13 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  dirty_0_14 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  dirty_0_15 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  dirty_0_16 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  dirty_0_17 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  dirty_0_18 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  dirty_0_19 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  dirty_0_20 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  dirty_0_21 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  dirty_0_22 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  dirty_0_23 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  dirty_0_24 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  dirty_0_25 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  dirty_0_26 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  dirty_0_27 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  dirty_0_28 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  dirty_0_29 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  dirty_0_30 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  dirty_0_31 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  dirty_0_32 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  dirty_0_33 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  dirty_0_34 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  dirty_0_35 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  dirty_0_36 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  dirty_0_37 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  dirty_0_38 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  dirty_0_39 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  dirty_0_40 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  dirty_0_41 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  dirty_0_42 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  dirty_0_43 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  dirty_0_44 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  dirty_0_45 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  dirty_0_46 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  dirty_0_47 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  dirty_0_48 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  dirty_0_49 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  dirty_0_50 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  dirty_0_51 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  dirty_0_52 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  dirty_0_53 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  dirty_0_54 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  dirty_0_55 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  dirty_0_56 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  dirty_0_57 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  dirty_0_58 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  dirty_0_59 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  dirty_0_60 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  dirty_0_61 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  dirty_0_62 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  dirty_0_63 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  dirty_0_64 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  dirty_0_65 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  dirty_0_66 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  dirty_0_67 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  dirty_0_68 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  dirty_0_69 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  dirty_0_70 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  dirty_0_71 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  dirty_0_72 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  dirty_0_73 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  dirty_0_74 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  dirty_0_75 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  dirty_0_76 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  dirty_0_77 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  dirty_0_78 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  dirty_0_79 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  dirty_0_80 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  dirty_0_81 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  dirty_0_82 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  dirty_0_83 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  dirty_0_84 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  dirty_0_85 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  dirty_0_86 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  dirty_0_87 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  dirty_0_88 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  dirty_0_89 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  dirty_0_90 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  dirty_0_91 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  dirty_0_92 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  dirty_0_93 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  dirty_0_94 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  dirty_0_95 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  dirty_0_96 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  dirty_0_97 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  dirty_0_98 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  dirty_0_99 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  dirty_0_100 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  dirty_0_101 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  dirty_0_102 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  dirty_0_103 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  dirty_0_104 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  dirty_0_105 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  dirty_0_106 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  dirty_0_107 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  dirty_0_108 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  dirty_0_109 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  dirty_0_110 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  dirty_0_111 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  dirty_0_112 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  dirty_0_113 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  dirty_0_114 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  dirty_0_115 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  dirty_0_116 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  dirty_0_117 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  dirty_0_118 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  dirty_0_119 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  dirty_0_120 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  dirty_0_121 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  dirty_0_122 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  dirty_0_123 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  dirty_0_124 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  dirty_0_125 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  dirty_0_126 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  dirty_0_127 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  dirty_1_0 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  dirty_1_1 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  dirty_1_2 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  dirty_1_3 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  dirty_1_4 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  dirty_1_5 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  dirty_1_6 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  dirty_1_7 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  dirty_1_8 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  dirty_1_9 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  dirty_1_10 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  dirty_1_11 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  dirty_1_12 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  dirty_1_13 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  dirty_1_14 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  dirty_1_15 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  dirty_1_16 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  dirty_1_17 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  dirty_1_18 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  dirty_1_19 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  dirty_1_20 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  dirty_1_21 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  dirty_1_22 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  dirty_1_23 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  dirty_1_24 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  dirty_1_25 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  dirty_1_26 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  dirty_1_27 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  dirty_1_28 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  dirty_1_29 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  dirty_1_30 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  dirty_1_31 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  dirty_1_32 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  dirty_1_33 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  dirty_1_34 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  dirty_1_35 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  dirty_1_36 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  dirty_1_37 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  dirty_1_38 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  dirty_1_39 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  dirty_1_40 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  dirty_1_41 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  dirty_1_42 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  dirty_1_43 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  dirty_1_44 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  dirty_1_45 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  dirty_1_46 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  dirty_1_47 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  dirty_1_48 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  dirty_1_49 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  dirty_1_50 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  dirty_1_51 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  dirty_1_52 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  dirty_1_53 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  dirty_1_54 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  dirty_1_55 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  dirty_1_56 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  dirty_1_57 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  dirty_1_58 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  dirty_1_59 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  dirty_1_60 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  dirty_1_61 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  dirty_1_62 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  dirty_1_63 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  dirty_1_64 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  dirty_1_65 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  dirty_1_66 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  dirty_1_67 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  dirty_1_68 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  dirty_1_69 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  dirty_1_70 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  dirty_1_71 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  dirty_1_72 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  dirty_1_73 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  dirty_1_74 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  dirty_1_75 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  dirty_1_76 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  dirty_1_77 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  dirty_1_78 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  dirty_1_79 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  dirty_1_80 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  dirty_1_81 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  dirty_1_82 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  dirty_1_83 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  dirty_1_84 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  dirty_1_85 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  dirty_1_86 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  dirty_1_87 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  dirty_1_88 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  dirty_1_89 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  dirty_1_90 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  dirty_1_91 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  dirty_1_92 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  dirty_1_93 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  dirty_1_94 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  dirty_1_95 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  dirty_1_96 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  dirty_1_97 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  dirty_1_98 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  dirty_1_99 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  dirty_1_100 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  dirty_1_101 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  dirty_1_102 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  dirty_1_103 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  dirty_1_104 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  dirty_1_105 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  dirty_1_106 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  dirty_1_107 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  dirty_1_108 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  dirty_1_109 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  dirty_1_110 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  dirty_1_111 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  dirty_1_112 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  dirty_1_113 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  dirty_1_114 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  dirty_1_115 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  dirty_1_116 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  dirty_1_117 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  dirty_1_118 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  dirty_1_119 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  dirty_1_120 = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  dirty_1_121 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  dirty_1_122 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  dirty_1_123 = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  dirty_1_124 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  dirty_1_125 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  dirty_1_126 = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  dirty_1_127 = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  way0_hit = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  way1_hit = _RAND_1025[0:0];
  _RAND_1026 = {2{`RANDOM}};
  write_back_data = _RAND_1026[63:0];
  _RAND_1027 = {1{`RANDOM}};
  write_back_addr = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  unuse_way = _RAND_1028[1:0];
  _RAND_1029 = {2{`RANDOM}};
  receive_data = _RAND_1029[63:0];
  _RAND_1030 = {1{`RANDOM}};
  quene = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  state = _RAND_1031[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
