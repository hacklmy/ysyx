module D_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_lsu_araddr,
  input         io_from_lsu_arvalid,
  input  [31:0] io_from_lsu_awaddr,
  input         io_from_lsu_awvalid,
  input  [63:0] io_from_lsu_wdata,
  input  [7:0]  io_from_lsu_wstrb,
  input         io_from_lsu_wvalid,
  output [63:0] io_to_lsu_rdata,
  output        io_to_lsu_rvalid,
  output        io_to_lsu_bvalid,
  output [31:0] io_to_axi_araddr,
  output [7:0]  io_to_axi_arlen,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  output [31:0] io_to_axi_awaddr,
  output [7:0]  io_to_axi_awlen,
  output        io_to_axi_awvalid,
  output [63:0] io_to_axi_wdata,
  output [7:0]  io_to_axi_wstrb,
  output        io_to_axi_wvalid,
  output        io_to_axi_bready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rlast,
  input         io_from_axi_rvalid,
  input         io_from_axi_wready,
  input         io_from_axi_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [127:0] _RAND_27;
  reg [127:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [127:0] _RAND_33;
  reg [127:0] _RAND_34;
  reg [127:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [127:0] _RAND_38;
  reg [127:0] _RAND_39;
  reg [127:0] _RAND_40;
  reg [127:0] _RAND_41;
  reg [127:0] _RAND_42;
  reg [127:0] _RAND_43;
  reg [127:0] _RAND_44;
  reg [127:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [127:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [127:0] _RAND_50;
  reg [127:0] _RAND_51;
  reg [127:0] _RAND_52;
  reg [127:0] _RAND_53;
  reg [127:0] _RAND_54;
  reg [127:0] _RAND_55;
  reg [127:0] _RAND_56;
  reg [127:0] _RAND_57;
  reg [127:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [127:0] _RAND_61;
  reg [127:0] _RAND_62;
  reg [127:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [127:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] ram_0_0; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_1; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_2; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_3; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_4; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_5; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_6; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_7; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_8; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_9; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_10; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_11; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_12; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_13; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_14; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_15; // @[d_cache.scala 19:24]
  reg [127:0] ram_1_0; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_1; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_2; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_3; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_4; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_5; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_6; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_7; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_8; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_9; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_10; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_11; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_12; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_13; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_14; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_15; // @[d_cache.scala 20:24]
  reg [127:0] ram_2_0; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_1; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_2; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_3; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_4; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_5; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_6; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_7; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_8; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_9; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_10; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_11; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_12; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_13; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_14; // @[d_cache.scala 21:24]
  reg [127:0] ram_2_15; // @[d_cache.scala 21:24]
  reg [127:0] ram_3_0; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_1; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_2; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_3; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_4; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_5; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_6; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_7; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_8; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_9; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_10; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_11; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_12; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_13; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_14; // @[d_cache.scala 22:24]
  reg [127:0] ram_3_15; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_0; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_1; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_2; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_3; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_4; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_5; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_6; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_7; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_8; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_9; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_10; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_11; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_12; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_13; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_14; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_15; // @[d_cache.scala 24:24]
  reg [31:0] tag_1_0; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_1; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_2; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_3; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_4; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_5; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_6; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_7; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_8; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_9; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_10; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_11; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_12; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_13; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_14; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_15; // @[d_cache.scala 25:24]
  reg [31:0] tag_2_0; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_1; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_2; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_3; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_4; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_5; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_6; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_7; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_8; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_9; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_10; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_11; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_12; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_13; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_14; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_15; // @[d_cache.scala 26:24]
  reg [31:0] tag_3_0; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_1; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_2; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_3; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_4; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_5; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_6; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_7; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_8; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_9; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_10; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_11; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_12; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_13; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_14; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_15; // @[d_cache.scala 27:24]
  reg  valid_0_0; // @[d_cache.scala 28:26]
  reg  valid_0_1; // @[d_cache.scala 28:26]
  reg  valid_0_2; // @[d_cache.scala 28:26]
  reg  valid_0_3; // @[d_cache.scala 28:26]
  reg  valid_0_4; // @[d_cache.scala 28:26]
  reg  valid_0_5; // @[d_cache.scala 28:26]
  reg  valid_0_6; // @[d_cache.scala 28:26]
  reg  valid_0_7; // @[d_cache.scala 28:26]
  reg  valid_0_8; // @[d_cache.scala 28:26]
  reg  valid_0_9; // @[d_cache.scala 28:26]
  reg  valid_0_10; // @[d_cache.scala 28:26]
  reg  valid_0_11; // @[d_cache.scala 28:26]
  reg  valid_0_12; // @[d_cache.scala 28:26]
  reg  valid_0_13; // @[d_cache.scala 28:26]
  reg  valid_0_14; // @[d_cache.scala 28:26]
  reg  valid_0_15; // @[d_cache.scala 28:26]
  reg  valid_1_0; // @[d_cache.scala 29:26]
  reg  valid_1_1; // @[d_cache.scala 29:26]
  reg  valid_1_2; // @[d_cache.scala 29:26]
  reg  valid_1_3; // @[d_cache.scala 29:26]
  reg  valid_1_4; // @[d_cache.scala 29:26]
  reg  valid_1_5; // @[d_cache.scala 29:26]
  reg  valid_1_6; // @[d_cache.scala 29:26]
  reg  valid_1_7; // @[d_cache.scala 29:26]
  reg  valid_1_8; // @[d_cache.scala 29:26]
  reg  valid_1_9; // @[d_cache.scala 29:26]
  reg  valid_1_10; // @[d_cache.scala 29:26]
  reg  valid_1_11; // @[d_cache.scala 29:26]
  reg  valid_1_12; // @[d_cache.scala 29:26]
  reg  valid_1_13; // @[d_cache.scala 29:26]
  reg  valid_1_14; // @[d_cache.scala 29:26]
  reg  valid_1_15; // @[d_cache.scala 29:26]
  reg  valid_2_0; // @[d_cache.scala 30:26]
  reg  valid_2_1; // @[d_cache.scala 30:26]
  reg  valid_2_2; // @[d_cache.scala 30:26]
  reg  valid_2_3; // @[d_cache.scala 30:26]
  reg  valid_2_4; // @[d_cache.scala 30:26]
  reg  valid_2_5; // @[d_cache.scala 30:26]
  reg  valid_2_6; // @[d_cache.scala 30:26]
  reg  valid_2_7; // @[d_cache.scala 30:26]
  reg  valid_2_8; // @[d_cache.scala 30:26]
  reg  valid_2_9; // @[d_cache.scala 30:26]
  reg  valid_2_10; // @[d_cache.scala 30:26]
  reg  valid_2_11; // @[d_cache.scala 30:26]
  reg  valid_2_12; // @[d_cache.scala 30:26]
  reg  valid_2_13; // @[d_cache.scala 30:26]
  reg  valid_2_14; // @[d_cache.scala 30:26]
  reg  valid_2_15; // @[d_cache.scala 30:26]
  reg  valid_3_0; // @[d_cache.scala 31:26]
  reg  valid_3_1; // @[d_cache.scala 31:26]
  reg  valid_3_2; // @[d_cache.scala 31:26]
  reg  valid_3_3; // @[d_cache.scala 31:26]
  reg  valid_3_4; // @[d_cache.scala 31:26]
  reg  valid_3_5; // @[d_cache.scala 31:26]
  reg  valid_3_6; // @[d_cache.scala 31:26]
  reg  valid_3_7; // @[d_cache.scala 31:26]
  reg  valid_3_8; // @[d_cache.scala 31:26]
  reg  valid_3_9; // @[d_cache.scala 31:26]
  reg  valid_3_10; // @[d_cache.scala 31:26]
  reg  valid_3_11; // @[d_cache.scala 31:26]
  reg  valid_3_12; // @[d_cache.scala 31:26]
  reg  valid_3_13; // @[d_cache.scala 31:26]
  reg  valid_3_14; // @[d_cache.scala 31:26]
  reg  valid_3_15; // @[d_cache.scala 31:26]
  reg  dirty_0_0; // @[d_cache.scala 32:26]
  reg  dirty_0_1; // @[d_cache.scala 32:26]
  reg  dirty_0_2; // @[d_cache.scala 32:26]
  reg  dirty_0_3; // @[d_cache.scala 32:26]
  reg  dirty_0_4; // @[d_cache.scala 32:26]
  reg  dirty_0_5; // @[d_cache.scala 32:26]
  reg  dirty_0_6; // @[d_cache.scala 32:26]
  reg  dirty_0_7; // @[d_cache.scala 32:26]
  reg  dirty_0_8; // @[d_cache.scala 32:26]
  reg  dirty_0_9; // @[d_cache.scala 32:26]
  reg  dirty_0_10; // @[d_cache.scala 32:26]
  reg  dirty_0_11; // @[d_cache.scala 32:26]
  reg  dirty_0_12; // @[d_cache.scala 32:26]
  reg  dirty_0_13; // @[d_cache.scala 32:26]
  reg  dirty_0_14; // @[d_cache.scala 32:26]
  reg  dirty_0_15; // @[d_cache.scala 32:26]
  reg  dirty_3_0; // @[d_cache.scala 35:26]
  reg  dirty_3_1; // @[d_cache.scala 35:26]
  reg  dirty_3_2; // @[d_cache.scala 35:26]
  reg  dirty_3_3; // @[d_cache.scala 35:26]
  reg  dirty_3_4; // @[d_cache.scala 35:26]
  reg  dirty_3_5; // @[d_cache.scala 35:26]
  reg  dirty_3_6; // @[d_cache.scala 35:26]
  reg  dirty_3_7; // @[d_cache.scala 35:26]
  reg  dirty_3_8; // @[d_cache.scala 35:26]
  reg  dirty_3_9; // @[d_cache.scala 35:26]
  reg  dirty_3_10; // @[d_cache.scala 35:26]
  reg  dirty_3_11; // @[d_cache.scala 35:26]
  reg  dirty_3_12; // @[d_cache.scala 35:26]
  reg  dirty_3_13; // @[d_cache.scala 35:26]
  reg  dirty_3_14; // @[d_cache.scala 35:26]
  reg  dirty_3_15; // @[d_cache.scala 35:26]
  reg [127:0] write_back_data; // @[d_cache.scala 41:34]
  reg [31:0] write_back_addr; // @[d_cache.scala 42:34]
  reg [63:0] receive_data_0; // @[d_cache.scala 47:31]
  reg [63:0] receive_data_1; // @[d_cache.scala 47:31]
  reg [2:0] receive_num; // @[d_cache.scala 48:30]
  reg [7:0] quene_0; // @[d_cache.scala 49:24]
  reg [7:0] quene_1; // @[d_cache.scala 49:24]
  reg [7:0] quene_2; // @[d_cache.scala 49:24]
  reg [7:0] quene_3; // @[d_cache.scala 49:24]
  reg [7:0] quene_4; // @[d_cache.scala 49:24]
  reg [7:0] quene_5; // @[d_cache.scala 49:24]
  reg [7:0] quene_6; // @[d_cache.scala 49:24]
  reg [7:0] quene_7; // @[d_cache.scala 49:24]
  reg [7:0] quene_8; // @[d_cache.scala 49:24]
  reg [7:0] quene_9; // @[d_cache.scala 49:24]
  reg [7:0] quene_10; // @[d_cache.scala 49:24]
  reg [7:0] quene_11; // @[d_cache.scala 49:24]
  reg [7:0] quene_12; // @[d_cache.scala 49:24]
  reg [7:0] quene_13; // @[d_cache.scala 49:24]
  reg [7:0] quene_14; // @[d_cache.scala 49:24]
  reg [7:0] quene_15; // @[d_cache.scala 49:24]
  wire [3:0] offset = io_from_lsu_araddr[3:0]; // @[d_cache.scala 51:36]
  wire [3:0] index = io_from_lsu_araddr[7:4]; // @[d_cache.scala 52:35]
  wire [23:0] tag = io_from_lsu_araddr[31:8]; // @[d_cache.scala 53:33]
  wire [6:0] shift_bit = {offset, 3'h0}; // @[d_cache.scala 55:28]
  wire [63:0] _wmask_T_4 = io_from_lsu_wstrb == 8'hff ? 64'hffffffffffffffff : 64'h0; // @[d_cache.scala 61:20]
  wire [63:0] _wmask_T_5 = io_from_lsu_wstrb == 8'hf ? 64'hffffffff : _wmask_T_4; // @[d_cache.scala 60:20]
  wire [63:0] _wmask_T_6 = io_from_lsu_wstrb == 8'h3 ? 64'hffff : _wmask_T_5; // @[d_cache.scala 59:20]
  wire [63:0] wmask = io_from_lsu_wstrb == 8'h1 ? 64'hff : _wmask_T_6; // @[d_cache.scala 58:20]
  wire [31:0] _GEN_1 = 4'h1 == index ? tag_0_1 : tag_0_0; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_2 = 4'h2 == index ? tag_0_2 : _GEN_1; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_3 = 4'h3 == index ? tag_0_3 : _GEN_2; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_4 = 4'h4 == index ? tag_0_4 : _GEN_3; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_5 = 4'h5 == index ? tag_0_5 : _GEN_4; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_6 = 4'h6 == index ? tag_0_6 : _GEN_5; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_7 = 4'h7 == index ? tag_0_7 : _GEN_6; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_8 = 4'h8 == index ? tag_0_8 : _GEN_7; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_9 = 4'h9 == index ? tag_0_9 : _GEN_8; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_10 = 4'ha == index ? tag_0_10 : _GEN_9; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_11 = 4'hb == index ? tag_0_11 : _GEN_10; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_12 = 4'hc == index ? tag_0_12 : _GEN_11; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_13 = 4'hd == index ? tag_0_13 : _GEN_12; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_14 = 4'he == index ? tag_0_14 : _GEN_13; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_15 = 4'hf == index ? tag_0_15 : _GEN_14; // @[d_cache.scala 63:{31,31}]
  wire [31:0] _GEN_215 = {{8'd0}, tag}; // @[d_cache.scala 63:31]
  wire  _GEN_17 = 4'h1 == index ? valid_0_1 : valid_0_0; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_18 = 4'h2 == index ? valid_0_2 : _GEN_17; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_19 = 4'h3 == index ? valid_0_3 : _GEN_18; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_20 = 4'h4 == index ? valid_0_4 : _GEN_19; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_21 = 4'h5 == index ? valid_0_5 : _GEN_20; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_22 = 4'h6 == index ? valid_0_6 : _GEN_21; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_23 = 4'h7 == index ? valid_0_7 : _GEN_22; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_24 = 4'h8 == index ? valid_0_8 : _GEN_23; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_25 = 4'h9 == index ? valid_0_9 : _GEN_24; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_26 = 4'ha == index ? valid_0_10 : _GEN_25; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_27 = 4'hb == index ? valid_0_11 : _GEN_26; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_28 = 4'hc == index ? valid_0_12 : _GEN_27; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_29 = 4'hd == index ? valid_0_13 : _GEN_28; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_30 = 4'he == index ? valid_0_14 : _GEN_29; // @[d_cache.scala 63:{57,57}]
  wire  _GEN_31 = 4'hf == index ? valid_0_15 : _GEN_30; // @[d_cache.scala 63:{57,57}]
  wire  way0_hit = _GEN_15 == _GEN_215 & _GEN_31; // @[d_cache.scala 63:40]
  wire [31:0] _GEN_33 = 4'h1 == index ? tag_1_1 : tag_1_0; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_34 = 4'h2 == index ? tag_1_2 : _GEN_33; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_35 = 4'h3 == index ? tag_1_3 : _GEN_34; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_36 = 4'h4 == index ? tag_1_4 : _GEN_35; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_37 = 4'h5 == index ? tag_1_5 : _GEN_36; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_38 = 4'h6 == index ? tag_1_6 : _GEN_37; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_39 = 4'h7 == index ? tag_1_7 : _GEN_38; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_40 = 4'h8 == index ? tag_1_8 : _GEN_39; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_41 = 4'h9 == index ? tag_1_9 : _GEN_40; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_42 = 4'ha == index ? tag_1_10 : _GEN_41; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_43 = 4'hb == index ? tag_1_11 : _GEN_42; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_44 = 4'hc == index ? tag_1_12 : _GEN_43; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_45 = 4'hd == index ? tag_1_13 : _GEN_44; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_46 = 4'he == index ? tag_1_14 : _GEN_45; // @[d_cache.scala 65:{31,31}]
  wire [31:0] _GEN_47 = 4'hf == index ? tag_1_15 : _GEN_46; // @[d_cache.scala 65:{31,31}]
  wire  _GEN_49 = 4'h1 == index ? valid_1_1 : valid_1_0; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_50 = 4'h2 == index ? valid_1_2 : _GEN_49; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_51 = 4'h3 == index ? valid_1_3 : _GEN_50; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_52 = 4'h4 == index ? valid_1_4 : _GEN_51; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_53 = 4'h5 == index ? valid_1_5 : _GEN_52; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_54 = 4'h6 == index ? valid_1_6 : _GEN_53; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_55 = 4'h7 == index ? valid_1_7 : _GEN_54; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_56 = 4'h8 == index ? valid_1_8 : _GEN_55; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_57 = 4'h9 == index ? valid_1_9 : _GEN_56; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_58 = 4'ha == index ? valid_1_10 : _GEN_57; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_59 = 4'hb == index ? valid_1_11 : _GEN_58; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_60 = 4'hc == index ? valid_1_12 : _GEN_59; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_61 = 4'hd == index ? valid_1_13 : _GEN_60; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_62 = 4'he == index ? valid_1_14 : _GEN_61; // @[d_cache.scala 65:{57,57}]
  wire  _GEN_63 = 4'hf == index ? valid_1_15 : _GEN_62; // @[d_cache.scala 65:{57,57}]
  wire  way1_hit = _GEN_47 == _GEN_215 & _GEN_63; // @[d_cache.scala 65:40]
  wire [31:0] _GEN_65 = 4'h1 == index ? tag_2_1 : tag_2_0; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_66 = 4'h2 == index ? tag_2_2 : _GEN_65; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_67 = 4'h3 == index ? tag_2_3 : _GEN_66; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_68 = 4'h4 == index ? tag_2_4 : _GEN_67; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_69 = 4'h5 == index ? tag_2_5 : _GEN_68; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_70 = 4'h6 == index ? tag_2_6 : _GEN_69; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_71 = 4'h7 == index ? tag_2_7 : _GEN_70; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_72 = 4'h8 == index ? tag_2_8 : _GEN_71; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_73 = 4'h9 == index ? tag_2_9 : _GEN_72; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_74 = 4'ha == index ? tag_2_10 : _GEN_73; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_75 = 4'hb == index ? tag_2_11 : _GEN_74; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_76 = 4'hc == index ? tag_2_12 : _GEN_75; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_77 = 4'hd == index ? tag_2_13 : _GEN_76; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_78 = 4'he == index ? tag_2_14 : _GEN_77; // @[d_cache.scala 66:{31,31}]
  wire [31:0] _GEN_79 = 4'hf == index ? tag_2_15 : _GEN_78; // @[d_cache.scala 66:{31,31}]
  wire  _GEN_81 = 4'h1 == index ? valid_2_1 : valid_2_0; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_82 = 4'h2 == index ? valid_2_2 : _GEN_81; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_83 = 4'h3 == index ? valid_2_3 : _GEN_82; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_84 = 4'h4 == index ? valid_2_4 : _GEN_83; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_85 = 4'h5 == index ? valid_2_5 : _GEN_84; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_86 = 4'h6 == index ? valid_2_6 : _GEN_85; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_87 = 4'h7 == index ? valid_2_7 : _GEN_86; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_88 = 4'h8 == index ? valid_2_8 : _GEN_87; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_89 = 4'h9 == index ? valid_2_9 : _GEN_88; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_90 = 4'ha == index ? valid_2_10 : _GEN_89; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_91 = 4'hb == index ? valid_2_11 : _GEN_90; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_92 = 4'hc == index ? valid_2_12 : _GEN_91; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_93 = 4'hd == index ? valid_2_13 : _GEN_92; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_94 = 4'he == index ? valid_2_14 : _GEN_93; // @[d_cache.scala 66:{57,57}]
  wire  _GEN_95 = 4'hf == index ? valid_2_15 : _GEN_94; // @[d_cache.scala 66:{57,57}]
  wire  way2_hit = _GEN_79 == _GEN_215 & _GEN_95; // @[d_cache.scala 66:40]
  wire [31:0] _GEN_97 = 4'h1 == index ? tag_3_1 : tag_3_0; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_98 = 4'h2 == index ? tag_3_2 : _GEN_97; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_99 = 4'h3 == index ? tag_3_3 : _GEN_98; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_100 = 4'h4 == index ? tag_3_4 : _GEN_99; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_101 = 4'h5 == index ? tag_3_5 : _GEN_100; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_102 = 4'h6 == index ? tag_3_6 : _GEN_101; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_103 = 4'h7 == index ? tag_3_7 : _GEN_102; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_104 = 4'h8 == index ? tag_3_8 : _GEN_103; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_105 = 4'h9 == index ? tag_3_9 : _GEN_104; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_106 = 4'ha == index ? tag_3_10 : _GEN_105; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_107 = 4'hb == index ? tag_3_11 : _GEN_106; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_108 = 4'hc == index ? tag_3_12 : _GEN_107; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_109 = 4'hd == index ? tag_3_13 : _GEN_108; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_110 = 4'he == index ? tag_3_14 : _GEN_109; // @[d_cache.scala 67:{31,31}]
  wire [31:0] _GEN_111 = 4'hf == index ? tag_3_15 : _GEN_110; // @[d_cache.scala 67:{31,31}]
  wire  _GEN_113 = 4'h1 == index ? valid_3_1 : valid_3_0; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_114 = 4'h2 == index ? valid_3_2 : _GEN_113; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_115 = 4'h3 == index ? valid_3_3 : _GEN_114; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_116 = 4'h4 == index ? valid_3_4 : _GEN_115; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_117 = 4'h5 == index ? valid_3_5 : _GEN_116; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_118 = 4'h6 == index ? valid_3_6 : _GEN_117; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_119 = 4'h7 == index ? valid_3_7 : _GEN_118; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_120 = 4'h8 == index ? valid_3_8 : _GEN_119; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_121 = 4'h9 == index ? valid_3_9 : _GEN_120; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_122 = 4'ha == index ? valid_3_10 : _GEN_121; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_123 = 4'hb == index ? valid_3_11 : _GEN_122; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_124 = 4'hc == index ? valid_3_12 : _GEN_123; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_125 = 4'hd == index ? valid_3_13 : _GEN_124; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_126 = 4'he == index ? valid_3_14 : _GEN_125; // @[d_cache.scala 67:{57,57}]
  wire  _GEN_127 = 4'hf == index ? valid_3_15 : _GEN_126; // @[d_cache.scala 67:{57,57}]
  wire  way3_hit = _GEN_111 == _GEN_215 & _GEN_127; // @[d_cache.scala 67:40]
  wire [2:0] _unuse_way_T_4 = ~_GEN_127 ? 3'h4 : 3'h0; // @[d_cache.scala 69:108]
  wire [2:0] _unuse_way_T_5 = ~_GEN_95 ? 3'h3 : _unuse_way_T_4; // @[d_cache.scala 69:79]
  wire [2:0] _unuse_way_T_6 = ~_GEN_63 ? 3'h2 : _unuse_way_T_5; // @[d_cache.scala 69:50]
  wire [2:0] unuse_way = ~_GEN_31 ? 3'h1 : _unuse_way_T_6; // @[d_cache.scala 69:21]
  reg [3:0] state; // @[d_cache.scala 71:24]
  wire  _T_5 = (io_from_lsu_arvalid | io_from_lsu_awvalid) & io_from_lsu_araddr >= 32'ha0000000; // @[d_cache.scala 78:60]
  wire [3:0] _GEN_128 = io_from_lsu_awvalid ? 4'h2 : state; // @[d_cache.scala 82:44 83:23 71:24]
  wire  _T_9 = way0_hit | way1_hit | way2_hit | way3_hit; // @[d_cache.scala 87:46]
  wire [63:0] _ram_0_T = io_from_lsu_wdata & wmask; // @[d_cache.scala 101:53]
  wire [190:0] _GEN_1364 = {{127'd0}, _ram_0_T}; // @[d_cache.scala 101:62]
  wire [190:0] _ram_0_T_1 = _GEN_1364 << shift_bit; // @[d_cache.scala 101:62]
  wire [190:0] _GEN_1365 = {{127'd0}, wmask}; // @[d_cache.scala 101:102]
  wire [190:0] _ram_0_T_2 = _GEN_1365 << shift_bit; // @[d_cache.scala 101:102]
  wire [190:0] _ram_0_T_3 = ~_ram_0_T_2; // @[d_cache.scala 101:94]
  wire [127:0] _GEN_136 = 4'h1 == index ? ram_0_1 : ram_0_0; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_137 = 4'h2 == index ? ram_0_2 : _GEN_136; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_138 = 4'h3 == index ? ram_0_3 : _GEN_137; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_139 = 4'h4 == index ? ram_0_4 : _GEN_138; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_140 = 4'h5 == index ? ram_0_5 : _GEN_139; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_141 = 4'h6 == index ? ram_0_6 : _GEN_140; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_142 = 4'h7 == index ? ram_0_7 : _GEN_141; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_143 = 4'h8 == index ? ram_0_8 : _GEN_142; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_144 = 4'h9 == index ? ram_0_9 : _GEN_143; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_145 = 4'ha == index ? ram_0_10 : _GEN_144; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_146 = 4'hb == index ? ram_0_11 : _GEN_145; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_147 = 4'hc == index ? ram_0_12 : _GEN_146; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_148 = 4'hd == index ? ram_0_13 : _GEN_147; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_149 = 4'he == index ? ram_0_14 : _GEN_148; // @[d_cache.scala 101:{92,92}]
  wire [127:0] _GEN_150 = 4'hf == index ? ram_0_15 : _GEN_149; // @[d_cache.scala 101:{92,92}]
  wire [190:0] _GEN_219 = {{63'd0}, _GEN_150}; // @[d_cache.scala 101:92]
  wire [190:0] _ram_0_T_4 = _GEN_219 & _ram_0_T_3; // @[d_cache.scala 101:92]
  wire [190:0] _ram_0_T_5 = _ram_0_T_1 | _ram_0_T_4; // @[d_cache.scala 101:76]
  wire [127:0] _GEN_151 = 4'h0 == index ? _ram_0_T_5[127:0] : ram_0_0; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_152 = 4'h1 == index ? _ram_0_T_5[127:0] : ram_0_1; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_153 = 4'h2 == index ? _ram_0_T_5[127:0] : ram_0_2; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_154 = 4'h3 == index ? _ram_0_T_5[127:0] : ram_0_3; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_155 = 4'h4 == index ? _ram_0_T_5[127:0] : ram_0_4; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_156 = 4'h5 == index ? _ram_0_T_5[127:0] : ram_0_5; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_157 = 4'h6 == index ? _ram_0_T_5[127:0] : ram_0_6; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_158 = 4'h7 == index ? _ram_0_T_5[127:0] : ram_0_7; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_159 = 4'h8 == index ? _ram_0_T_5[127:0] : ram_0_8; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_160 = 4'h9 == index ? _ram_0_T_5[127:0] : ram_0_9; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_161 = 4'ha == index ? _ram_0_T_5[127:0] : ram_0_10; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_162 = 4'hb == index ? _ram_0_T_5[127:0] : ram_0_11; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_163 = 4'hc == index ? _ram_0_T_5[127:0] : ram_0_12; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_164 = 4'hd == index ? _ram_0_T_5[127:0] : ram_0_13; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_165 = 4'he == index ? _ram_0_T_5[127:0] : ram_0_14; // @[d_cache.scala 101:{30,30} 19:24]
  wire [127:0] _GEN_166 = 4'hf == index ? _ram_0_T_5[127:0] : ram_0_15; // @[d_cache.scala 101:{30,30} 19:24]
  wire  _GEN_220 = 4'h0 == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_167 = 4'h0 == index | dirty_0_0; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_221 = 4'h1 == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_168 = 4'h1 == index | dirty_0_1; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_222 = 4'h2 == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_169 = 4'h2 == index | dirty_0_2; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_223 = 4'h3 == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_170 = 4'h3 == index | dirty_0_3; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_224 = 4'h4 == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_171 = 4'h4 == index | dirty_0_4; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_225 = 4'h5 == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_172 = 4'h5 == index | dirty_0_5; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_226 = 4'h6 == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_173 = 4'h6 == index | dirty_0_6; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_227 = 4'h7 == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_174 = 4'h7 == index | dirty_0_7; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_228 = 4'h8 == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_175 = 4'h8 == index | dirty_0_8; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_229 = 4'h9 == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_176 = 4'h9 == index | dirty_0_9; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_230 = 4'ha == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_177 = 4'ha == index | dirty_0_10; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_263 = 4'hb == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_178 = 4'hb == index | dirty_0_11; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_264 = 4'hc == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_179 = 4'hc == index | dirty_0_12; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_265 = 4'hd == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_180 = 4'hd == index | dirty_0_13; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_266 = 4'he == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_181 = 4'he == index | dirty_0_14; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_267 = 4'hf == index; // @[d_cache.scala 102:{32,32} 32:26]
  wire  _GEN_182 = 4'hf == index | dirty_0_15; // @[d_cache.scala 102:{32,32} 32:26]
  wire [127:0] _GEN_184 = 4'h1 == index ? ram_1_1 : ram_1_0; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_185 = 4'h2 == index ? ram_1_2 : _GEN_184; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_186 = 4'h3 == index ? ram_1_3 : _GEN_185; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_187 = 4'h4 == index ? ram_1_4 : _GEN_186; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_188 = 4'h5 == index ? ram_1_5 : _GEN_187; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_189 = 4'h6 == index ? ram_1_6 : _GEN_188; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_190 = 4'h7 == index ? ram_1_7 : _GEN_189; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_191 = 4'h8 == index ? ram_1_8 : _GEN_190; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_192 = 4'h9 == index ? ram_1_9 : _GEN_191; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_193 = 4'ha == index ? ram_1_10 : _GEN_192; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_194 = 4'hb == index ? ram_1_11 : _GEN_193; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_195 = 4'hc == index ? ram_1_12 : _GEN_194; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_196 = 4'hd == index ? ram_1_13 : _GEN_195; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_197 = 4'he == index ? ram_1_14 : _GEN_196; // @[d_cache.scala 109:{92,92}]
  wire [127:0] _GEN_198 = 4'hf == index ? ram_1_15 : _GEN_197; // @[d_cache.scala 109:{92,92}]
  wire [190:0] _GEN_268 = {{63'd0}, _GEN_198}; // @[d_cache.scala 109:92]
  wire [190:0] _ram_1_T_4 = _GEN_268 & _ram_0_T_3; // @[d_cache.scala 109:92]
  wire [190:0] _ram_1_T_5 = _ram_0_T_1 | _ram_1_T_4; // @[d_cache.scala 109:76]
  wire [127:0] _GEN_199 = 4'h0 == index ? _ram_1_T_5[127:0] : ram_1_0; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_200 = 4'h1 == index ? _ram_1_T_5[127:0] : ram_1_1; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_201 = 4'h2 == index ? _ram_1_T_5[127:0] : ram_1_2; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_202 = 4'h3 == index ? _ram_1_T_5[127:0] : ram_1_3; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_203 = 4'h4 == index ? _ram_1_T_5[127:0] : ram_1_4; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_204 = 4'h5 == index ? _ram_1_T_5[127:0] : ram_1_5; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_205 = 4'h6 == index ? _ram_1_T_5[127:0] : ram_1_6; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_206 = 4'h7 == index ? _ram_1_T_5[127:0] : ram_1_7; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_207 = 4'h8 == index ? _ram_1_T_5[127:0] : ram_1_8; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_208 = 4'h9 == index ? _ram_1_T_5[127:0] : ram_1_9; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_209 = 4'ha == index ? _ram_1_T_5[127:0] : ram_1_10; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_210 = 4'hb == index ? _ram_1_T_5[127:0] : ram_1_11; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_211 = 4'hc == index ? _ram_1_T_5[127:0] : ram_1_12; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_212 = 4'hd == index ? _ram_1_T_5[127:0] : ram_1_13; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_213 = 4'he == index ? _ram_1_T_5[127:0] : ram_1_14; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_214 = 4'hf == index ? _ram_1_T_5[127:0] : ram_1_15; // @[d_cache.scala 109:{30,30} 20:24]
  wire [127:0] _GEN_232 = 4'h1 == index ? ram_2_1 : ram_2_0; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_233 = 4'h2 == index ? ram_2_2 : _GEN_232; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_234 = 4'h3 == index ? ram_2_3 : _GEN_233; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_235 = 4'h4 == index ? ram_2_4 : _GEN_234; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_236 = 4'h5 == index ? ram_2_5 : _GEN_235; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_237 = 4'h6 == index ? ram_2_6 : _GEN_236; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_238 = 4'h7 == index ? ram_2_7 : _GEN_237; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_239 = 4'h8 == index ? ram_2_8 : _GEN_238; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_240 = 4'h9 == index ? ram_2_9 : _GEN_239; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_241 = 4'ha == index ? ram_2_10 : _GEN_240; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_242 = 4'hb == index ? ram_2_11 : _GEN_241; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_243 = 4'hc == index ? ram_2_12 : _GEN_242; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_244 = 4'hd == index ? ram_2_13 : _GEN_243; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_245 = 4'he == index ? ram_2_14 : _GEN_244; // @[d_cache.scala 116:{92,92}]
  wire [127:0] _GEN_246 = 4'hf == index ? ram_2_15 : _GEN_245; // @[d_cache.scala 116:{92,92}]
  wire [190:0] _GEN_269 = {{63'd0}, _GEN_246}; // @[d_cache.scala 116:92]
  wire [190:0] _ram_2_T_4 = _GEN_269 & _ram_0_T_3; // @[d_cache.scala 116:92]
  wire [190:0] _ram_2_T_5 = _ram_0_T_1 | _ram_2_T_4; // @[d_cache.scala 116:76]
  wire [127:0] _GEN_247 = 4'h0 == index ? _ram_2_T_5[127:0] : ram_2_0; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_248 = 4'h1 == index ? _ram_2_T_5[127:0] : ram_2_1; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_249 = 4'h2 == index ? _ram_2_T_5[127:0] : ram_2_2; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_250 = 4'h3 == index ? _ram_2_T_5[127:0] : ram_2_3; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_251 = 4'h4 == index ? _ram_2_T_5[127:0] : ram_2_4; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_252 = 4'h5 == index ? _ram_2_T_5[127:0] : ram_2_5; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_253 = 4'h6 == index ? _ram_2_T_5[127:0] : ram_2_6; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_254 = 4'h7 == index ? _ram_2_T_5[127:0] : ram_2_7; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_255 = 4'h8 == index ? _ram_2_T_5[127:0] : ram_2_8; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_256 = 4'h9 == index ? _ram_2_T_5[127:0] : ram_2_9; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_257 = 4'ha == index ? _ram_2_T_5[127:0] : ram_2_10; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_258 = 4'hb == index ? _ram_2_T_5[127:0] : ram_2_11; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_259 = 4'hc == index ? _ram_2_T_5[127:0] : ram_2_12; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_260 = 4'hd == index ? _ram_2_T_5[127:0] : ram_2_13; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_261 = 4'he == index ? _ram_2_T_5[127:0] : ram_2_14; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_262 = 4'hf == index ? _ram_2_T_5[127:0] : ram_2_15; // @[d_cache.scala 116:{30,30} 21:24]
  wire [127:0] _GEN_280 = 4'h1 == index ? ram_3_1 : ram_3_0; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_281 = 4'h2 == index ? ram_3_2 : _GEN_280; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_282 = 4'h3 == index ? ram_3_3 : _GEN_281; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_283 = 4'h4 == index ? ram_3_4 : _GEN_282; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_284 = 4'h5 == index ? ram_3_5 : _GEN_283; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_285 = 4'h6 == index ? ram_3_6 : _GEN_284; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_286 = 4'h7 == index ? ram_3_7 : _GEN_285; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_287 = 4'h8 == index ? ram_3_8 : _GEN_286; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_288 = 4'h9 == index ? ram_3_9 : _GEN_287; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_289 = 4'ha == index ? ram_3_10 : _GEN_288; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_290 = 4'hb == index ? ram_3_11 : _GEN_289; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_291 = 4'hc == index ? ram_3_12 : _GEN_290; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_292 = 4'hd == index ? ram_3_13 : _GEN_291; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_293 = 4'he == index ? ram_3_14 : _GEN_292; // @[d_cache.scala 123:{92,92}]
  wire [127:0] _GEN_294 = 4'hf == index ? ram_3_15 : _GEN_293; // @[d_cache.scala 123:{92,92}]
  wire [190:0] _GEN_270 = {{63'd0}, _GEN_294}; // @[d_cache.scala 123:92]
  wire [190:0] _ram_3_T_4 = _GEN_270 & _ram_0_T_3; // @[d_cache.scala 123:92]
  wire [190:0] _ram_3_T_5 = _ram_0_T_1 | _ram_3_T_4; // @[d_cache.scala 123:76]
  wire [127:0] _GEN_295 = 4'h0 == index ? _ram_3_T_5[127:0] : ram_3_0; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_296 = 4'h1 == index ? _ram_3_T_5[127:0] : ram_3_1; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_297 = 4'h2 == index ? _ram_3_T_5[127:0] : ram_3_2; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_298 = 4'h3 == index ? _ram_3_T_5[127:0] : ram_3_3; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_299 = 4'h4 == index ? _ram_3_T_5[127:0] : ram_3_4; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_300 = 4'h5 == index ? _ram_3_T_5[127:0] : ram_3_5; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_301 = 4'h6 == index ? _ram_3_T_5[127:0] : ram_3_6; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_302 = 4'h7 == index ? _ram_3_T_5[127:0] : ram_3_7; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_303 = 4'h8 == index ? _ram_3_T_5[127:0] : ram_3_8; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_304 = 4'h9 == index ? _ram_3_T_5[127:0] : ram_3_9; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_305 = 4'ha == index ? _ram_3_T_5[127:0] : ram_3_10; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_306 = 4'hb == index ? _ram_3_T_5[127:0] : ram_3_11; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_307 = 4'hc == index ? _ram_3_T_5[127:0] : ram_3_12; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_308 = 4'hd == index ? _ram_3_T_5[127:0] : ram_3_13; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_309 = 4'he == index ? _ram_3_T_5[127:0] : ram_3_14; // @[d_cache.scala 123:{30,30} 22:24]
  wire [127:0] _GEN_310 = 4'hf == index ? _ram_3_T_5[127:0] : ram_3_15; // @[d_cache.scala 123:{30,30} 22:24]
  wire  _GEN_311 = _GEN_220 | dirty_3_0; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_312 = _GEN_221 | dirty_3_1; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_313 = _GEN_222 | dirty_3_2; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_314 = _GEN_223 | dirty_3_3; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_315 = _GEN_224 | dirty_3_4; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_316 = _GEN_225 | dirty_3_5; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_317 = _GEN_226 | dirty_3_6; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_318 = _GEN_227 | dirty_3_7; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_319 = _GEN_228 | dirty_3_8; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_320 = _GEN_229 | dirty_3_9; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_321 = _GEN_230 | dirty_3_10; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_322 = _GEN_263 | dirty_3_11; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_323 = _GEN_264 | dirty_3_12; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_324 = _GEN_265 | dirty_3_13; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_325 = _GEN_266 | dirty_3_14; // @[d_cache.scala 124:{32,32} 35:26]
  wire  _GEN_326 = _GEN_267 | dirty_3_15; // @[d_cache.scala 124:{32,32} 35:26]
  wire [3:0] _GEN_327 = way3_hit ? 4'h0 : 4'h4; // @[d_cache.scala 118:33 126:23]
  wire [127:0] _GEN_328 = way3_hit ? _GEN_295 : ram_3_0; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_329 = way3_hit ? _GEN_296 : ram_3_1; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_330 = way3_hit ? _GEN_297 : ram_3_2; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_331 = way3_hit ? _GEN_298 : ram_3_3; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_332 = way3_hit ? _GEN_299 : ram_3_4; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_333 = way3_hit ? _GEN_300 : ram_3_5; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_334 = way3_hit ? _GEN_301 : ram_3_6; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_335 = way3_hit ? _GEN_302 : ram_3_7; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_336 = way3_hit ? _GEN_303 : ram_3_8; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_337 = way3_hit ? _GEN_304 : ram_3_9; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_338 = way3_hit ? _GEN_305 : ram_3_10; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_339 = way3_hit ? _GEN_306 : ram_3_11; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_340 = way3_hit ? _GEN_307 : ram_3_12; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_341 = way3_hit ? _GEN_308 : ram_3_13; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_342 = way3_hit ? _GEN_309 : ram_3_14; // @[d_cache.scala 118:33 22:24]
  wire [127:0] _GEN_343 = way3_hit ? _GEN_310 : ram_3_15; // @[d_cache.scala 118:33 22:24]
  wire  _GEN_344 = way3_hit ? _GEN_311 : dirty_3_0; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_345 = way3_hit ? _GEN_312 : dirty_3_1; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_346 = way3_hit ? _GEN_313 : dirty_3_2; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_347 = way3_hit ? _GEN_314 : dirty_3_3; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_348 = way3_hit ? _GEN_315 : dirty_3_4; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_349 = way3_hit ? _GEN_316 : dirty_3_5; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_350 = way3_hit ? _GEN_317 : dirty_3_6; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_351 = way3_hit ? _GEN_318 : dirty_3_7; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_352 = way3_hit ? _GEN_319 : dirty_3_8; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_353 = way3_hit ? _GEN_320 : dirty_3_9; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_354 = way3_hit ? _GEN_321 : dirty_3_10; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_355 = way3_hit ? _GEN_322 : dirty_3_11; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_356 = way3_hit ? _GEN_323 : dirty_3_12; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_357 = way3_hit ? _GEN_324 : dirty_3_13; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_358 = way3_hit ? _GEN_325 : dirty_3_14; // @[d_cache.scala 118:33 35:26]
  wire  _GEN_359 = way3_hit ? _GEN_326 : dirty_3_15; // @[d_cache.scala 118:33 35:26]
  wire [3:0] _GEN_360 = way2_hit ? 4'h0 : _GEN_327; // @[d_cache.scala 111:34]
  wire [127:0] _GEN_361 = way2_hit ? _GEN_247 : ram_2_0; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_362 = way2_hit ? _GEN_248 : ram_2_1; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_363 = way2_hit ? _GEN_249 : ram_2_2; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_364 = way2_hit ? _GEN_250 : ram_2_3; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_365 = way2_hit ? _GEN_251 : ram_2_4; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_366 = way2_hit ? _GEN_252 : ram_2_5; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_367 = way2_hit ? _GEN_253 : ram_2_6; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_368 = way2_hit ? _GEN_254 : ram_2_7; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_369 = way2_hit ? _GEN_255 : ram_2_8; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_370 = way2_hit ? _GEN_256 : ram_2_9; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_371 = way2_hit ? _GEN_257 : ram_2_10; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_372 = way2_hit ? _GEN_258 : ram_2_11; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_373 = way2_hit ? _GEN_259 : ram_2_12; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_374 = way2_hit ? _GEN_260 : ram_2_13; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_375 = way2_hit ? _GEN_261 : ram_2_14; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_376 = way2_hit ? _GEN_262 : ram_2_15; // @[d_cache.scala 111:34 21:24]
  wire [127:0] _GEN_393 = way2_hit ? ram_3_0 : _GEN_328; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_394 = way2_hit ? ram_3_1 : _GEN_329; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_395 = way2_hit ? ram_3_2 : _GEN_330; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_396 = way2_hit ? ram_3_3 : _GEN_331; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_397 = way2_hit ? ram_3_4 : _GEN_332; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_398 = way2_hit ? ram_3_5 : _GEN_333; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_399 = way2_hit ? ram_3_6 : _GEN_334; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_400 = way2_hit ? ram_3_7 : _GEN_335; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_401 = way2_hit ? ram_3_8 : _GEN_336; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_402 = way2_hit ? ram_3_9 : _GEN_337; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_403 = way2_hit ? ram_3_10 : _GEN_338; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_404 = way2_hit ? ram_3_11 : _GEN_339; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_405 = way2_hit ? ram_3_12 : _GEN_340; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_406 = way2_hit ? ram_3_13 : _GEN_341; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_407 = way2_hit ? ram_3_14 : _GEN_342; // @[d_cache.scala 111:34 22:24]
  wire [127:0] _GEN_408 = way2_hit ? ram_3_15 : _GEN_343; // @[d_cache.scala 111:34 22:24]
  wire  _GEN_409 = way2_hit ? dirty_3_0 : _GEN_344; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_410 = way2_hit ? dirty_3_1 : _GEN_345; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_411 = way2_hit ? dirty_3_2 : _GEN_346; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_412 = way2_hit ? dirty_3_3 : _GEN_347; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_413 = way2_hit ? dirty_3_4 : _GEN_348; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_414 = way2_hit ? dirty_3_5 : _GEN_349; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_415 = way2_hit ? dirty_3_6 : _GEN_350; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_416 = way2_hit ? dirty_3_7 : _GEN_351; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_417 = way2_hit ? dirty_3_8 : _GEN_352; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_418 = way2_hit ? dirty_3_9 : _GEN_353; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_419 = way2_hit ? dirty_3_10 : _GEN_354; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_420 = way2_hit ? dirty_3_11 : _GEN_355; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_421 = way2_hit ? dirty_3_12 : _GEN_356; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_422 = way2_hit ? dirty_3_13 : _GEN_357; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_423 = way2_hit ? dirty_3_14 : _GEN_358; // @[d_cache.scala 111:34 35:26]
  wire  _GEN_424 = way2_hit ? dirty_3_15 : _GEN_359; // @[d_cache.scala 111:34 35:26]
  wire [3:0] _GEN_425 = way1_hit ? 4'h0 : _GEN_360; // @[d_cache.scala 104:33]
  wire [127:0] _GEN_426 = way1_hit ? _GEN_199 : ram_1_0; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_427 = way1_hit ? _GEN_200 : ram_1_1; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_428 = way1_hit ? _GEN_201 : ram_1_2; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_429 = way1_hit ? _GEN_202 : ram_1_3; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_430 = way1_hit ? _GEN_203 : ram_1_4; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_431 = way1_hit ? _GEN_204 : ram_1_5; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_432 = way1_hit ? _GEN_205 : ram_1_6; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_433 = way1_hit ? _GEN_206 : ram_1_7; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_434 = way1_hit ? _GEN_207 : ram_1_8; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_435 = way1_hit ? _GEN_208 : ram_1_9; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_436 = way1_hit ? _GEN_209 : ram_1_10; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_437 = way1_hit ? _GEN_210 : ram_1_11; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_438 = way1_hit ? _GEN_211 : ram_1_12; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_439 = way1_hit ? _GEN_212 : ram_1_13; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_440 = way1_hit ? _GEN_213 : ram_1_14; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_441 = way1_hit ? _GEN_214 : ram_1_15; // @[d_cache.scala 104:33 20:24]
  wire [127:0] _GEN_458 = way1_hit ? ram_2_0 : _GEN_361; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_459 = way1_hit ? ram_2_1 : _GEN_362; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_460 = way1_hit ? ram_2_2 : _GEN_363; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_461 = way1_hit ? ram_2_3 : _GEN_364; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_462 = way1_hit ? ram_2_4 : _GEN_365; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_463 = way1_hit ? ram_2_5 : _GEN_366; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_464 = way1_hit ? ram_2_6 : _GEN_367; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_465 = way1_hit ? ram_2_7 : _GEN_368; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_466 = way1_hit ? ram_2_8 : _GEN_369; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_467 = way1_hit ? ram_2_9 : _GEN_370; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_468 = way1_hit ? ram_2_10 : _GEN_371; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_469 = way1_hit ? ram_2_11 : _GEN_372; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_470 = way1_hit ? ram_2_12 : _GEN_373; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_471 = way1_hit ? ram_2_13 : _GEN_374; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_472 = way1_hit ? ram_2_14 : _GEN_375; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_473 = way1_hit ? ram_2_15 : _GEN_376; // @[d_cache.scala 104:33 21:24]
  wire [127:0] _GEN_490 = way1_hit ? ram_3_0 : _GEN_393; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_491 = way1_hit ? ram_3_1 : _GEN_394; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_492 = way1_hit ? ram_3_2 : _GEN_395; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_493 = way1_hit ? ram_3_3 : _GEN_396; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_494 = way1_hit ? ram_3_4 : _GEN_397; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_495 = way1_hit ? ram_3_5 : _GEN_398; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_496 = way1_hit ? ram_3_6 : _GEN_399; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_497 = way1_hit ? ram_3_7 : _GEN_400; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_498 = way1_hit ? ram_3_8 : _GEN_401; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_499 = way1_hit ? ram_3_9 : _GEN_402; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_500 = way1_hit ? ram_3_10 : _GEN_403; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_501 = way1_hit ? ram_3_11 : _GEN_404; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_502 = way1_hit ? ram_3_12 : _GEN_405; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_503 = way1_hit ? ram_3_13 : _GEN_406; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_504 = way1_hit ? ram_3_14 : _GEN_407; // @[d_cache.scala 104:33 22:24]
  wire [127:0] _GEN_505 = way1_hit ? ram_3_15 : _GEN_408; // @[d_cache.scala 104:33 22:24]
  wire  _GEN_506 = way1_hit ? dirty_3_0 : _GEN_409; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_507 = way1_hit ? dirty_3_1 : _GEN_410; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_508 = way1_hit ? dirty_3_2 : _GEN_411; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_509 = way1_hit ? dirty_3_3 : _GEN_412; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_510 = way1_hit ? dirty_3_4 : _GEN_413; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_511 = way1_hit ? dirty_3_5 : _GEN_414; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_512 = way1_hit ? dirty_3_6 : _GEN_415; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_513 = way1_hit ? dirty_3_7 : _GEN_416; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_514 = way1_hit ? dirty_3_8 : _GEN_417; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_515 = way1_hit ? dirty_3_9 : _GEN_418; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_516 = way1_hit ? dirty_3_10 : _GEN_419; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_517 = way1_hit ? dirty_3_11 : _GEN_420; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_518 = way1_hit ? dirty_3_12 : _GEN_421; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_519 = way1_hit ? dirty_3_13 : _GEN_422; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_520 = way1_hit ? dirty_3_14 : _GEN_423; // @[d_cache.scala 104:33 35:26]
  wire  _GEN_521 = way1_hit ? dirty_3_15 : _GEN_424; // @[d_cache.scala 104:33 35:26]
  wire [3:0] _GEN_522 = way0_hit ? 4'h0 : _GEN_425; // @[d_cache.scala 97:27]
  wire [127:0] _GEN_523 = way0_hit ? _GEN_151 : ram_0_0; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_524 = way0_hit ? _GEN_152 : ram_0_1; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_525 = way0_hit ? _GEN_153 : ram_0_2; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_526 = way0_hit ? _GEN_154 : ram_0_3; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_527 = way0_hit ? _GEN_155 : ram_0_4; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_528 = way0_hit ? _GEN_156 : ram_0_5; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_529 = way0_hit ? _GEN_157 : ram_0_6; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_530 = way0_hit ? _GEN_158 : ram_0_7; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_531 = way0_hit ? _GEN_159 : ram_0_8; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_532 = way0_hit ? _GEN_160 : ram_0_9; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_533 = way0_hit ? _GEN_161 : ram_0_10; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_534 = way0_hit ? _GEN_162 : ram_0_11; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_535 = way0_hit ? _GEN_163 : ram_0_12; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_536 = way0_hit ? _GEN_164 : ram_0_13; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_537 = way0_hit ? _GEN_165 : ram_0_14; // @[d_cache.scala 19:24 97:27]
  wire [127:0] _GEN_538 = way0_hit ? _GEN_166 : ram_0_15; // @[d_cache.scala 19:24 97:27]
  wire  _GEN_539 = way0_hit ? _GEN_167 : dirty_0_0; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_540 = way0_hit ? _GEN_168 : dirty_0_1; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_541 = way0_hit ? _GEN_169 : dirty_0_2; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_542 = way0_hit ? _GEN_170 : dirty_0_3; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_543 = way0_hit ? _GEN_171 : dirty_0_4; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_544 = way0_hit ? _GEN_172 : dirty_0_5; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_545 = way0_hit ? _GEN_173 : dirty_0_6; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_546 = way0_hit ? _GEN_174 : dirty_0_7; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_547 = way0_hit ? _GEN_175 : dirty_0_8; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_548 = way0_hit ? _GEN_176 : dirty_0_9; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_549 = way0_hit ? _GEN_177 : dirty_0_10; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_550 = way0_hit ? _GEN_178 : dirty_0_11; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_551 = way0_hit ? _GEN_179 : dirty_0_12; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_552 = way0_hit ? _GEN_180 : dirty_0_13; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_553 = way0_hit ? _GEN_181 : dirty_0_14; // @[d_cache.scala 32:26 97:27]
  wire  _GEN_554 = way0_hit ? _GEN_182 : dirty_0_15; // @[d_cache.scala 32:26 97:27]
  wire [127:0] _GEN_555 = way0_hit ? ram_1_0 : _GEN_426; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_556 = way0_hit ? ram_1_1 : _GEN_427; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_557 = way0_hit ? ram_1_2 : _GEN_428; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_558 = way0_hit ? ram_1_3 : _GEN_429; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_559 = way0_hit ? ram_1_4 : _GEN_430; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_560 = way0_hit ? ram_1_5 : _GEN_431; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_561 = way0_hit ? ram_1_6 : _GEN_432; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_562 = way0_hit ? ram_1_7 : _GEN_433; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_563 = way0_hit ? ram_1_8 : _GEN_434; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_564 = way0_hit ? ram_1_9 : _GEN_435; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_565 = way0_hit ? ram_1_10 : _GEN_436; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_566 = way0_hit ? ram_1_11 : _GEN_437; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_567 = way0_hit ? ram_1_12 : _GEN_438; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_568 = way0_hit ? ram_1_13 : _GEN_439; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_569 = way0_hit ? ram_1_14 : _GEN_440; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_570 = way0_hit ? ram_1_15 : _GEN_441; // @[d_cache.scala 20:24 97:27]
  wire [127:0] _GEN_587 = way0_hit ? ram_2_0 : _GEN_458; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_588 = way0_hit ? ram_2_1 : _GEN_459; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_589 = way0_hit ? ram_2_2 : _GEN_460; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_590 = way0_hit ? ram_2_3 : _GEN_461; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_591 = way0_hit ? ram_2_4 : _GEN_462; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_592 = way0_hit ? ram_2_5 : _GEN_463; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_593 = way0_hit ? ram_2_6 : _GEN_464; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_594 = way0_hit ? ram_2_7 : _GEN_465; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_595 = way0_hit ? ram_2_8 : _GEN_466; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_596 = way0_hit ? ram_2_9 : _GEN_467; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_597 = way0_hit ? ram_2_10 : _GEN_468; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_598 = way0_hit ? ram_2_11 : _GEN_469; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_599 = way0_hit ? ram_2_12 : _GEN_470; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_600 = way0_hit ? ram_2_13 : _GEN_471; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_601 = way0_hit ? ram_2_14 : _GEN_472; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_602 = way0_hit ? ram_2_15 : _GEN_473; // @[d_cache.scala 21:24 97:27]
  wire [127:0] _GEN_619 = way0_hit ? ram_3_0 : _GEN_490; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_620 = way0_hit ? ram_3_1 : _GEN_491; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_621 = way0_hit ? ram_3_2 : _GEN_492; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_622 = way0_hit ? ram_3_3 : _GEN_493; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_623 = way0_hit ? ram_3_4 : _GEN_494; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_624 = way0_hit ? ram_3_5 : _GEN_495; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_625 = way0_hit ? ram_3_6 : _GEN_496; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_626 = way0_hit ? ram_3_7 : _GEN_497; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_627 = way0_hit ? ram_3_8 : _GEN_498; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_628 = way0_hit ? ram_3_9 : _GEN_499; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_629 = way0_hit ? ram_3_10 : _GEN_500; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_630 = way0_hit ? ram_3_11 : _GEN_501; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_631 = way0_hit ? ram_3_12 : _GEN_502; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_632 = way0_hit ? ram_3_13 : _GEN_503; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_633 = way0_hit ? ram_3_14 : _GEN_504; // @[d_cache.scala 22:24 97:27]
  wire [127:0] _GEN_634 = way0_hit ? ram_3_15 : _GEN_505; // @[d_cache.scala 22:24 97:27]
  wire  _GEN_635 = way0_hit ? dirty_3_0 : _GEN_506; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_636 = way0_hit ? dirty_3_1 : _GEN_507; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_637 = way0_hit ? dirty_3_2 : _GEN_508; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_638 = way0_hit ? dirty_3_3 : _GEN_509; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_639 = way0_hit ? dirty_3_4 : _GEN_510; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_640 = way0_hit ? dirty_3_5 : _GEN_511; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_641 = way0_hit ? dirty_3_6 : _GEN_512; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_642 = way0_hit ? dirty_3_7 : _GEN_513; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_643 = way0_hit ? dirty_3_8 : _GEN_514; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_644 = way0_hit ? dirty_3_9 : _GEN_515; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_645 = way0_hit ? dirty_3_10 : _GEN_516; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_646 = way0_hit ? dirty_3_11 : _GEN_517; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_647 = way0_hit ? dirty_3_12 : _GEN_518; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_648 = way0_hit ? dirty_3_13 : _GEN_519; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_649 = way0_hit ? dirty_3_14 : _GEN_520; // @[d_cache.scala 35:26 97:27]
  wire  _GEN_650 = way0_hit ? dirty_3_15 : _GEN_521; // @[d_cache.scala 35:26 97:27]
  wire [63:0] _GEN_651 = ~receive_num[0] ? io_from_axi_rdata : receive_data_0; // @[d_cache.scala 131:{43,43} 47:31]
  wire [63:0] _GEN_652 = receive_num[0] ? io_from_axi_rdata : receive_data_1; // @[d_cache.scala 131:{43,43} 47:31]
  wire [2:0] _receive_num_T_1 = receive_num + 3'h1; // @[d_cache.scala 132:44]
  wire [3:0] _GEN_653 = io_from_axi_rlast ? 4'h5 : state; // @[d_cache.scala 133:40 134:27 71:24]
  wire [63:0] _GEN_654 = io_from_axi_rvalid ? _GEN_651 : receive_data_0; // @[d_cache.scala 130:37 47:31]
  wire [63:0] _GEN_655 = io_from_axi_rvalid ? _GEN_652 : receive_data_1; // @[d_cache.scala 130:37 47:31]
  wire [2:0] _GEN_656 = io_from_axi_rvalid ? _receive_num_T_1 : receive_num; // @[d_cache.scala 130:37 132:29 48:30]
  wire [3:0] _GEN_657 = io_from_axi_rvalid ? _GEN_653 : state; // @[d_cache.scala 130:37 71:24]
  wire [3:0] _GEN_658 = io_from_axi_bvalid ? 4'h0 : state; // @[d_cache.scala 139:59 140:23 71:24]
  wire [127:0] _ram_0_T_6 = {receive_data_1,receive_data_0}; // @[Cat.scala 31:58]
  wire [127:0] _GEN_659 = 4'h0 == index ? _ram_0_T_6 : ram_0_0; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_660 = 4'h1 == index ? _ram_0_T_6 : ram_0_1; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_661 = 4'h2 == index ? _ram_0_T_6 : ram_0_2; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_662 = 4'h3 == index ? _ram_0_T_6 : ram_0_3; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_663 = 4'h4 == index ? _ram_0_T_6 : ram_0_4; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_664 = 4'h5 == index ? _ram_0_T_6 : ram_0_5; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_665 = 4'h6 == index ? _ram_0_T_6 : ram_0_6; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_666 = 4'h7 == index ? _ram_0_T_6 : ram_0_7; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_667 = 4'h8 == index ? _ram_0_T_6 : ram_0_8; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_668 = 4'h9 == index ? _ram_0_T_6 : ram_0_9; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_669 = 4'ha == index ? _ram_0_T_6 : ram_0_10; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_670 = 4'hb == index ? _ram_0_T_6 : ram_0_11; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_671 = 4'hc == index ? _ram_0_T_6 : ram_0_12; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_672 = 4'hd == index ? _ram_0_T_6 : ram_0_13; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_673 = 4'he == index ? _ram_0_T_6 : ram_0_14; // @[d_cache.scala 146:{30,30} 19:24]
  wire [127:0] _GEN_674 = 4'hf == index ? _ram_0_T_6 : ram_0_15; // @[d_cache.scala 146:{30,30} 19:24]
  wire [31:0] _GEN_675 = 4'h0 == index ? _GEN_215 : tag_0_0; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_676 = 4'h1 == index ? _GEN_215 : tag_0_1; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_677 = 4'h2 == index ? _GEN_215 : tag_0_2; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_678 = 4'h3 == index ? _GEN_215 : tag_0_3; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_679 = 4'h4 == index ? _GEN_215 : tag_0_4; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_680 = 4'h5 == index ? _GEN_215 : tag_0_5; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_681 = 4'h6 == index ? _GEN_215 : tag_0_6; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_682 = 4'h7 == index ? _GEN_215 : tag_0_7; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_683 = 4'h8 == index ? _GEN_215 : tag_0_8; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_684 = 4'h9 == index ? _GEN_215 : tag_0_9; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_685 = 4'ha == index ? _GEN_215 : tag_0_10; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_686 = 4'hb == index ? _GEN_215 : tag_0_11; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_687 = 4'hc == index ? _GEN_215 : tag_0_12; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_688 = 4'hd == index ? _GEN_215 : tag_0_13; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_689 = 4'he == index ? _GEN_215 : tag_0_14; // @[d_cache.scala 147:{30,30} 24:24]
  wire [31:0] _GEN_690 = 4'hf == index ? _GEN_215 : tag_0_15; // @[d_cache.scala 147:{30,30} 24:24]
  wire  _GEN_691 = _GEN_220 | valid_0_0; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_692 = _GEN_221 | valid_0_1; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_693 = _GEN_222 | valid_0_2; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_694 = _GEN_223 | valid_0_3; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_695 = _GEN_224 | valid_0_4; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_696 = _GEN_225 | valid_0_5; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_697 = _GEN_226 | valid_0_6; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_698 = _GEN_227 | valid_0_7; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_699 = _GEN_228 | valid_0_8; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_700 = _GEN_229 | valid_0_9; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_701 = _GEN_230 | valid_0_10; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_702 = _GEN_263 | valid_0_11; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_703 = _GEN_264 | valid_0_12; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_704 = _GEN_265 | valid_0_13; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_705 = _GEN_266 | valid_0_14; // @[d_cache.scala 148:{32,32} 28:26]
  wire  _GEN_706 = _GEN_267 | valid_0_15; // @[d_cache.scala 148:{32,32} 28:26]
  wire [7:0] _GEN_708 = 4'h1 == index ? quene_1 : quene_0; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_709 = 4'h2 == index ? quene_2 : _GEN_708; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_710 = 4'h3 == index ? quene_3 : _GEN_709; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_711 = 4'h4 == index ? quene_4 : _GEN_710; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_712 = 4'h5 == index ? quene_5 : _GEN_711; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_713 = 4'h6 == index ? quene_6 : _GEN_712; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_714 = 4'h7 == index ? quene_7 : _GEN_713; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_715 = 4'h8 == index ? quene_8 : _GEN_714; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_716 = 4'h9 == index ? quene_9 : _GEN_715; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_717 = 4'ha == index ? quene_10 : _GEN_716; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_718 = 4'hb == index ? quene_11 : _GEN_717; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_719 = 4'hc == index ? quene_12 : _GEN_718; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_720 = 4'hd == index ? quene_13 : _GEN_719; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_721 = 4'he == index ? quene_14 : _GEN_720; // @[d_cache.scala 149:{46,46}]
  wire [7:0] _GEN_722 = 4'hf == index ? quene_15 : _GEN_721; // @[d_cache.scala 149:{46,46}]
  wire [9:0] _GEN_450 = {_GEN_722, 2'h0}; // @[d_cache.scala 149:46]
  wire [10:0] _quene_T = {{1'd0}, _GEN_450}; // @[d_cache.scala 149:46]
  wire [7:0] _GEN_723 = 4'h0 == index ? _quene_T[7:0] : quene_0; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_724 = 4'h1 == index ? _quene_T[7:0] : quene_1; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_725 = 4'h2 == index ? _quene_T[7:0] : quene_2; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_726 = 4'h3 == index ? _quene_T[7:0] : quene_3; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_727 = 4'h4 == index ? _quene_T[7:0] : quene_4; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_728 = 4'h5 == index ? _quene_T[7:0] : quene_5; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_729 = 4'h6 == index ? _quene_T[7:0] : quene_6; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_730 = 4'h7 == index ? _quene_T[7:0] : quene_7; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_731 = 4'h8 == index ? _quene_T[7:0] : quene_8; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_732 = 4'h9 == index ? _quene_T[7:0] : quene_9; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_733 = 4'ha == index ? _quene_T[7:0] : quene_10; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_734 = 4'hb == index ? _quene_T[7:0] : quene_11; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_735 = 4'hc == index ? _quene_T[7:0] : quene_12; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_736 = 4'hd == index ? _quene_T[7:0] : quene_13; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_737 = 4'he == index ? _quene_T[7:0] : quene_14; // @[d_cache.scala 149:{30,30} 49:24]
  wire [7:0] _GEN_738 = 4'hf == index ? _quene_T[7:0] : quene_15; // @[d_cache.scala 149:{30,30} 49:24]
  wire [127:0] _GEN_739 = 4'h0 == index ? _ram_0_T_6 : ram_1_0; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_740 = 4'h1 == index ? _ram_0_T_6 : ram_1_1; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_741 = 4'h2 == index ? _ram_0_T_6 : ram_1_2; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_742 = 4'h3 == index ? _ram_0_T_6 : ram_1_3; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_743 = 4'h4 == index ? _ram_0_T_6 : ram_1_4; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_744 = 4'h5 == index ? _ram_0_T_6 : ram_1_5; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_745 = 4'h6 == index ? _ram_0_T_6 : ram_1_6; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_746 = 4'h7 == index ? _ram_0_T_6 : ram_1_7; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_747 = 4'h8 == index ? _ram_0_T_6 : ram_1_8; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_748 = 4'h9 == index ? _ram_0_T_6 : ram_1_9; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_749 = 4'ha == index ? _ram_0_T_6 : ram_1_10; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_750 = 4'hb == index ? _ram_0_T_6 : ram_1_11; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_751 = 4'hc == index ? _ram_0_T_6 : ram_1_12; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_752 = 4'hd == index ? _ram_0_T_6 : ram_1_13; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_753 = 4'he == index ? _ram_0_T_6 : ram_1_14; // @[d_cache.scala 152:{30,30} 20:24]
  wire [127:0] _GEN_754 = 4'hf == index ? _ram_0_T_6 : ram_1_15; // @[d_cache.scala 152:{30,30} 20:24]
  wire [31:0] _GEN_755 = 4'h0 == index ? _GEN_215 : tag_1_0; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_756 = 4'h1 == index ? _GEN_215 : tag_1_1; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_757 = 4'h2 == index ? _GEN_215 : tag_1_2; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_758 = 4'h3 == index ? _GEN_215 : tag_1_3; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_759 = 4'h4 == index ? _GEN_215 : tag_1_4; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_760 = 4'h5 == index ? _GEN_215 : tag_1_5; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_761 = 4'h6 == index ? _GEN_215 : tag_1_6; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_762 = 4'h7 == index ? _GEN_215 : tag_1_7; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_763 = 4'h8 == index ? _GEN_215 : tag_1_8; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_764 = 4'h9 == index ? _GEN_215 : tag_1_9; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_765 = 4'ha == index ? _GEN_215 : tag_1_10; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_766 = 4'hb == index ? _GEN_215 : tag_1_11; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_767 = 4'hc == index ? _GEN_215 : tag_1_12; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_768 = 4'hd == index ? _GEN_215 : tag_1_13; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_769 = 4'he == index ? _GEN_215 : tag_1_14; // @[d_cache.scala 153:{30,30} 25:24]
  wire [31:0] _GEN_770 = 4'hf == index ? _GEN_215 : tag_1_15; // @[d_cache.scala 153:{30,30} 25:24]
  wire  _GEN_771 = _GEN_220 | valid_1_0; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_772 = _GEN_221 | valid_1_1; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_773 = _GEN_222 | valid_1_2; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_774 = _GEN_223 | valid_1_3; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_775 = _GEN_224 | valid_1_4; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_776 = _GEN_225 | valid_1_5; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_777 = _GEN_226 | valid_1_6; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_778 = _GEN_227 | valid_1_7; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_779 = _GEN_228 | valid_1_8; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_780 = _GEN_229 | valid_1_9; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_781 = _GEN_230 | valid_1_10; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_782 = _GEN_263 | valid_1_11; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_783 = _GEN_264 | valid_1_12; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_784 = _GEN_265 | valid_1_13; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_785 = _GEN_266 | valid_1_14; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_786 = _GEN_267 | valid_1_15; // @[d_cache.scala 154:{32,32} 29:26]
  wire [10:0] _quene_T_2 = _quene_T | 11'h1; // @[d_cache.scala 155:55]
  wire [7:0] _GEN_787 = 4'h0 == index ? _quene_T_2[7:0] : quene_0; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_788 = 4'h1 == index ? _quene_T_2[7:0] : quene_1; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_789 = 4'h2 == index ? _quene_T_2[7:0] : quene_2; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_790 = 4'h3 == index ? _quene_T_2[7:0] : quene_3; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_791 = 4'h4 == index ? _quene_T_2[7:0] : quene_4; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_792 = 4'h5 == index ? _quene_T_2[7:0] : quene_5; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_793 = 4'h6 == index ? _quene_T_2[7:0] : quene_6; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_794 = 4'h7 == index ? _quene_T_2[7:0] : quene_7; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_795 = 4'h8 == index ? _quene_T_2[7:0] : quene_8; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_796 = 4'h9 == index ? _quene_T_2[7:0] : quene_9; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_797 = 4'ha == index ? _quene_T_2[7:0] : quene_10; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_798 = 4'hb == index ? _quene_T_2[7:0] : quene_11; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_799 = 4'hc == index ? _quene_T_2[7:0] : quene_12; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_800 = 4'hd == index ? _quene_T_2[7:0] : quene_13; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_801 = 4'he == index ? _quene_T_2[7:0] : quene_14; // @[d_cache.scala 155:{30,30} 49:24]
  wire [7:0] _GEN_802 = 4'hf == index ? _quene_T_2[7:0] : quene_15; // @[d_cache.scala 155:{30,30} 49:24]
  wire [127:0] _GEN_803 = 4'h0 == index ? _ram_0_T_6 : ram_2_0; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_804 = 4'h1 == index ? _ram_0_T_6 : ram_2_1; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_805 = 4'h2 == index ? _ram_0_T_6 : ram_2_2; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_806 = 4'h3 == index ? _ram_0_T_6 : ram_2_3; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_807 = 4'h4 == index ? _ram_0_T_6 : ram_2_4; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_808 = 4'h5 == index ? _ram_0_T_6 : ram_2_5; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_809 = 4'h6 == index ? _ram_0_T_6 : ram_2_6; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_810 = 4'h7 == index ? _ram_0_T_6 : ram_2_7; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_811 = 4'h8 == index ? _ram_0_T_6 : ram_2_8; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_812 = 4'h9 == index ? _ram_0_T_6 : ram_2_9; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_813 = 4'ha == index ? _ram_0_T_6 : ram_2_10; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_814 = 4'hb == index ? _ram_0_T_6 : ram_2_11; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_815 = 4'hc == index ? _ram_0_T_6 : ram_2_12; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_816 = 4'hd == index ? _ram_0_T_6 : ram_2_13; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_817 = 4'he == index ? _ram_0_T_6 : ram_2_14; // @[d_cache.scala 158:{30,30} 21:24]
  wire [127:0] _GEN_818 = 4'hf == index ? _ram_0_T_6 : ram_2_15; // @[d_cache.scala 158:{30,30} 21:24]
  wire [31:0] _GEN_819 = 4'h0 == index ? _GEN_215 : tag_2_0; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_820 = 4'h1 == index ? _GEN_215 : tag_2_1; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_821 = 4'h2 == index ? _GEN_215 : tag_2_2; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_822 = 4'h3 == index ? _GEN_215 : tag_2_3; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_823 = 4'h4 == index ? _GEN_215 : tag_2_4; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_824 = 4'h5 == index ? _GEN_215 : tag_2_5; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_825 = 4'h6 == index ? _GEN_215 : tag_2_6; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_826 = 4'h7 == index ? _GEN_215 : tag_2_7; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_827 = 4'h8 == index ? _GEN_215 : tag_2_8; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_828 = 4'h9 == index ? _GEN_215 : tag_2_9; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_829 = 4'ha == index ? _GEN_215 : tag_2_10; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_830 = 4'hb == index ? _GEN_215 : tag_2_11; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_831 = 4'hc == index ? _GEN_215 : tag_2_12; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_832 = 4'hd == index ? _GEN_215 : tag_2_13; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_833 = 4'he == index ? _GEN_215 : tag_2_14; // @[d_cache.scala 159:{30,30} 26:24]
  wire [31:0] _GEN_834 = 4'hf == index ? _GEN_215 : tag_2_15; // @[d_cache.scala 159:{30,30} 26:24]
  wire  _GEN_835 = _GEN_220 | valid_2_0; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_836 = _GEN_221 | valid_2_1; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_837 = _GEN_222 | valid_2_2; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_838 = _GEN_223 | valid_2_3; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_839 = _GEN_224 | valid_2_4; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_840 = _GEN_225 | valid_2_5; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_841 = _GEN_226 | valid_2_6; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_842 = _GEN_227 | valid_2_7; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_843 = _GEN_228 | valid_2_8; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_844 = _GEN_229 | valid_2_9; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_845 = _GEN_230 | valid_2_10; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_846 = _GEN_263 | valid_2_11; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_847 = _GEN_264 | valid_2_12; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_848 = _GEN_265 | valid_2_13; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_849 = _GEN_266 | valid_2_14; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_850 = _GEN_267 | valid_2_15; // @[d_cache.scala 160:{32,32} 30:26]
  wire [10:0] _quene_T_4 = _quene_T | 11'h2; // @[d_cache.scala 161:55]
  wire [7:0] _GEN_851 = 4'h0 == index ? _quene_T_4[7:0] : quene_0; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_852 = 4'h1 == index ? _quene_T_4[7:0] : quene_1; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_853 = 4'h2 == index ? _quene_T_4[7:0] : quene_2; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_854 = 4'h3 == index ? _quene_T_4[7:0] : quene_3; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_855 = 4'h4 == index ? _quene_T_4[7:0] : quene_4; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_856 = 4'h5 == index ? _quene_T_4[7:0] : quene_5; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_857 = 4'h6 == index ? _quene_T_4[7:0] : quene_6; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_858 = 4'h7 == index ? _quene_T_4[7:0] : quene_7; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_859 = 4'h8 == index ? _quene_T_4[7:0] : quene_8; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_860 = 4'h9 == index ? _quene_T_4[7:0] : quene_9; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_861 = 4'ha == index ? _quene_T_4[7:0] : quene_10; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_862 = 4'hb == index ? _quene_T_4[7:0] : quene_11; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_863 = 4'hc == index ? _quene_T_4[7:0] : quene_12; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_864 = 4'hd == index ? _quene_T_4[7:0] : quene_13; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_865 = 4'he == index ? _quene_T_4[7:0] : quene_14; // @[d_cache.scala 161:{30,30} 49:24]
  wire [7:0] _GEN_866 = 4'hf == index ? _quene_T_4[7:0] : quene_15; // @[d_cache.scala 161:{30,30} 49:24]
  wire [127:0] _GEN_867 = 4'h0 == index ? _ram_0_T_6 : ram_3_0; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_868 = 4'h1 == index ? _ram_0_T_6 : ram_3_1; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_869 = 4'h2 == index ? _ram_0_T_6 : ram_3_2; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_870 = 4'h3 == index ? _ram_0_T_6 : ram_3_3; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_871 = 4'h4 == index ? _ram_0_T_6 : ram_3_4; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_872 = 4'h5 == index ? _ram_0_T_6 : ram_3_5; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_873 = 4'h6 == index ? _ram_0_T_6 : ram_3_6; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_874 = 4'h7 == index ? _ram_0_T_6 : ram_3_7; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_875 = 4'h8 == index ? _ram_0_T_6 : ram_3_8; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_876 = 4'h9 == index ? _ram_0_T_6 : ram_3_9; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_877 = 4'ha == index ? _ram_0_T_6 : ram_3_10; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_878 = 4'hb == index ? _ram_0_T_6 : ram_3_11; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_879 = 4'hc == index ? _ram_0_T_6 : ram_3_12; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_880 = 4'hd == index ? _ram_0_T_6 : ram_3_13; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_881 = 4'he == index ? _ram_0_T_6 : ram_3_14; // @[d_cache.scala 164:{30,30} 22:24]
  wire [127:0] _GEN_882 = 4'hf == index ? _ram_0_T_6 : ram_3_15; // @[d_cache.scala 164:{30,30} 22:24]
  wire [31:0] _GEN_883 = 4'h0 == index ? _GEN_215 : tag_3_0; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_884 = 4'h1 == index ? _GEN_215 : tag_3_1; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_885 = 4'h2 == index ? _GEN_215 : tag_3_2; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_886 = 4'h3 == index ? _GEN_215 : tag_3_3; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_887 = 4'h4 == index ? _GEN_215 : tag_3_4; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_888 = 4'h5 == index ? _GEN_215 : tag_3_5; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_889 = 4'h6 == index ? _GEN_215 : tag_3_6; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_890 = 4'h7 == index ? _GEN_215 : tag_3_7; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_891 = 4'h8 == index ? _GEN_215 : tag_3_8; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_892 = 4'h9 == index ? _GEN_215 : tag_3_9; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_893 = 4'ha == index ? _GEN_215 : tag_3_10; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_894 = 4'hb == index ? _GEN_215 : tag_3_11; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_895 = 4'hc == index ? _GEN_215 : tag_3_12; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_896 = 4'hd == index ? _GEN_215 : tag_3_13; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_897 = 4'he == index ? _GEN_215 : tag_3_14; // @[d_cache.scala 165:{30,30} 27:24]
  wire [31:0] _GEN_898 = 4'hf == index ? _GEN_215 : tag_3_15; // @[d_cache.scala 165:{30,30} 27:24]
  wire  _GEN_899 = _GEN_220 | valid_3_0; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_900 = _GEN_221 | valid_3_1; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_901 = _GEN_222 | valid_3_2; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_902 = _GEN_223 | valid_3_3; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_903 = _GEN_224 | valid_3_4; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_904 = _GEN_225 | valid_3_5; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_905 = _GEN_226 | valid_3_6; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_906 = _GEN_227 | valid_3_7; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_907 = _GEN_228 | valid_3_8; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_908 = _GEN_229 | valid_3_9; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_909 = _GEN_230 | valid_3_10; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_910 = _GEN_263 | valid_3_11; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_911 = _GEN_264 | valid_3_12; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_912 = _GEN_265 | valid_3_13; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_913 = _GEN_266 | valid_3_14; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_914 = _GEN_267 | valid_3_15; // @[d_cache.scala 166:{32,32} 31:26]
  wire [10:0] _quene_T_6 = _quene_T | 11'h3; // @[d_cache.scala 167:55]
  wire [7:0] _GEN_915 = 4'h0 == index ? _quene_T_6[7:0] : quene_0; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_916 = 4'h1 == index ? _quene_T_6[7:0] : quene_1; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_917 = 4'h2 == index ? _quene_T_6[7:0] : quene_2; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_918 = 4'h3 == index ? _quene_T_6[7:0] : quene_3; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_919 = 4'h4 == index ? _quene_T_6[7:0] : quene_4; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_920 = 4'h5 == index ? _quene_T_6[7:0] : quene_5; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_921 = 4'h6 == index ? _quene_T_6[7:0] : quene_6; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_922 = 4'h7 == index ? _quene_T_6[7:0] : quene_7; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_923 = 4'h8 == index ? _quene_T_6[7:0] : quene_8; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_924 = 4'h9 == index ? _quene_T_6[7:0] : quene_9; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_925 = 4'ha == index ? _quene_T_6[7:0] : quene_10; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_926 = 4'hb == index ? _quene_T_6[7:0] : quene_11; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_927 = 4'hc == index ? _quene_T_6[7:0] : quene_12; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_928 = 4'hd == index ? _quene_T_6[7:0] : quene_13; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_929 = 4'he == index ? _quene_T_6[7:0] : quene_14; // @[d_cache.scala 167:{30,30} 49:24]
  wire [7:0] _GEN_930 = 4'hf == index ? _quene_T_6[7:0] : quene_15; // @[d_cache.scala 167:{30,30} 49:24]
  wire  _GEN_932 = 4'h1 == index ? dirty_0_1 : dirty_0_0; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_933 = 4'h2 == index ? dirty_0_2 : _GEN_932; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_934 = 4'h3 == index ? dirty_0_3 : _GEN_933; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_935 = 4'h4 == index ? dirty_0_4 : _GEN_934; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_936 = 4'h5 == index ? dirty_0_5 : _GEN_935; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_937 = 4'h6 == index ? dirty_0_6 : _GEN_936; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_938 = 4'h7 == index ? dirty_0_7 : _GEN_937; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_939 = 4'h8 == index ? dirty_0_8 : _GEN_938; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_940 = 4'h9 == index ? dirty_0_9 : _GEN_939; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_941 = 4'ha == index ? dirty_0_10 : _GEN_940; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_942 = 4'hb == index ? dirty_0_11 : _GEN_941; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_943 = 4'hc == index ? dirty_0_12 : _GEN_942; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_944 = 4'hd == index ? dirty_0_13 : _GEN_943; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_945 = 4'he == index ? dirty_0_14 : _GEN_944; // @[d_cache.scala 171:{40,40}]
  wire  _GEN_946 = 4'hf == index ? dirty_0_15 : _GEN_945; // @[d_cache.scala 171:{40,40}]
  wire [39:0] _write_back_addr_T_1 = {_GEN_15,index,4'h0}; // @[Cat.scala 31:58]
  wire  _GEN_947 = 4'h0 == index ? 1'h0 : dirty_0_0; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_948 = 4'h1 == index ? 1'h0 : dirty_0_1; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_949 = 4'h2 == index ? 1'h0 : dirty_0_2; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_950 = 4'h3 == index ? 1'h0 : dirty_0_3; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_951 = 4'h4 == index ? 1'h0 : dirty_0_4; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_952 = 4'h5 == index ? 1'h0 : dirty_0_5; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_953 = 4'h6 == index ? 1'h0 : dirty_0_6; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_954 = 4'h7 == index ? 1'h0 : dirty_0_7; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_955 = 4'h8 == index ? 1'h0 : dirty_0_8; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_956 = 4'h9 == index ? 1'h0 : dirty_0_9; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_957 = 4'ha == index ? 1'h0 : dirty_0_10; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_958 = 4'hb == index ? 1'h0 : dirty_0_11; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_959 = 4'hc == index ? 1'h0 : dirty_0_12; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_960 = 4'hd == index ? 1'h0 : dirty_0_13; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_961 = 4'he == index ? 1'h0 : dirty_0_14; // @[d_cache.scala 174:{40,40} 32:26]
  wire  _GEN_962 = 4'hf == index ? 1'h0 : dirty_0_15; // @[d_cache.scala 174:{40,40} 32:26]
  wire [127:0] _GEN_963 = _GEN_946 ? _GEN_150 : write_back_data; // @[d_cache.scala 171:47 172:41 41:34]
  wire [39:0] _GEN_964 = _GEN_946 ? _write_back_addr_T_1 : {{8'd0}, write_back_addr}; // @[d_cache.scala 171:47 173:41 42:34]
  wire  _GEN_965 = _GEN_946 ? _GEN_947 : dirty_0_0; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_966 = _GEN_946 ? _GEN_948 : dirty_0_1; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_967 = _GEN_946 ? _GEN_949 : dirty_0_2; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_968 = _GEN_946 ? _GEN_950 : dirty_0_3; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_969 = _GEN_946 ? _GEN_951 : dirty_0_4; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_970 = _GEN_946 ? _GEN_952 : dirty_0_5; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_971 = _GEN_946 ? _GEN_953 : dirty_0_6; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_972 = _GEN_946 ? _GEN_954 : dirty_0_7; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_973 = _GEN_946 ? _GEN_955 : dirty_0_8; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_974 = _GEN_946 ? _GEN_956 : dirty_0_9; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_975 = _GEN_946 ? _GEN_957 : dirty_0_10; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_976 = _GEN_946 ? _GEN_958 : dirty_0_11; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_977 = _GEN_946 ? _GEN_959 : dirty_0_12; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_978 = _GEN_946 ? _GEN_960 : dirty_0_13; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_979 = _GEN_946 ? _GEN_961 : dirty_0_14; // @[d_cache.scala 171:47 32:26]
  wire  _GEN_980 = _GEN_946 ? _GEN_962 : dirty_0_15; // @[d_cache.scala 171:47 32:26]
  wire [3:0] _GEN_981 = _GEN_946 ? 4'h6 : 4'h1; // @[d_cache.scala 171:47 175:31 177:31]
  wire [39:0] _write_back_addr_T_3 = {_GEN_47,index,4'h0}; // @[Cat.scala 31:58]
  wire [127:0] _GEN_1062 = _GEN_946 ? _GEN_198 : write_back_data; // @[d_cache.scala 184:47 185:41 41:34]
  wire [39:0] _GEN_1063 = _GEN_946 ? _write_back_addr_T_3 : {{8'd0}, write_back_addr}; // @[d_cache.scala 184:47 186:41 42:34]
  wire [39:0] _write_back_addr_T_5 = {_GEN_79,index,4'h0}; // @[Cat.scala 31:58]
  wire [127:0] _GEN_1161 = _GEN_946 ? _GEN_246 : write_back_data; // @[d_cache.scala 197:47 198:41 41:34]
  wire [39:0] _GEN_1162 = _GEN_946 ? _write_back_addr_T_5 : {{8'd0}, write_back_addr}; // @[d_cache.scala 197:47 199:41 42:34]
  wire  _GEN_1245 = 4'h1 == index ? dirty_3_1 : dirty_3_0; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1246 = 4'h2 == index ? dirty_3_2 : _GEN_1245; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1247 = 4'h3 == index ? dirty_3_3 : _GEN_1246; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1248 = 4'h4 == index ? dirty_3_4 : _GEN_1247; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1249 = 4'h5 == index ? dirty_3_5 : _GEN_1248; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1250 = 4'h6 == index ? dirty_3_6 : _GEN_1249; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1251 = 4'h7 == index ? dirty_3_7 : _GEN_1250; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1252 = 4'h8 == index ? dirty_3_8 : _GEN_1251; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1253 = 4'h9 == index ? dirty_3_9 : _GEN_1252; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1254 = 4'ha == index ? dirty_3_10 : _GEN_1253; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1255 = 4'hb == index ? dirty_3_11 : _GEN_1254; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1256 = 4'hc == index ? dirty_3_12 : _GEN_1255; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1257 = 4'hd == index ? dirty_3_13 : _GEN_1256; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1258 = 4'he == index ? dirty_3_14 : _GEN_1257; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1259 = 4'hf == index ? dirty_3_15 : _GEN_1258; // @[d_cache.scala 210:{40,40}]
  wire [39:0] _write_back_addr_T_7 = {_GEN_111,index,4'h0}; // @[Cat.scala 31:58]
  wire  _GEN_1260 = 4'h0 == index ? 1'h0 : dirty_3_0; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1261 = 4'h1 == index ? 1'h0 : dirty_3_1; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1262 = 4'h2 == index ? 1'h0 : dirty_3_2; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1263 = 4'h3 == index ? 1'h0 : dirty_3_3; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1264 = 4'h4 == index ? 1'h0 : dirty_3_4; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1265 = 4'h5 == index ? 1'h0 : dirty_3_5; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1266 = 4'h6 == index ? 1'h0 : dirty_3_6; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1267 = 4'h7 == index ? 1'h0 : dirty_3_7; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1268 = 4'h8 == index ? 1'h0 : dirty_3_8; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1269 = 4'h9 == index ? 1'h0 : dirty_3_9; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1270 = 4'ha == index ? 1'h0 : dirty_3_10; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1271 = 4'hb == index ? 1'h0 : dirty_3_11; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1272 = 4'hc == index ? 1'h0 : dirty_3_12; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1273 = 4'hd == index ? 1'h0 : dirty_3_13; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1274 = 4'he == index ? 1'h0 : dirty_3_14; // @[d_cache.scala 213:{40,40} 35:26]
  wire  _GEN_1275 = 4'hf == index ? 1'h0 : dirty_3_15; // @[d_cache.scala 213:{40,40} 35:26]
  wire [127:0] _GEN_1276 = _GEN_1259 ? _GEN_294 : write_back_data; // @[d_cache.scala 210:47 211:41 41:34]
  wire [39:0] _GEN_1277 = _GEN_1259 ? _write_back_addr_T_7 : {{8'd0}, write_back_addr}; // @[d_cache.scala 210:47 212:41 42:34]
  wire  _GEN_1278 = _GEN_1259 ? _GEN_1260 : dirty_3_0; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1279 = _GEN_1259 ? _GEN_1261 : dirty_3_1; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1280 = _GEN_1259 ? _GEN_1262 : dirty_3_2; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1281 = _GEN_1259 ? _GEN_1263 : dirty_3_3; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1282 = _GEN_1259 ? _GEN_1264 : dirty_3_4; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1283 = _GEN_1259 ? _GEN_1265 : dirty_3_5; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1284 = _GEN_1259 ? _GEN_1266 : dirty_3_6; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1285 = _GEN_1259 ? _GEN_1267 : dirty_3_7; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1286 = _GEN_1259 ? _GEN_1268 : dirty_3_8; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1287 = _GEN_1259 ? _GEN_1269 : dirty_3_9; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1288 = _GEN_1259 ? _GEN_1270 : dirty_3_10; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1289 = _GEN_1259 ? _GEN_1271 : dirty_3_11; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1290 = _GEN_1259 ? _GEN_1272 : dirty_3_12; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1291 = _GEN_1259 ? _GEN_1273 : dirty_3_13; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1292 = _GEN_1259 ? _GEN_1274 : dirty_3_14; // @[d_cache.scala 210:47 35:26]
  wire  _GEN_1293 = _GEN_1259 ? _GEN_1275 : dirty_3_15; // @[d_cache.scala 210:47 35:26]
  wire [3:0] _GEN_1294 = _GEN_1259 ? 4'h6 : 4'h1; // @[d_cache.scala 210:47 214:31 216:31]
  wire [127:0] _GEN_1359 = _GEN_722[7:6] == 2'h2 ? _GEN_1161 : _GEN_1276; // @[d_cache.scala 196:52]
  wire [39:0] _GEN_1360 = _GEN_722[7:6] == 2'h2 ? _GEN_1162 : _GEN_1277; // @[d_cache.scala 196:52]
  wire [3:0] _GEN_1377 = _GEN_722[7:6] == 2'h2 ? _GEN_981 : _GEN_1294; // @[d_cache.scala 196:52]
  wire [127:0] _GEN_1378 = _GEN_722[7:6] == 2'h2 ? _GEN_803 : ram_2_0; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1379 = _GEN_722[7:6] == 2'h2 ? _GEN_804 : ram_2_1; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1380 = _GEN_722[7:6] == 2'h2 ? _GEN_805 : ram_2_2; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1381 = _GEN_722[7:6] == 2'h2 ? _GEN_806 : ram_2_3; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1382 = _GEN_722[7:6] == 2'h2 ? _GEN_807 : ram_2_4; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1383 = _GEN_722[7:6] == 2'h2 ? _GEN_808 : ram_2_5; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1384 = _GEN_722[7:6] == 2'h2 ? _GEN_809 : ram_2_6; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1385 = _GEN_722[7:6] == 2'h2 ? _GEN_810 : ram_2_7; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1386 = _GEN_722[7:6] == 2'h2 ? _GEN_811 : ram_2_8; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1387 = _GEN_722[7:6] == 2'h2 ? _GEN_812 : ram_2_9; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1388 = _GEN_722[7:6] == 2'h2 ? _GEN_813 : ram_2_10; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1389 = _GEN_722[7:6] == 2'h2 ? _GEN_814 : ram_2_11; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1390 = _GEN_722[7:6] == 2'h2 ? _GEN_815 : ram_2_12; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1391 = _GEN_722[7:6] == 2'h2 ? _GEN_816 : ram_2_13; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1392 = _GEN_722[7:6] == 2'h2 ? _GEN_817 : ram_2_14; // @[d_cache.scala 196:52 21:24]
  wire [127:0] _GEN_1393 = _GEN_722[7:6] == 2'h2 ? _GEN_818 : ram_2_15; // @[d_cache.scala 196:52 21:24]
  wire [31:0] _GEN_1394 = _GEN_722[7:6] == 2'h2 ? _GEN_819 : tag_2_0; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1395 = _GEN_722[7:6] == 2'h2 ? _GEN_820 : tag_2_1; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1396 = _GEN_722[7:6] == 2'h2 ? _GEN_821 : tag_2_2; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1397 = _GEN_722[7:6] == 2'h2 ? _GEN_822 : tag_2_3; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1398 = _GEN_722[7:6] == 2'h2 ? _GEN_823 : tag_2_4; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1399 = _GEN_722[7:6] == 2'h2 ? _GEN_824 : tag_2_5; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1400 = _GEN_722[7:6] == 2'h2 ? _GEN_825 : tag_2_6; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1401 = _GEN_722[7:6] == 2'h2 ? _GEN_826 : tag_2_7; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1402 = _GEN_722[7:6] == 2'h2 ? _GEN_827 : tag_2_8; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1403 = _GEN_722[7:6] == 2'h2 ? _GEN_828 : tag_2_9; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1404 = _GEN_722[7:6] == 2'h2 ? _GEN_829 : tag_2_10; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1405 = _GEN_722[7:6] == 2'h2 ? _GEN_830 : tag_2_11; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1406 = _GEN_722[7:6] == 2'h2 ? _GEN_831 : tag_2_12; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1407 = _GEN_722[7:6] == 2'h2 ? _GEN_832 : tag_2_13; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1408 = _GEN_722[7:6] == 2'h2 ? _GEN_833 : tag_2_14; // @[d_cache.scala 196:52 26:24]
  wire [31:0] _GEN_1409 = _GEN_722[7:6] == 2'h2 ? _GEN_834 : tag_2_15; // @[d_cache.scala 196:52 26:24]
  wire  _GEN_1410 = _GEN_722[7:6] == 2'h2 ? _GEN_835 : valid_2_0; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1411 = _GEN_722[7:6] == 2'h2 ? _GEN_836 : valid_2_1; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1412 = _GEN_722[7:6] == 2'h2 ? _GEN_837 : valid_2_2; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1413 = _GEN_722[7:6] == 2'h2 ? _GEN_838 : valid_2_3; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1414 = _GEN_722[7:6] == 2'h2 ? _GEN_839 : valid_2_4; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1415 = _GEN_722[7:6] == 2'h2 ? _GEN_840 : valid_2_5; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1416 = _GEN_722[7:6] == 2'h2 ? _GEN_841 : valid_2_6; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1417 = _GEN_722[7:6] == 2'h2 ? _GEN_842 : valid_2_7; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1418 = _GEN_722[7:6] == 2'h2 ? _GEN_843 : valid_2_8; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1419 = _GEN_722[7:6] == 2'h2 ? _GEN_844 : valid_2_9; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1420 = _GEN_722[7:6] == 2'h2 ? _GEN_845 : valid_2_10; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1421 = _GEN_722[7:6] == 2'h2 ? _GEN_846 : valid_2_11; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1422 = _GEN_722[7:6] == 2'h2 ? _GEN_847 : valid_2_12; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1423 = _GEN_722[7:6] == 2'h2 ? _GEN_848 : valid_2_13; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1424 = _GEN_722[7:6] == 2'h2 ? _GEN_849 : valid_2_14; // @[d_cache.scala 196:52 30:26]
  wire  _GEN_1425 = _GEN_722[7:6] == 2'h2 ? _GEN_850 : valid_2_15; // @[d_cache.scala 196:52 30:26]
  wire [7:0] _GEN_1426 = _GEN_722[7:6] == 2'h2 ? _GEN_851 : _GEN_915; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1427 = _GEN_722[7:6] == 2'h2 ? _GEN_852 : _GEN_916; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1428 = _GEN_722[7:6] == 2'h2 ? _GEN_853 : _GEN_917; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1429 = _GEN_722[7:6] == 2'h2 ? _GEN_854 : _GEN_918; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1430 = _GEN_722[7:6] == 2'h2 ? _GEN_855 : _GEN_919; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1431 = _GEN_722[7:6] == 2'h2 ? _GEN_856 : _GEN_920; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1432 = _GEN_722[7:6] == 2'h2 ? _GEN_857 : _GEN_921; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1433 = _GEN_722[7:6] == 2'h2 ? _GEN_858 : _GEN_922; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1434 = _GEN_722[7:6] == 2'h2 ? _GEN_859 : _GEN_923; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1435 = _GEN_722[7:6] == 2'h2 ? _GEN_860 : _GEN_924; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1436 = _GEN_722[7:6] == 2'h2 ? _GEN_861 : _GEN_925; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1437 = _GEN_722[7:6] == 2'h2 ? _GEN_862 : _GEN_926; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1438 = _GEN_722[7:6] == 2'h2 ? _GEN_863 : _GEN_927; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1439 = _GEN_722[7:6] == 2'h2 ? _GEN_864 : _GEN_928; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1440 = _GEN_722[7:6] == 2'h2 ? _GEN_865 : _GEN_929; // @[d_cache.scala 196:52]
  wire [7:0] _GEN_1441 = _GEN_722[7:6] == 2'h2 ? _GEN_866 : _GEN_930; // @[d_cache.scala 196:52]
  wire  _GEN_1442 = _GEN_722[7:6] == 2'h2 ? dirty_3_0 : _GEN_1278; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1443 = _GEN_722[7:6] == 2'h2 ? dirty_3_1 : _GEN_1279; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1444 = _GEN_722[7:6] == 2'h2 ? dirty_3_2 : _GEN_1280; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1445 = _GEN_722[7:6] == 2'h2 ? dirty_3_3 : _GEN_1281; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1446 = _GEN_722[7:6] == 2'h2 ? dirty_3_4 : _GEN_1282; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1447 = _GEN_722[7:6] == 2'h2 ? dirty_3_5 : _GEN_1283; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1448 = _GEN_722[7:6] == 2'h2 ? dirty_3_6 : _GEN_1284; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1449 = _GEN_722[7:6] == 2'h2 ? dirty_3_7 : _GEN_1285; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1450 = _GEN_722[7:6] == 2'h2 ? dirty_3_8 : _GEN_1286; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1451 = _GEN_722[7:6] == 2'h2 ? dirty_3_9 : _GEN_1287; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1452 = _GEN_722[7:6] == 2'h2 ? dirty_3_10 : _GEN_1288; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1453 = _GEN_722[7:6] == 2'h2 ? dirty_3_11 : _GEN_1289; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1454 = _GEN_722[7:6] == 2'h2 ? dirty_3_12 : _GEN_1290; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1455 = _GEN_722[7:6] == 2'h2 ? dirty_3_13 : _GEN_1291; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1456 = _GEN_722[7:6] == 2'h2 ? dirty_3_14 : _GEN_1292; // @[d_cache.scala 196:52 35:26]
  wire  _GEN_1457 = _GEN_722[7:6] == 2'h2 ? dirty_3_15 : _GEN_1293; // @[d_cache.scala 196:52 35:26]
  wire [127:0] _GEN_1458 = _GEN_722[7:6] == 2'h2 ? ram_3_0 : _GEN_867; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1459 = _GEN_722[7:6] == 2'h2 ? ram_3_1 : _GEN_868; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1460 = _GEN_722[7:6] == 2'h2 ? ram_3_2 : _GEN_869; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1461 = _GEN_722[7:6] == 2'h2 ? ram_3_3 : _GEN_870; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1462 = _GEN_722[7:6] == 2'h2 ? ram_3_4 : _GEN_871; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1463 = _GEN_722[7:6] == 2'h2 ? ram_3_5 : _GEN_872; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1464 = _GEN_722[7:6] == 2'h2 ? ram_3_6 : _GEN_873; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1465 = _GEN_722[7:6] == 2'h2 ? ram_3_7 : _GEN_874; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1466 = _GEN_722[7:6] == 2'h2 ? ram_3_8 : _GEN_875; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1467 = _GEN_722[7:6] == 2'h2 ? ram_3_9 : _GEN_876; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1468 = _GEN_722[7:6] == 2'h2 ? ram_3_10 : _GEN_877; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1469 = _GEN_722[7:6] == 2'h2 ? ram_3_11 : _GEN_878; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1470 = _GEN_722[7:6] == 2'h2 ? ram_3_12 : _GEN_879; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1471 = _GEN_722[7:6] == 2'h2 ? ram_3_13 : _GEN_880; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1472 = _GEN_722[7:6] == 2'h2 ? ram_3_14 : _GEN_881; // @[d_cache.scala 196:52 22:24]
  wire [127:0] _GEN_1473 = _GEN_722[7:6] == 2'h2 ? ram_3_15 : _GEN_882; // @[d_cache.scala 196:52 22:24]
  wire [31:0] _GEN_1474 = _GEN_722[7:6] == 2'h2 ? tag_3_0 : _GEN_883; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1475 = _GEN_722[7:6] == 2'h2 ? tag_3_1 : _GEN_884; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1476 = _GEN_722[7:6] == 2'h2 ? tag_3_2 : _GEN_885; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1477 = _GEN_722[7:6] == 2'h2 ? tag_3_3 : _GEN_886; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1478 = _GEN_722[7:6] == 2'h2 ? tag_3_4 : _GEN_887; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1479 = _GEN_722[7:6] == 2'h2 ? tag_3_5 : _GEN_888; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1480 = _GEN_722[7:6] == 2'h2 ? tag_3_6 : _GEN_889; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1481 = _GEN_722[7:6] == 2'h2 ? tag_3_7 : _GEN_890; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1482 = _GEN_722[7:6] == 2'h2 ? tag_3_8 : _GEN_891; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1483 = _GEN_722[7:6] == 2'h2 ? tag_3_9 : _GEN_892; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1484 = _GEN_722[7:6] == 2'h2 ? tag_3_10 : _GEN_893; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1485 = _GEN_722[7:6] == 2'h2 ? tag_3_11 : _GEN_894; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1486 = _GEN_722[7:6] == 2'h2 ? tag_3_12 : _GEN_895; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1487 = _GEN_722[7:6] == 2'h2 ? tag_3_13 : _GEN_896; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1488 = _GEN_722[7:6] == 2'h2 ? tag_3_14 : _GEN_897; // @[d_cache.scala 196:52 27:24]
  wire [31:0] _GEN_1489 = _GEN_722[7:6] == 2'h2 ? tag_3_15 : _GEN_898; // @[d_cache.scala 196:52 27:24]
  wire  _GEN_1490 = _GEN_722[7:6] == 2'h2 ? valid_3_0 : _GEN_899; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1491 = _GEN_722[7:6] == 2'h2 ? valid_3_1 : _GEN_900; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1492 = _GEN_722[7:6] == 2'h2 ? valid_3_2 : _GEN_901; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1493 = _GEN_722[7:6] == 2'h2 ? valid_3_3 : _GEN_902; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1494 = _GEN_722[7:6] == 2'h2 ? valid_3_4 : _GEN_903; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1495 = _GEN_722[7:6] == 2'h2 ? valid_3_5 : _GEN_904; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1496 = _GEN_722[7:6] == 2'h2 ? valid_3_6 : _GEN_905; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1497 = _GEN_722[7:6] == 2'h2 ? valid_3_7 : _GEN_906; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1498 = _GEN_722[7:6] == 2'h2 ? valid_3_8 : _GEN_907; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1499 = _GEN_722[7:6] == 2'h2 ? valid_3_9 : _GEN_908; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1500 = _GEN_722[7:6] == 2'h2 ? valid_3_10 : _GEN_909; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1501 = _GEN_722[7:6] == 2'h2 ? valid_3_11 : _GEN_910; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1502 = _GEN_722[7:6] == 2'h2 ? valid_3_12 : _GEN_911; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1503 = _GEN_722[7:6] == 2'h2 ? valid_3_13 : _GEN_912; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1504 = _GEN_722[7:6] == 2'h2 ? valid_3_14 : _GEN_913; // @[d_cache.scala 196:52 31:26]
  wire  _GEN_1505 = _GEN_722[7:6] == 2'h2 ? valid_3_15 : _GEN_914; // @[d_cache.scala 196:52 31:26]
  wire [127:0] _GEN_1506 = _GEN_722[7:6] == 2'h1 ? _GEN_1062 : _GEN_1359; // @[d_cache.scala 183:52]
  wire [39:0] _GEN_1507 = _GEN_722[7:6] == 2'h1 ? _GEN_1063 : _GEN_1360; // @[d_cache.scala 183:52]
  wire [3:0] _GEN_1524 = _GEN_722[7:6] == 2'h1 ? _GEN_981 : _GEN_1377; // @[d_cache.scala 183:52]
  wire [127:0] _GEN_1525 = _GEN_722[7:6] == 2'h1 ? _GEN_739 : ram_1_0; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1526 = _GEN_722[7:6] == 2'h1 ? _GEN_740 : ram_1_1; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1527 = _GEN_722[7:6] == 2'h1 ? _GEN_741 : ram_1_2; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1528 = _GEN_722[7:6] == 2'h1 ? _GEN_742 : ram_1_3; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1529 = _GEN_722[7:6] == 2'h1 ? _GEN_743 : ram_1_4; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1530 = _GEN_722[7:6] == 2'h1 ? _GEN_744 : ram_1_5; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1531 = _GEN_722[7:6] == 2'h1 ? _GEN_745 : ram_1_6; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1532 = _GEN_722[7:6] == 2'h1 ? _GEN_746 : ram_1_7; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1533 = _GEN_722[7:6] == 2'h1 ? _GEN_747 : ram_1_8; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1534 = _GEN_722[7:6] == 2'h1 ? _GEN_748 : ram_1_9; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1535 = _GEN_722[7:6] == 2'h1 ? _GEN_749 : ram_1_10; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1536 = _GEN_722[7:6] == 2'h1 ? _GEN_750 : ram_1_11; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1537 = _GEN_722[7:6] == 2'h1 ? _GEN_751 : ram_1_12; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1538 = _GEN_722[7:6] == 2'h1 ? _GEN_752 : ram_1_13; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1539 = _GEN_722[7:6] == 2'h1 ? _GEN_753 : ram_1_14; // @[d_cache.scala 183:52 20:24]
  wire [127:0] _GEN_1540 = _GEN_722[7:6] == 2'h1 ? _GEN_754 : ram_1_15; // @[d_cache.scala 183:52 20:24]
  wire [31:0] _GEN_1541 = _GEN_722[7:6] == 2'h1 ? _GEN_755 : tag_1_0; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1542 = _GEN_722[7:6] == 2'h1 ? _GEN_756 : tag_1_1; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1543 = _GEN_722[7:6] == 2'h1 ? _GEN_757 : tag_1_2; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1544 = _GEN_722[7:6] == 2'h1 ? _GEN_758 : tag_1_3; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1545 = _GEN_722[7:6] == 2'h1 ? _GEN_759 : tag_1_4; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1546 = _GEN_722[7:6] == 2'h1 ? _GEN_760 : tag_1_5; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1547 = _GEN_722[7:6] == 2'h1 ? _GEN_761 : tag_1_6; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1548 = _GEN_722[7:6] == 2'h1 ? _GEN_762 : tag_1_7; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1549 = _GEN_722[7:6] == 2'h1 ? _GEN_763 : tag_1_8; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1550 = _GEN_722[7:6] == 2'h1 ? _GEN_764 : tag_1_9; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1551 = _GEN_722[7:6] == 2'h1 ? _GEN_765 : tag_1_10; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1552 = _GEN_722[7:6] == 2'h1 ? _GEN_766 : tag_1_11; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1553 = _GEN_722[7:6] == 2'h1 ? _GEN_767 : tag_1_12; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1554 = _GEN_722[7:6] == 2'h1 ? _GEN_768 : tag_1_13; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1555 = _GEN_722[7:6] == 2'h1 ? _GEN_769 : tag_1_14; // @[d_cache.scala 183:52 25:24]
  wire [31:0] _GEN_1556 = _GEN_722[7:6] == 2'h1 ? _GEN_770 : tag_1_15; // @[d_cache.scala 183:52 25:24]
  wire  _GEN_1557 = _GEN_722[7:6] == 2'h1 ? _GEN_771 : valid_1_0; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1558 = _GEN_722[7:6] == 2'h1 ? _GEN_772 : valid_1_1; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1559 = _GEN_722[7:6] == 2'h1 ? _GEN_773 : valid_1_2; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1560 = _GEN_722[7:6] == 2'h1 ? _GEN_774 : valid_1_3; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1561 = _GEN_722[7:6] == 2'h1 ? _GEN_775 : valid_1_4; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1562 = _GEN_722[7:6] == 2'h1 ? _GEN_776 : valid_1_5; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1563 = _GEN_722[7:6] == 2'h1 ? _GEN_777 : valid_1_6; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1564 = _GEN_722[7:6] == 2'h1 ? _GEN_778 : valid_1_7; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1565 = _GEN_722[7:6] == 2'h1 ? _GEN_779 : valid_1_8; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1566 = _GEN_722[7:6] == 2'h1 ? _GEN_780 : valid_1_9; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1567 = _GEN_722[7:6] == 2'h1 ? _GEN_781 : valid_1_10; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1568 = _GEN_722[7:6] == 2'h1 ? _GEN_782 : valid_1_11; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1569 = _GEN_722[7:6] == 2'h1 ? _GEN_783 : valid_1_12; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1570 = _GEN_722[7:6] == 2'h1 ? _GEN_784 : valid_1_13; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1571 = _GEN_722[7:6] == 2'h1 ? _GEN_785 : valid_1_14; // @[d_cache.scala 183:52 29:26]
  wire  _GEN_1572 = _GEN_722[7:6] == 2'h1 ? _GEN_786 : valid_1_15; // @[d_cache.scala 183:52 29:26]
  wire [7:0] _GEN_1573 = _GEN_722[7:6] == 2'h1 ? _GEN_787 : _GEN_1426; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1574 = _GEN_722[7:6] == 2'h1 ? _GEN_788 : _GEN_1427; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1575 = _GEN_722[7:6] == 2'h1 ? _GEN_789 : _GEN_1428; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1576 = _GEN_722[7:6] == 2'h1 ? _GEN_790 : _GEN_1429; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1577 = _GEN_722[7:6] == 2'h1 ? _GEN_791 : _GEN_1430; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1578 = _GEN_722[7:6] == 2'h1 ? _GEN_792 : _GEN_1431; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1579 = _GEN_722[7:6] == 2'h1 ? _GEN_793 : _GEN_1432; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1580 = _GEN_722[7:6] == 2'h1 ? _GEN_794 : _GEN_1433; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1581 = _GEN_722[7:6] == 2'h1 ? _GEN_795 : _GEN_1434; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1582 = _GEN_722[7:6] == 2'h1 ? _GEN_796 : _GEN_1435; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1583 = _GEN_722[7:6] == 2'h1 ? _GEN_797 : _GEN_1436; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1584 = _GEN_722[7:6] == 2'h1 ? _GEN_798 : _GEN_1437; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1585 = _GEN_722[7:6] == 2'h1 ? _GEN_799 : _GEN_1438; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1586 = _GEN_722[7:6] == 2'h1 ? _GEN_800 : _GEN_1439; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1587 = _GEN_722[7:6] == 2'h1 ? _GEN_801 : _GEN_1440; // @[d_cache.scala 183:52]
  wire [7:0] _GEN_1588 = _GEN_722[7:6] == 2'h1 ? _GEN_802 : _GEN_1441; // @[d_cache.scala 183:52]
  wire [127:0] _GEN_1605 = _GEN_722[7:6] == 2'h1 ? ram_2_0 : _GEN_1378; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1606 = _GEN_722[7:6] == 2'h1 ? ram_2_1 : _GEN_1379; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1607 = _GEN_722[7:6] == 2'h1 ? ram_2_2 : _GEN_1380; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1608 = _GEN_722[7:6] == 2'h1 ? ram_2_3 : _GEN_1381; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1609 = _GEN_722[7:6] == 2'h1 ? ram_2_4 : _GEN_1382; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1610 = _GEN_722[7:6] == 2'h1 ? ram_2_5 : _GEN_1383; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1611 = _GEN_722[7:6] == 2'h1 ? ram_2_6 : _GEN_1384; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1612 = _GEN_722[7:6] == 2'h1 ? ram_2_7 : _GEN_1385; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1613 = _GEN_722[7:6] == 2'h1 ? ram_2_8 : _GEN_1386; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1614 = _GEN_722[7:6] == 2'h1 ? ram_2_9 : _GEN_1387; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1615 = _GEN_722[7:6] == 2'h1 ? ram_2_10 : _GEN_1388; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1616 = _GEN_722[7:6] == 2'h1 ? ram_2_11 : _GEN_1389; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1617 = _GEN_722[7:6] == 2'h1 ? ram_2_12 : _GEN_1390; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1618 = _GEN_722[7:6] == 2'h1 ? ram_2_13 : _GEN_1391; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1619 = _GEN_722[7:6] == 2'h1 ? ram_2_14 : _GEN_1392; // @[d_cache.scala 183:52 21:24]
  wire [127:0] _GEN_1620 = _GEN_722[7:6] == 2'h1 ? ram_2_15 : _GEN_1393; // @[d_cache.scala 183:52 21:24]
  wire [31:0] _GEN_1621 = _GEN_722[7:6] == 2'h1 ? tag_2_0 : _GEN_1394; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1622 = _GEN_722[7:6] == 2'h1 ? tag_2_1 : _GEN_1395; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1623 = _GEN_722[7:6] == 2'h1 ? tag_2_2 : _GEN_1396; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1624 = _GEN_722[7:6] == 2'h1 ? tag_2_3 : _GEN_1397; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1625 = _GEN_722[7:6] == 2'h1 ? tag_2_4 : _GEN_1398; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1626 = _GEN_722[7:6] == 2'h1 ? tag_2_5 : _GEN_1399; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1627 = _GEN_722[7:6] == 2'h1 ? tag_2_6 : _GEN_1400; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1628 = _GEN_722[7:6] == 2'h1 ? tag_2_7 : _GEN_1401; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1629 = _GEN_722[7:6] == 2'h1 ? tag_2_8 : _GEN_1402; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1630 = _GEN_722[7:6] == 2'h1 ? tag_2_9 : _GEN_1403; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1631 = _GEN_722[7:6] == 2'h1 ? tag_2_10 : _GEN_1404; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1632 = _GEN_722[7:6] == 2'h1 ? tag_2_11 : _GEN_1405; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1633 = _GEN_722[7:6] == 2'h1 ? tag_2_12 : _GEN_1406; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1634 = _GEN_722[7:6] == 2'h1 ? tag_2_13 : _GEN_1407; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1635 = _GEN_722[7:6] == 2'h1 ? tag_2_14 : _GEN_1408; // @[d_cache.scala 183:52 26:24]
  wire [31:0] _GEN_1636 = _GEN_722[7:6] == 2'h1 ? tag_2_15 : _GEN_1409; // @[d_cache.scala 183:52 26:24]
  wire  _GEN_1637 = _GEN_722[7:6] == 2'h1 ? valid_2_0 : _GEN_1410; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1638 = _GEN_722[7:6] == 2'h1 ? valid_2_1 : _GEN_1411; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1639 = _GEN_722[7:6] == 2'h1 ? valid_2_2 : _GEN_1412; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1640 = _GEN_722[7:6] == 2'h1 ? valid_2_3 : _GEN_1413; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1641 = _GEN_722[7:6] == 2'h1 ? valid_2_4 : _GEN_1414; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1642 = _GEN_722[7:6] == 2'h1 ? valid_2_5 : _GEN_1415; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1643 = _GEN_722[7:6] == 2'h1 ? valid_2_6 : _GEN_1416; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1644 = _GEN_722[7:6] == 2'h1 ? valid_2_7 : _GEN_1417; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1645 = _GEN_722[7:6] == 2'h1 ? valid_2_8 : _GEN_1418; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1646 = _GEN_722[7:6] == 2'h1 ? valid_2_9 : _GEN_1419; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1647 = _GEN_722[7:6] == 2'h1 ? valid_2_10 : _GEN_1420; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1648 = _GEN_722[7:6] == 2'h1 ? valid_2_11 : _GEN_1421; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1649 = _GEN_722[7:6] == 2'h1 ? valid_2_12 : _GEN_1422; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1650 = _GEN_722[7:6] == 2'h1 ? valid_2_13 : _GEN_1423; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1651 = _GEN_722[7:6] == 2'h1 ? valid_2_14 : _GEN_1424; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1652 = _GEN_722[7:6] == 2'h1 ? valid_2_15 : _GEN_1425; // @[d_cache.scala 183:52 30:26]
  wire  _GEN_1653 = _GEN_722[7:6] == 2'h1 ? dirty_3_0 : _GEN_1442; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1654 = _GEN_722[7:6] == 2'h1 ? dirty_3_1 : _GEN_1443; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1655 = _GEN_722[7:6] == 2'h1 ? dirty_3_2 : _GEN_1444; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1656 = _GEN_722[7:6] == 2'h1 ? dirty_3_3 : _GEN_1445; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1657 = _GEN_722[7:6] == 2'h1 ? dirty_3_4 : _GEN_1446; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1658 = _GEN_722[7:6] == 2'h1 ? dirty_3_5 : _GEN_1447; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1659 = _GEN_722[7:6] == 2'h1 ? dirty_3_6 : _GEN_1448; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1660 = _GEN_722[7:6] == 2'h1 ? dirty_3_7 : _GEN_1449; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1661 = _GEN_722[7:6] == 2'h1 ? dirty_3_8 : _GEN_1450; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1662 = _GEN_722[7:6] == 2'h1 ? dirty_3_9 : _GEN_1451; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1663 = _GEN_722[7:6] == 2'h1 ? dirty_3_10 : _GEN_1452; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1664 = _GEN_722[7:6] == 2'h1 ? dirty_3_11 : _GEN_1453; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1665 = _GEN_722[7:6] == 2'h1 ? dirty_3_12 : _GEN_1454; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1666 = _GEN_722[7:6] == 2'h1 ? dirty_3_13 : _GEN_1455; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1667 = _GEN_722[7:6] == 2'h1 ? dirty_3_14 : _GEN_1456; // @[d_cache.scala 183:52 35:26]
  wire  _GEN_1668 = _GEN_722[7:6] == 2'h1 ? dirty_3_15 : _GEN_1457; // @[d_cache.scala 183:52 35:26]
  wire [127:0] _GEN_1669 = _GEN_722[7:6] == 2'h1 ? ram_3_0 : _GEN_1458; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1670 = _GEN_722[7:6] == 2'h1 ? ram_3_1 : _GEN_1459; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1671 = _GEN_722[7:6] == 2'h1 ? ram_3_2 : _GEN_1460; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1672 = _GEN_722[7:6] == 2'h1 ? ram_3_3 : _GEN_1461; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1673 = _GEN_722[7:6] == 2'h1 ? ram_3_4 : _GEN_1462; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1674 = _GEN_722[7:6] == 2'h1 ? ram_3_5 : _GEN_1463; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1675 = _GEN_722[7:6] == 2'h1 ? ram_3_6 : _GEN_1464; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1676 = _GEN_722[7:6] == 2'h1 ? ram_3_7 : _GEN_1465; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1677 = _GEN_722[7:6] == 2'h1 ? ram_3_8 : _GEN_1466; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1678 = _GEN_722[7:6] == 2'h1 ? ram_3_9 : _GEN_1467; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1679 = _GEN_722[7:6] == 2'h1 ? ram_3_10 : _GEN_1468; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1680 = _GEN_722[7:6] == 2'h1 ? ram_3_11 : _GEN_1469; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1681 = _GEN_722[7:6] == 2'h1 ? ram_3_12 : _GEN_1470; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1682 = _GEN_722[7:6] == 2'h1 ? ram_3_13 : _GEN_1471; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1683 = _GEN_722[7:6] == 2'h1 ? ram_3_14 : _GEN_1472; // @[d_cache.scala 183:52 22:24]
  wire [127:0] _GEN_1684 = _GEN_722[7:6] == 2'h1 ? ram_3_15 : _GEN_1473; // @[d_cache.scala 183:52 22:24]
  wire [31:0] _GEN_1685 = _GEN_722[7:6] == 2'h1 ? tag_3_0 : _GEN_1474; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1686 = _GEN_722[7:6] == 2'h1 ? tag_3_1 : _GEN_1475; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1687 = _GEN_722[7:6] == 2'h1 ? tag_3_2 : _GEN_1476; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1688 = _GEN_722[7:6] == 2'h1 ? tag_3_3 : _GEN_1477; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1689 = _GEN_722[7:6] == 2'h1 ? tag_3_4 : _GEN_1478; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1690 = _GEN_722[7:6] == 2'h1 ? tag_3_5 : _GEN_1479; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1691 = _GEN_722[7:6] == 2'h1 ? tag_3_6 : _GEN_1480; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1692 = _GEN_722[7:6] == 2'h1 ? tag_3_7 : _GEN_1481; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1693 = _GEN_722[7:6] == 2'h1 ? tag_3_8 : _GEN_1482; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1694 = _GEN_722[7:6] == 2'h1 ? tag_3_9 : _GEN_1483; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1695 = _GEN_722[7:6] == 2'h1 ? tag_3_10 : _GEN_1484; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1696 = _GEN_722[7:6] == 2'h1 ? tag_3_11 : _GEN_1485; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1697 = _GEN_722[7:6] == 2'h1 ? tag_3_12 : _GEN_1486; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1698 = _GEN_722[7:6] == 2'h1 ? tag_3_13 : _GEN_1487; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1699 = _GEN_722[7:6] == 2'h1 ? tag_3_14 : _GEN_1488; // @[d_cache.scala 183:52 27:24]
  wire [31:0] _GEN_1700 = _GEN_722[7:6] == 2'h1 ? tag_3_15 : _GEN_1489; // @[d_cache.scala 183:52 27:24]
  wire  _GEN_1701 = _GEN_722[7:6] == 2'h1 ? valid_3_0 : _GEN_1490; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1702 = _GEN_722[7:6] == 2'h1 ? valid_3_1 : _GEN_1491; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1703 = _GEN_722[7:6] == 2'h1 ? valid_3_2 : _GEN_1492; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1704 = _GEN_722[7:6] == 2'h1 ? valid_3_3 : _GEN_1493; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1705 = _GEN_722[7:6] == 2'h1 ? valid_3_4 : _GEN_1494; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1706 = _GEN_722[7:6] == 2'h1 ? valid_3_5 : _GEN_1495; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1707 = _GEN_722[7:6] == 2'h1 ? valid_3_6 : _GEN_1496; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1708 = _GEN_722[7:6] == 2'h1 ? valid_3_7 : _GEN_1497; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1709 = _GEN_722[7:6] == 2'h1 ? valid_3_8 : _GEN_1498; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1710 = _GEN_722[7:6] == 2'h1 ? valid_3_9 : _GEN_1499; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1711 = _GEN_722[7:6] == 2'h1 ? valid_3_10 : _GEN_1500; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1712 = _GEN_722[7:6] == 2'h1 ? valid_3_11 : _GEN_1501; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1713 = _GEN_722[7:6] == 2'h1 ? valid_3_12 : _GEN_1502; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1714 = _GEN_722[7:6] == 2'h1 ? valid_3_13 : _GEN_1503; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1715 = _GEN_722[7:6] == 2'h1 ? valid_3_14 : _GEN_1504; // @[d_cache.scala 183:52 31:26]
  wire  _GEN_1716 = _GEN_722[7:6] == 2'h1 ? valid_3_15 : _GEN_1505; // @[d_cache.scala 183:52 31:26]
  wire [127:0] _GEN_1717 = _GEN_722[7:6] == 2'h0 ? _GEN_963 : _GEN_1506; // @[d_cache.scala 169:46]
  wire [39:0] _GEN_1718 = _GEN_722[7:6] == 2'h0 ? _GEN_964 : _GEN_1507; // @[d_cache.scala 169:46]
  wire  _GEN_1719 = _GEN_722[7:6] == 2'h0 ? _GEN_965 : dirty_0_0; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1720 = _GEN_722[7:6] == 2'h0 ? _GEN_966 : dirty_0_1; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1721 = _GEN_722[7:6] == 2'h0 ? _GEN_967 : dirty_0_2; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1722 = _GEN_722[7:6] == 2'h0 ? _GEN_968 : dirty_0_3; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1723 = _GEN_722[7:6] == 2'h0 ? _GEN_969 : dirty_0_4; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1724 = _GEN_722[7:6] == 2'h0 ? _GEN_970 : dirty_0_5; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1725 = _GEN_722[7:6] == 2'h0 ? _GEN_971 : dirty_0_6; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1726 = _GEN_722[7:6] == 2'h0 ? _GEN_972 : dirty_0_7; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1727 = _GEN_722[7:6] == 2'h0 ? _GEN_973 : dirty_0_8; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1728 = _GEN_722[7:6] == 2'h0 ? _GEN_974 : dirty_0_9; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1729 = _GEN_722[7:6] == 2'h0 ? _GEN_975 : dirty_0_10; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1730 = _GEN_722[7:6] == 2'h0 ? _GEN_976 : dirty_0_11; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1731 = _GEN_722[7:6] == 2'h0 ? _GEN_977 : dirty_0_12; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1732 = _GEN_722[7:6] == 2'h0 ? _GEN_978 : dirty_0_13; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1733 = _GEN_722[7:6] == 2'h0 ? _GEN_979 : dirty_0_14; // @[d_cache.scala 169:46 32:26]
  wire  _GEN_1734 = _GEN_722[7:6] == 2'h0 ? _GEN_980 : dirty_0_15; // @[d_cache.scala 169:46 32:26]
  wire [3:0] _GEN_1735 = _GEN_722[7:6] == 2'h0 ? _GEN_981 : _GEN_1524; // @[d_cache.scala 169:46]
  wire [127:0] _GEN_1736 = _GEN_722[7:6] == 2'h0 ? _GEN_659 : ram_0_0; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1737 = _GEN_722[7:6] == 2'h0 ? _GEN_660 : ram_0_1; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1738 = _GEN_722[7:6] == 2'h0 ? _GEN_661 : ram_0_2; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1739 = _GEN_722[7:6] == 2'h0 ? _GEN_662 : ram_0_3; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1740 = _GEN_722[7:6] == 2'h0 ? _GEN_663 : ram_0_4; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1741 = _GEN_722[7:6] == 2'h0 ? _GEN_664 : ram_0_5; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1742 = _GEN_722[7:6] == 2'h0 ? _GEN_665 : ram_0_6; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1743 = _GEN_722[7:6] == 2'h0 ? _GEN_666 : ram_0_7; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1744 = _GEN_722[7:6] == 2'h0 ? _GEN_667 : ram_0_8; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1745 = _GEN_722[7:6] == 2'h0 ? _GEN_668 : ram_0_9; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1746 = _GEN_722[7:6] == 2'h0 ? _GEN_669 : ram_0_10; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1747 = _GEN_722[7:6] == 2'h0 ? _GEN_670 : ram_0_11; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1748 = _GEN_722[7:6] == 2'h0 ? _GEN_671 : ram_0_12; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1749 = _GEN_722[7:6] == 2'h0 ? _GEN_672 : ram_0_13; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1750 = _GEN_722[7:6] == 2'h0 ? _GEN_673 : ram_0_14; // @[d_cache.scala 169:46 19:24]
  wire [127:0] _GEN_1751 = _GEN_722[7:6] == 2'h0 ? _GEN_674 : ram_0_15; // @[d_cache.scala 169:46 19:24]
  wire [31:0] _GEN_1752 = _GEN_722[7:6] == 2'h0 ? _GEN_675 : tag_0_0; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1753 = _GEN_722[7:6] == 2'h0 ? _GEN_676 : tag_0_1; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1754 = _GEN_722[7:6] == 2'h0 ? _GEN_677 : tag_0_2; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1755 = _GEN_722[7:6] == 2'h0 ? _GEN_678 : tag_0_3; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1756 = _GEN_722[7:6] == 2'h0 ? _GEN_679 : tag_0_4; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1757 = _GEN_722[7:6] == 2'h0 ? _GEN_680 : tag_0_5; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1758 = _GEN_722[7:6] == 2'h0 ? _GEN_681 : tag_0_6; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1759 = _GEN_722[7:6] == 2'h0 ? _GEN_682 : tag_0_7; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1760 = _GEN_722[7:6] == 2'h0 ? _GEN_683 : tag_0_8; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1761 = _GEN_722[7:6] == 2'h0 ? _GEN_684 : tag_0_9; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1762 = _GEN_722[7:6] == 2'h0 ? _GEN_685 : tag_0_10; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1763 = _GEN_722[7:6] == 2'h0 ? _GEN_686 : tag_0_11; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1764 = _GEN_722[7:6] == 2'h0 ? _GEN_687 : tag_0_12; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1765 = _GEN_722[7:6] == 2'h0 ? _GEN_688 : tag_0_13; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1766 = _GEN_722[7:6] == 2'h0 ? _GEN_689 : tag_0_14; // @[d_cache.scala 169:46 24:24]
  wire [31:0] _GEN_1767 = _GEN_722[7:6] == 2'h0 ? _GEN_690 : tag_0_15; // @[d_cache.scala 169:46 24:24]
  wire  _GEN_1768 = _GEN_722[7:6] == 2'h0 ? _GEN_691 : valid_0_0; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1769 = _GEN_722[7:6] == 2'h0 ? _GEN_692 : valid_0_1; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1770 = _GEN_722[7:6] == 2'h0 ? _GEN_693 : valid_0_2; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1771 = _GEN_722[7:6] == 2'h0 ? _GEN_694 : valid_0_3; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1772 = _GEN_722[7:6] == 2'h0 ? _GEN_695 : valid_0_4; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1773 = _GEN_722[7:6] == 2'h0 ? _GEN_696 : valid_0_5; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1774 = _GEN_722[7:6] == 2'h0 ? _GEN_697 : valid_0_6; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1775 = _GEN_722[7:6] == 2'h0 ? _GEN_698 : valid_0_7; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1776 = _GEN_722[7:6] == 2'h0 ? _GEN_699 : valid_0_8; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1777 = _GEN_722[7:6] == 2'h0 ? _GEN_700 : valid_0_9; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1778 = _GEN_722[7:6] == 2'h0 ? _GEN_701 : valid_0_10; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1779 = _GEN_722[7:6] == 2'h0 ? _GEN_702 : valid_0_11; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1780 = _GEN_722[7:6] == 2'h0 ? _GEN_703 : valid_0_12; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1781 = _GEN_722[7:6] == 2'h0 ? _GEN_704 : valid_0_13; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1782 = _GEN_722[7:6] == 2'h0 ? _GEN_705 : valid_0_14; // @[d_cache.scala 169:46 28:26]
  wire  _GEN_1783 = _GEN_722[7:6] == 2'h0 ? _GEN_706 : valid_0_15; // @[d_cache.scala 169:46 28:26]
  wire [7:0] _GEN_1784 = _GEN_722[7:6] == 2'h0 ? _GEN_723 : _GEN_1573; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1785 = _GEN_722[7:6] == 2'h0 ? _GEN_724 : _GEN_1574; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1786 = _GEN_722[7:6] == 2'h0 ? _GEN_725 : _GEN_1575; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1787 = _GEN_722[7:6] == 2'h0 ? _GEN_726 : _GEN_1576; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1788 = _GEN_722[7:6] == 2'h0 ? _GEN_727 : _GEN_1577; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1789 = _GEN_722[7:6] == 2'h0 ? _GEN_728 : _GEN_1578; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1790 = _GEN_722[7:6] == 2'h0 ? _GEN_729 : _GEN_1579; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1791 = _GEN_722[7:6] == 2'h0 ? _GEN_730 : _GEN_1580; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1792 = _GEN_722[7:6] == 2'h0 ? _GEN_731 : _GEN_1581; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1793 = _GEN_722[7:6] == 2'h0 ? _GEN_732 : _GEN_1582; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1794 = _GEN_722[7:6] == 2'h0 ? _GEN_733 : _GEN_1583; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1795 = _GEN_722[7:6] == 2'h0 ? _GEN_734 : _GEN_1584; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1796 = _GEN_722[7:6] == 2'h0 ? _GEN_735 : _GEN_1585; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1797 = _GEN_722[7:6] == 2'h0 ? _GEN_736 : _GEN_1586; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1798 = _GEN_722[7:6] == 2'h0 ? _GEN_737 : _GEN_1587; // @[d_cache.scala 169:46]
  wire [7:0] _GEN_1799 = _GEN_722[7:6] == 2'h0 ? _GEN_738 : _GEN_1588; // @[d_cache.scala 169:46]
  wire [127:0] _GEN_1816 = _GEN_722[7:6] == 2'h0 ? ram_1_0 : _GEN_1525; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1817 = _GEN_722[7:6] == 2'h0 ? ram_1_1 : _GEN_1526; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1818 = _GEN_722[7:6] == 2'h0 ? ram_1_2 : _GEN_1527; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1819 = _GEN_722[7:6] == 2'h0 ? ram_1_3 : _GEN_1528; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1820 = _GEN_722[7:6] == 2'h0 ? ram_1_4 : _GEN_1529; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1821 = _GEN_722[7:6] == 2'h0 ? ram_1_5 : _GEN_1530; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1822 = _GEN_722[7:6] == 2'h0 ? ram_1_6 : _GEN_1531; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1823 = _GEN_722[7:6] == 2'h0 ? ram_1_7 : _GEN_1532; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1824 = _GEN_722[7:6] == 2'h0 ? ram_1_8 : _GEN_1533; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1825 = _GEN_722[7:6] == 2'h0 ? ram_1_9 : _GEN_1534; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1826 = _GEN_722[7:6] == 2'h0 ? ram_1_10 : _GEN_1535; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1827 = _GEN_722[7:6] == 2'h0 ? ram_1_11 : _GEN_1536; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1828 = _GEN_722[7:6] == 2'h0 ? ram_1_12 : _GEN_1537; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1829 = _GEN_722[7:6] == 2'h0 ? ram_1_13 : _GEN_1538; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1830 = _GEN_722[7:6] == 2'h0 ? ram_1_14 : _GEN_1539; // @[d_cache.scala 169:46 20:24]
  wire [127:0] _GEN_1831 = _GEN_722[7:6] == 2'h0 ? ram_1_15 : _GEN_1540; // @[d_cache.scala 169:46 20:24]
  wire [31:0] _GEN_1832 = _GEN_722[7:6] == 2'h0 ? tag_1_0 : _GEN_1541; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1833 = _GEN_722[7:6] == 2'h0 ? tag_1_1 : _GEN_1542; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1834 = _GEN_722[7:6] == 2'h0 ? tag_1_2 : _GEN_1543; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1835 = _GEN_722[7:6] == 2'h0 ? tag_1_3 : _GEN_1544; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1836 = _GEN_722[7:6] == 2'h0 ? tag_1_4 : _GEN_1545; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1837 = _GEN_722[7:6] == 2'h0 ? tag_1_5 : _GEN_1546; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1838 = _GEN_722[7:6] == 2'h0 ? tag_1_6 : _GEN_1547; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1839 = _GEN_722[7:6] == 2'h0 ? tag_1_7 : _GEN_1548; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1840 = _GEN_722[7:6] == 2'h0 ? tag_1_8 : _GEN_1549; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1841 = _GEN_722[7:6] == 2'h0 ? tag_1_9 : _GEN_1550; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1842 = _GEN_722[7:6] == 2'h0 ? tag_1_10 : _GEN_1551; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1843 = _GEN_722[7:6] == 2'h0 ? tag_1_11 : _GEN_1552; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1844 = _GEN_722[7:6] == 2'h0 ? tag_1_12 : _GEN_1553; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1845 = _GEN_722[7:6] == 2'h0 ? tag_1_13 : _GEN_1554; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1846 = _GEN_722[7:6] == 2'h0 ? tag_1_14 : _GEN_1555; // @[d_cache.scala 169:46 25:24]
  wire [31:0] _GEN_1847 = _GEN_722[7:6] == 2'h0 ? tag_1_15 : _GEN_1556; // @[d_cache.scala 169:46 25:24]
  wire  _GEN_1848 = _GEN_722[7:6] == 2'h0 ? valid_1_0 : _GEN_1557; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1849 = _GEN_722[7:6] == 2'h0 ? valid_1_1 : _GEN_1558; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1850 = _GEN_722[7:6] == 2'h0 ? valid_1_2 : _GEN_1559; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1851 = _GEN_722[7:6] == 2'h0 ? valid_1_3 : _GEN_1560; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1852 = _GEN_722[7:6] == 2'h0 ? valid_1_4 : _GEN_1561; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1853 = _GEN_722[7:6] == 2'h0 ? valid_1_5 : _GEN_1562; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1854 = _GEN_722[7:6] == 2'h0 ? valid_1_6 : _GEN_1563; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1855 = _GEN_722[7:6] == 2'h0 ? valid_1_7 : _GEN_1564; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1856 = _GEN_722[7:6] == 2'h0 ? valid_1_8 : _GEN_1565; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1857 = _GEN_722[7:6] == 2'h0 ? valid_1_9 : _GEN_1566; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1858 = _GEN_722[7:6] == 2'h0 ? valid_1_10 : _GEN_1567; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1859 = _GEN_722[7:6] == 2'h0 ? valid_1_11 : _GEN_1568; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1860 = _GEN_722[7:6] == 2'h0 ? valid_1_12 : _GEN_1569; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1861 = _GEN_722[7:6] == 2'h0 ? valid_1_13 : _GEN_1570; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1862 = _GEN_722[7:6] == 2'h0 ? valid_1_14 : _GEN_1571; // @[d_cache.scala 169:46 29:26]
  wire  _GEN_1863 = _GEN_722[7:6] == 2'h0 ? valid_1_15 : _GEN_1572; // @[d_cache.scala 169:46 29:26]
  wire [127:0] _GEN_1880 = _GEN_722[7:6] == 2'h0 ? ram_2_0 : _GEN_1605; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1881 = _GEN_722[7:6] == 2'h0 ? ram_2_1 : _GEN_1606; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1882 = _GEN_722[7:6] == 2'h0 ? ram_2_2 : _GEN_1607; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1883 = _GEN_722[7:6] == 2'h0 ? ram_2_3 : _GEN_1608; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1884 = _GEN_722[7:6] == 2'h0 ? ram_2_4 : _GEN_1609; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1885 = _GEN_722[7:6] == 2'h0 ? ram_2_5 : _GEN_1610; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1886 = _GEN_722[7:6] == 2'h0 ? ram_2_6 : _GEN_1611; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1887 = _GEN_722[7:6] == 2'h0 ? ram_2_7 : _GEN_1612; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1888 = _GEN_722[7:6] == 2'h0 ? ram_2_8 : _GEN_1613; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1889 = _GEN_722[7:6] == 2'h0 ? ram_2_9 : _GEN_1614; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1890 = _GEN_722[7:6] == 2'h0 ? ram_2_10 : _GEN_1615; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1891 = _GEN_722[7:6] == 2'h0 ? ram_2_11 : _GEN_1616; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1892 = _GEN_722[7:6] == 2'h0 ? ram_2_12 : _GEN_1617; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1893 = _GEN_722[7:6] == 2'h0 ? ram_2_13 : _GEN_1618; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1894 = _GEN_722[7:6] == 2'h0 ? ram_2_14 : _GEN_1619; // @[d_cache.scala 169:46 21:24]
  wire [127:0] _GEN_1895 = _GEN_722[7:6] == 2'h0 ? ram_2_15 : _GEN_1620; // @[d_cache.scala 169:46 21:24]
  wire [31:0] _GEN_1896 = _GEN_722[7:6] == 2'h0 ? tag_2_0 : _GEN_1621; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1897 = _GEN_722[7:6] == 2'h0 ? tag_2_1 : _GEN_1622; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1898 = _GEN_722[7:6] == 2'h0 ? tag_2_2 : _GEN_1623; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1899 = _GEN_722[7:6] == 2'h0 ? tag_2_3 : _GEN_1624; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1900 = _GEN_722[7:6] == 2'h0 ? tag_2_4 : _GEN_1625; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1901 = _GEN_722[7:6] == 2'h0 ? tag_2_5 : _GEN_1626; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1902 = _GEN_722[7:6] == 2'h0 ? tag_2_6 : _GEN_1627; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1903 = _GEN_722[7:6] == 2'h0 ? tag_2_7 : _GEN_1628; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1904 = _GEN_722[7:6] == 2'h0 ? tag_2_8 : _GEN_1629; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1905 = _GEN_722[7:6] == 2'h0 ? tag_2_9 : _GEN_1630; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1906 = _GEN_722[7:6] == 2'h0 ? tag_2_10 : _GEN_1631; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1907 = _GEN_722[7:6] == 2'h0 ? tag_2_11 : _GEN_1632; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1908 = _GEN_722[7:6] == 2'h0 ? tag_2_12 : _GEN_1633; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1909 = _GEN_722[7:6] == 2'h0 ? tag_2_13 : _GEN_1634; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1910 = _GEN_722[7:6] == 2'h0 ? tag_2_14 : _GEN_1635; // @[d_cache.scala 169:46 26:24]
  wire [31:0] _GEN_1911 = _GEN_722[7:6] == 2'h0 ? tag_2_15 : _GEN_1636; // @[d_cache.scala 169:46 26:24]
  wire  _GEN_1912 = _GEN_722[7:6] == 2'h0 ? valid_2_0 : _GEN_1637; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1913 = _GEN_722[7:6] == 2'h0 ? valid_2_1 : _GEN_1638; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1914 = _GEN_722[7:6] == 2'h0 ? valid_2_2 : _GEN_1639; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1915 = _GEN_722[7:6] == 2'h0 ? valid_2_3 : _GEN_1640; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1916 = _GEN_722[7:6] == 2'h0 ? valid_2_4 : _GEN_1641; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1917 = _GEN_722[7:6] == 2'h0 ? valid_2_5 : _GEN_1642; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1918 = _GEN_722[7:6] == 2'h0 ? valid_2_6 : _GEN_1643; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1919 = _GEN_722[7:6] == 2'h0 ? valid_2_7 : _GEN_1644; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1920 = _GEN_722[7:6] == 2'h0 ? valid_2_8 : _GEN_1645; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1921 = _GEN_722[7:6] == 2'h0 ? valid_2_9 : _GEN_1646; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1922 = _GEN_722[7:6] == 2'h0 ? valid_2_10 : _GEN_1647; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1923 = _GEN_722[7:6] == 2'h0 ? valid_2_11 : _GEN_1648; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1924 = _GEN_722[7:6] == 2'h0 ? valid_2_12 : _GEN_1649; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1925 = _GEN_722[7:6] == 2'h0 ? valid_2_13 : _GEN_1650; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1926 = _GEN_722[7:6] == 2'h0 ? valid_2_14 : _GEN_1651; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1927 = _GEN_722[7:6] == 2'h0 ? valid_2_15 : _GEN_1652; // @[d_cache.scala 169:46 30:26]
  wire  _GEN_1928 = _GEN_722[7:6] == 2'h0 ? dirty_3_0 : _GEN_1653; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1929 = _GEN_722[7:6] == 2'h0 ? dirty_3_1 : _GEN_1654; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1930 = _GEN_722[7:6] == 2'h0 ? dirty_3_2 : _GEN_1655; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1931 = _GEN_722[7:6] == 2'h0 ? dirty_3_3 : _GEN_1656; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1932 = _GEN_722[7:6] == 2'h0 ? dirty_3_4 : _GEN_1657; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1933 = _GEN_722[7:6] == 2'h0 ? dirty_3_5 : _GEN_1658; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1934 = _GEN_722[7:6] == 2'h0 ? dirty_3_6 : _GEN_1659; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1935 = _GEN_722[7:6] == 2'h0 ? dirty_3_7 : _GEN_1660; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1936 = _GEN_722[7:6] == 2'h0 ? dirty_3_8 : _GEN_1661; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1937 = _GEN_722[7:6] == 2'h0 ? dirty_3_9 : _GEN_1662; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1938 = _GEN_722[7:6] == 2'h0 ? dirty_3_10 : _GEN_1663; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1939 = _GEN_722[7:6] == 2'h0 ? dirty_3_11 : _GEN_1664; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1940 = _GEN_722[7:6] == 2'h0 ? dirty_3_12 : _GEN_1665; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1941 = _GEN_722[7:6] == 2'h0 ? dirty_3_13 : _GEN_1666; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1942 = _GEN_722[7:6] == 2'h0 ? dirty_3_14 : _GEN_1667; // @[d_cache.scala 169:46 35:26]
  wire  _GEN_1943 = _GEN_722[7:6] == 2'h0 ? dirty_3_15 : _GEN_1668; // @[d_cache.scala 169:46 35:26]
  wire [127:0] _GEN_1944 = _GEN_722[7:6] == 2'h0 ? ram_3_0 : _GEN_1669; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1945 = _GEN_722[7:6] == 2'h0 ? ram_3_1 : _GEN_1670; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1946 = _GEN_722[7:6] == 2'h0 ? ram_3_2 : _GEN_1671; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1947 = _GEN_722[7:6] == 2'h0 ? ram_3_3 : _GEN_1672; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1948 = _GEN_722[7:6] == 2'h0 ? ram_3_4 : _GEN_1673; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1949 = _GEN_722[7:6] == 2'h0 ? ram_3_5 : _GEN_1674; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1950 = _GEN_722[7:6] == 2'h0 ? ram_3_6 : _GEN_1675; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1951 = _GEN_722[7:6] == 2'h0 ? ram_3_7 : _GEN_1676; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1952 = _GEN_722[7:6] == 2'h0 ? ram_3_8 : _GEN_1677; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1953 = _GEN_722[7:6] == 2'h0 ? ram_3_9 : _GEN_1678; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1954 = _GEN_722[7:6] == 2'h0 ? ram_3_10 : _GEN_1679; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1955 = _GEN_722[7:6] == 2'h0 ? ram_3_11 : _GEN_1680; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1956 = _GEN_722[7:6] == 2'h0 ? ram_3_12 : _GEN_1681; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1957 = _GEN_722[7:6] == 2'h0 ? ram_3_13 : _GEN_1682; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1958 = _GEN_722[7:6] == 2'h0 ? ram_3_14 : _GEN_1683; // @[d_cache.scala 169:46 22:24]
  wire [127:0] _GEN_1959 = _GEN_722[7:6] == 2'h0 ? ram_3_15 : _GEN_1684; // @[d_cache.scala 169:46 22:24]
  wire [31:0] _GEN_1960 = _GEN_722[7:6] == 2'h0 ? tag_3_0 : _GEN_1685; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1961 = _GEN_722[7:6] == 2'h0 ? tag_3_1 : _GEN_1686; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1962 = _GEN_722[7:6] == 2'h0 ? tag_3_2 : _GEN_1687; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1963 = _GEN_722[7:6] == 2'h0 ? tag_3_3 : _GEN_1688; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1964 = _GEN_722[7:6] == 2'h0 ? tag_3_4 : _GEN_1689; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1965 = _GEN_722[7:6] == 2'h0 ? tag_3_5 : _GEN_1690; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1966 = _GEN_722[7:6] == 2'h0 ? tag_3_6 : _GEN_1691; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1967 = _GEN_722[7:6] == 2'h0 ? tag_3_7 : _GEN_1692; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1968 = _GEN_722[7:6] == 2'h0 ? tag_3_8 : _GEN_1693; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1969 = _GEN_722[7:6] == 2'h0 ? tag_3_9 : _GEN_1694; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1970 = _GEN_722[7:6] == 2'h0 ? tag_3_10 : _GEN_1695; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1971 = _GEN_722[7:6] == 2'h0 ? tag_3_11 : _GEN_1696; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1972 = _GEN_722[7:6] == 2'h0 ? tag_3_12 : _GEN_1697; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1973 = _GEN_722[7:6] == 2'h0 ? tag_3_13 : _GEN_1698; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1974 = _GEN_722[7:6] == 2'h0 ? tag_3_14 : _GEN_1699; // @[d_cache.scala 169:46 27:24]
  wire [31:0] _GEN_1975 = _GEN_722[7:6] == 2'h0 ? tag_3_15 : _GEN_1700; // @[d_cache.scala 169:46 27:24]
  wire  _GEN_1976 = _GEN_722[7:6] == 2'h0 ? valid_3_0 : _GEN_1701; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1977 = _GEN_722[7:6] == 2'h0 ? valid_3_1 : _GEN_1702; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1978 = _GEN_722[7:6] == 2'h0 ? valid_3_2 : _GEN_1703; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1979 = _GEN_722[7:6] == 2'h0 ? valid_3_3 : _GEN_1704; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1980 = _GEN_722[7:6] == 2'h0 ? valid_3_4 : _GEN_1705; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1981 = _GEN_722[7:6] == 2'h0 ? valid_3_5 : _GEN_1706; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1982 = _GEN_722[7:6] == 2'h0 ? valid_3_6 : _GEN_1707; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1983 = _GEN_722[7:6] == 2'h0 ? valid_3_7 : _GEN_1708; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1984 = _GEN_722[7:6] == 2'h0 ? valid_3_8 : _GEN_1709; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1985 = _GEN_722[7:6] == 2'h0 ? valid_3_9 : _GEN_1710; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1986 = _GEN_722[7:6] == 2'h0 ? valid_3_10 : _GEN_1711; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1987 = _GEN_722[7:6] == 2'h0 ? valid_3_11 : _GEN_1712; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1988 = _GEN_722[7:6] == 2'h0 ? valid_3_12 : _GEN_1713; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1989 = _GEN_722[7:6] == 2'h0 ? valid_3_13 : _GEN_1714; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1990 = _GEN_722[7:6] == 2'h0 ? valid_3_14 : _GEN_1715; // @[d_cache.scala 169:46 31:26]
  wire  _GEN_1991 = _GEN_722[7:6] == 2'h0 ? valid_3_15 : _GEN_1716; // @[d_cache.scala 169:46 31:26]
  wire [3:0] _GEN_1992 = unuse_way == 3'h4 ? 4'h1 : _GEN_1735; // @[d_cache.scala 162:40 163:23]
  wire [127:0] _GEN_1993 = unuse_way == 3'h4 ? _GEN_867 : _GEN_1944; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_1994 = unuse_way == 3'h4 ? _GEN_868 : _GEN_1945; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_1995 = unuse_way == 3'h4 ? _GEN_869 : _GEN_1946; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_1996 = unuse_way == 3'h4 ? _GEN_870 : _GEN_1947; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_1997 = unuse_way == 3'h4 ? _GEN_871 : _GEN_1948; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_1998 = unuse_way == 3'h4 ? _GEN_872 : _GEN_1949; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_1999 = unuse_way == 3'h4 ? _GEN_873 : _GEN_1950; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_2000 = unuse_way == 3'h4 ? _GEN_874 : _GEN_1951; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_2001 = unuse_way == 3'h4 ? _GEN_875 : _GEN_1952; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_2002 = unuse_way == 3'h4 ? _GEN_876 : _GEN_1953; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_2003 = unuse_way == 3'h4 ? _GEN_877 : _GEN_1954; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_2004 = unuse_way == 3'h4 ? _GEN_878 : _GEN_1955; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_2005 = unuse_way == 3'h4 ? _GEN_879 : _GEN_1956; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_2006 = unuse_way == 3'h4 ? _GEN_880 : _GEN_1957; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_2007 = unuse_way == 3'h4 ? _GEN_881 : _GEN_1958; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_2008 = unuse_way == 3'h4 ? _GEN_882 : _GEN_1959; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2009 = unuse_way == 3'h4 ? _GEN_883 : _GEN_1960; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2010 = unuse_way == 3'h4 ? _GEN_884 : _GEN_1961; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2011 = unuse_way == 3'h4 ? _GEN_885 : _GEN_1962; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2012 = unuse_way == 3'h4 ? _GEN_886 : _GEN_1963; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2013 = unuse_way == 3'h4 ? _GEN_887 : _GEN_1964; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2014 = unuse_way == 3'h4 ? _GEN_888 : _GEN_1965; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2015 = unuse_way == 3'h4 ? _GEN_889 : _GEN_1966; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2016 = unuse_way == 3'h4 ? _GEN_890 : _GEN_1967; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2017 = unuse_way == 3'h4 ? _GEN_891 : _GEN_1968; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2018 = unuse_way == 3'h4 ? _GEN_892 : _GEN_1969; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2019 = unuse_way == 3'h4 ? _GEN_893 : _GEN_1970; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2020 = unuse_way == 3'h4 ? _GEN_894 : _GEN_1971; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2021 = unuse_way == 3'h4 ? _GEN_895 : _GEN_1972; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2022 = unuse_way == 3'h4 ? _GEN_896 : _GEN_1973; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2023 = unuse_way == 3'h4 ? _GEN_897 : _GEN_1974; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2024 = unuse_way == 3'h4 ? _GEN_898 : _GEN_1975; // @[d_cache.scala 162:40]
  wire  _GEN_2025 = unuse_way == 3'h4 ? _GEN_899 : _GEN_1976; // @[d_cache.scala 162:40]
  wire  _GEN_2026 = unuse_way == 3'h4 ? _GEN_900 : _GEN_1977; // @[d_cache.scala 162:40]
  wire  _GEN_2027 = unuse_way == 3'h4 ? _GEN_901 : _GEN_1978; // @[d_cache.scala 162:40]
  wire  _GEN_2028 = unuse_way == 3'h4 ? _GEN_902 : _GEN_1979; // @[d_cache.scala 162:40]
  wire  _GEN_2029 = unuse_way == 3'h4 ? _GEN_903 : _GEN_1980; // @[d_cache.scala 162:40]
  wire  _GEN_2030 = unuse_way == 3'h4 ? _GEN_904 : _GEN_1981; // @[d_cache.scala 162:40]
  wire  _GEN_2031 = unuse_way == 3'h4 ? _GEN_905 : _GEN_1982; // @[d_cache.scala 162:40]
  wire  _GEN_2032 = unuse_way == 3'h4 ? _GEN_906 : _GEN_1983; // @[d_cache.scala 162:40]
  wire  _GEN_2033 = unuse_way == 3'h4 ? _GEN_907 : _GEN_1984; // @[d_cache.scala 162:40]
  wire  _GEN_2034 = unuse_way == 3'h4 ? _GEN_908 : _GEN_1985; // @[d_cache.scala 162:40]
  wire  _GEN_2035 = unuse_way == 3'h4 ? _GEN_909 : _GEN_1986; // @[d_cache.scala 162:40]
  wire  _GEN_2036 = unuse_way == 3'h4 ? _GEN_910 : _GEN_1987; // @[d_cache.scala 162:40]
  wire  _GEN_2037 = unuse_way == 3'h4 ? _GEN_911 : _GEN_1988; // @[d_cache.scala 162:40]
  wire  _GEN_2038 = unuse_way == 3'h4 ? _GEN_912 : _GEN_1989; // @[d_cache.scala 162:40]
  wire  _GEN_2039 = unuse_way == 3'h4 ? _GEN_913 : _GEN_1990; // @[d_cache.scala 162:40]
  wire  _GEN_2040 = unuse_way == 3'h4 ? _GEN_914 : _GEN_1991; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2041 = unuse_way == 3'h4 ? _GEN_915 : _GEN_1784; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2042 = unuse_way == 3'h4 ? _GEN_916 : _GEN_1785; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2043 = unuse_way == 3'h4 ? _GEN_917 : _GEN_1786; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2044 = unuse_way == 3'h4 ? _GEN_918 : _GEN_1787; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2045 = unuse_way == 3'h4 ? _GEN_919 : _GEN_1788; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2046 = unuse_way == 3'h4 ? _GEN_920 : _GEN_1789; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2047 = unuse_way == 3'h4 ? _GEN_921 : _GEN_1790; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2048 = unuse_way == 3'h4 ? _GEN_922 : _GEN_1791; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2049 = unuse_way == 3'h4 ? _GEN_923 : _GEN_1792; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2050 = unuse_way == 3'h4 ? _GEN_924 : _GEN_1793; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2051 = unuse_way == 3'h4 ? _GEN_925 : _GEN_1794; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2052 = unuse_way == 3'h4 ? _GEN_926 : _GEN_1795; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2053 = unuse_way == 3'h4 ? _GEN_927 : _GEN_1796; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2054 = unuse_way == 3'h4 ? _GEN_928 : _GEN_1797; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2055 = unuse_way == 3'h4 ? _GEN_929 : _GEN_1798; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2056 = unuse_way == 3'h4 ? _GEN_930 : _GEN_1799; // @[d_cache.scala 162:40]
  wire [127:0] _GEN_2057 = unuse_way == 3'h4 ? write_back_data : _GEN_1717; // @[d_cache.scala 162:40 41:34]
  wire [39:0] _GEN_2058 = unuse_way == 3'h4 ? {{8'd0}, write_back_addr} : _GEN_1718; // @[d_cache.scala 162:40 42:34]
  wire  _GEN_2059 = unuse_way == 3'h4 ? dirty_0_0 : _GEN_1719; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2060 = unuse_way == 3'h4 ? dirty_0_1 : _GEN_1720; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2061 = unuse_way == 3'h4 ? dirty_0_2 : _GEN_1721; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2062 = unuse_way == 3'h4 ? dirty_0_3 : _GEN_1722; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2063 = unuse_way == 3'h4 ? dirty_0_4 : _GEN_1723; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2064 = unuse_way == 3'h4 ? dirty_0_5 : _GEN_1724; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2065 = unuse_way == 3'h4 ? dirty_0_6 : _GEN_1725; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2066 = unuse_way == 3'h4 ? dirty_0_7 : _GEN_1726; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2067 = unuse_way == 3'h4 ? dirty_0_8 : _GEN_1727; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2068 = unuse_way == 3'h4 ? dirty_0_9 : _GEN_1728; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2069 = unuse_way == 3'h4 ? dirty_0_10 : _GEN_1729; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2070 = unuse_way == 3'h4 ? dirty_0_11 : _GEN_1730; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2071 = unuse_way == 3'h4 ? dirty_0_12 : _GEN_1731; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2072 = unuse_way == 3'h4 ? dirty_0_13 : _GEN_1732; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2073 = unuse_way == 3'h4 ? dirty_0_14 : _GEN_1733; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2074 = unuse_way == 3'h4 ? dirty_0_15 : _GEN_1734; // @[d_cache.scala 162:40 32:26]
  wire [127:0] _GEN_2075 = unuse_way == 3'h4 ? ram_0_0 : _GEN_1736; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2076 = unuse_way == 3'h4 ? ram_0_1 : _GEN_1737; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2077 = unuse_way == 3'h4 ? ram_0_2 : _GEN_1738; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2078 = unuse_way == 3'h4 ? ram_0_3 : _GEN_1739; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2079 = unuse_way == 3'h4 ? ram_0_4 : _GEN_1740; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2080 = unuse_way == 3'h4 ? ram_0_5 : _GEN_1741; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2081 = unuse_way == 3'h4 ? ram_0_6 : _GEN_1742; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2082 = unuse_way == 3'h4 ? ram_0_7 : _GEN_1743; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2083 = unuse_way == 3'h4 ? ram_0_8 : _GEN_1744; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2084 = unuse_way == 3'h4 ? ram_0_9 : _GEN_1745; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2085 = unuse_way == 3'h4 ? ram_0_10 : _GEN_1746; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2086 = unuse_way == 3'h4 ? ram_0_11 : _GEN_1747; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2087 = unuse_way == 3'h4 ? ram_0_12 : _GEN_1748; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2088 = unuse_way == 3'h4 ? ram_0_13 : _GEN_1749; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2089 = unuse_way == 3'h4 ? ram_0_14 : _GEN_1750; // @[d_cache.scala 162:40 19:24]
  wire [127:0] _GEN_2090 = unuse_way == 3'h4 ? ram_0_15 : _GEN_1751; // @[d_cache.scala 162:40 19:24]
  wire [31:0] _GEN_2091 = unuse_way == 3'h4 ? tag_0_0 : _GEN_1752; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2092 = unuse_way == 3'h4 ? tag_0_1 : _GEN_1753; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2093 = unuse_way == 3'h4 ? tag_0_2 : _GEN_1754; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2094 = unuse_way == 3'h4 ? tag_0_3 : _GEN_1755; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2095 = unuse_way == 3'h4 ? tag_0_4 : _GEN_1756; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2096 = unuse_way == 3'h4 ? tag_0_5 : _GEN_1757; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2097 = unuse_way == 3'h4 ? tag_0_6 : _GEN_1758; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2098 = unuse_way == 3'h4 ? tag_0_7 : _GEN_1759; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2099 = unuse_way == 3'h4 ? tag_0_8 : _GEN_1760; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2100 = unuse_way == 3'h4 ? tag_0_9 : _GEN_1761; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2101 = unuse_way == 3'h4 ? tag_0_10 : _GEN_1762; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2102 = unuse_way == 3'h4 ? tag_0_11 : _GEN_1763; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2103 = unuse_way == 3'h4 ? tag_0_12 : _GEN_1764; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2104 = unuse_way == 3'h4 ? tag_0_13 : _GEN_1765; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2105 = unuse_way == 3'h4 ? tag_0_14 : _GEN_1766; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2106 = unuse_way == 3'h4 ? tag_0_15 : _GEN_1767; // @[d_cache.scala 162:40 24:24]
  wire  _GEN_2107 = unuse_way == 3'h4 ? valid_0_0 : _GEN_1768; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2108 = unuse_way == 3'h4 ? valid_0_1 : _GEN_1769; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2109 = unuse_way == 3'h4 ? valid_0_2 : _GEN_1770; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2110 = unuse_way == 3'h4 ? valid_0_3 : _GEN_1771; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2111 = unuse_way == 3'h4 ? valid_0_4 : _GEN_1772; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2112 = unuse_way == 3'h4 ? valid_0_5 : _GEN_1773; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2113 = unuse_way == 3'h4 ? valid_0_6 : _GEN_1774; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2114 = unuse_way == 3'h4 ? valid_0_7 : _GEN_1775; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2115 = unuse_way == 3'h4 ? valid_0_8 : _GEN_1776; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2116 = unuse_way == 3'h4 ? valid_0_9 : _GEN_1777; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2117 = unuse_way == 3'h4 ? valid_0_10 : _GEN_1778; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2118 = unuse_way == 3'h4 ? valid_0_11 : _GEN_1779; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2119 = unuse_way == 3'h4 ? valid_0_12 : _GEN_1780; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2120 = unuse_way == 3'h4 ? valid_0_13 : _GEN_1781; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2121 = unuse_way == 3'h4 ? valid_0_14 : _GEN_1782; // @[d_cache.scala 162:40 28:26]
  wire  _GEN_2122 = unuse_way == 3'h4 ? valid_0_15 : _GEN_1783; // @[d_cache.scala 162:40 28:26]
  wire [127:0] _GEN_2139 = unuse_way == 3'h4 ? ram_1_0 : _GEN_1816; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2140 = unuse_way == 3'h4 ? ram_1_1 : _GEN_1817; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2141 = unuse_way == 3'h4 ? ram_1_2 : _GEN_1818; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2142 = unuse_way == 3'h4 ? ram_1_3 : _GEN_1819; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2143 = unuse_way == 3'h4 ? ram_1_4 : _GEN_1820; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2144 = unuse_way == 3'h4 ? ram_1_5 : _GEN_1821; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2145 = unuse_way == 3'h4 ? ram_1_6 : _GEN_1822; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2146 = unuse_way == 3'h4 ? ram_1_7 : _GEN_1823; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2147 = unuse_way == 3'h4 ? ram_1_8 : _GEN_1824; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2148 = unuse_way == 3'h4 ? ram_1_9 : _GEN_1825; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2149 = unuse_way == 3'h4 ? ram_1_10 : _GEN_1826; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2150 = unuse_way == 3'h4 ? ram_1_11 : _GEN_1827; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2151 = unuse_way == 3'h4 ? ram_1_12 : _GEN_1828; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2152 = unuse_way == 3'h4 ? ram_1_13 : _GEN_1829; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2153 = unuse_way == 3'h4 ? ram_1_14 : _GEN_1830; // @[d_cache.scala 162:40 20:24]
  wire [127:0] _GEN_2154 = unuse_way == 3'h4 ? ram_1_15 : _GEN_1831; // @[d_cache.scala 162:40 20:24]
  wire [31:0] _GEN_2155 = unuse_way == 3'h4 ? tag_1_0 : _GEN_1832; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2156 = unuse_way == 3'h4 ? tag_1_1 : _GEN_1833; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2157 = unuse_way == 3'h4 ? tag_1_2 : _GEN_1834; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2158 = unuse_way == 3'h4 ? tag_1_3 : _GEN_1835; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2159 = unuse_way == 3'h4 ? tag_1_4 : _GEN_1836; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2160 = unuse_way == 3'h4 ? tag_1_5 : _GEN_1837; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2161 = unuse_way == 3'h4 ? tag_1_6 : _GEN_1838; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2162 = unuse_way == 3'h4 ? tag_1_7 : _GEN_1839; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2163 = unuse_way == 3'h4 ? tag_1_8 : _GEN_1840; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2164 = unuse_way == 3'h4 ? tag_1_9 : _GEN_1841; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2165 = unuse_way == 3'h4 ? tag_1_10 : _GEN_1842; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2166 = unuse_way == 3'h4 ? tag_1_11 : _GEN_1843; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2167 = unuse_way == 3'h4 ? tag_1_12 : _GEN_1844; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2168 = unuse_way == 3'h4 ? tag_1_13 : _GEN_1845; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2169 = unuse_way == 3'h4 ? tag_1_14 : _GEN_1846; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_2170 = unuse_way == 3'h4 ? tag_1_15 : _GEN_1847; // @[d_cache.scala 162:40 25:24]
  wire  _GEN_2171 = unuse_way == 3'h4 ? valid_1_0 : _GEN_1848; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2172 = unuse_way == 3'h4 ? valid_1_1 : _GEN_1849; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2173 = unuse_way == 3'h4 ? valid_1_2 : _GEN_1850; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2174 = unuse_way == 3'h4 ? valid_1_3 : _GEN_1851; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2175 = unuse_way == 3'h4 ? valid_1_4 : _GEN_1852; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2176 = unuse_way == 3'h4 ? valid_1_5 : _GEN_1853; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2177 = unuse_way == 3'h4 ? valid_1_6 : _GEN_1854; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2178 = unuse_way == 3'h4 ? valid_1_7 : _GEN_1855; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2179 = unuse_way == 3'h4 ? valid_1_8 : _GEN_1856; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2180 = unuse_way == 3'h4 ? valid_1_9 : _GEN_1857; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2181 = unuse_way == 3'h4 ? valid_1_10 : _GEN_1858; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2182 = unuse_way == 3'h4 ? valid_1_11 : _GEN_1859; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2183 = unuse_way == 3'h4 ? valid_1_12 : _GEN_1860; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2184 = unuse_way == 3'h4 ? valid_1_13 : _GEN_1861; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2185 = unuse_way == 3'h4 ? valid_1_14 : _GEN_1862; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2186 = unuse_way == 3'h4 ? valid_1_15 : _GEN_1863; // @[d_cache.scala 162:40 29:26]
  wire [127:0] _GEN_2203 = unuse_way == 3'h4 ? ram_2_0 : _GEN_1880; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2204 = unuse_way == 3'h4 ? ram_2_1 : _GEN_1881; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2205 = unuse_way == 3'h4 ? ram_2_2 : _GEN_1882; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2206 = unuse_way == 3'h4 ? ram_2_3 : _GEN_1883; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2207 = unuse_way == 3'h4 ? ram_2_4 : _GEN_1884; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2208 = unuse_way == 3'h4 ? ram_2_5 : _GEN_1885; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2209 = unuse_way == 3'h4 ? ram_2_6 : _GEN_1886; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2210 = unuse_way == 3'h4 ? ram_2_7 : _GEN_1887; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2211 = unuse_way == 3'h4 ? ram_2_8 : _GEN_1888; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2212 = unuse_way == 3'h4 ? ram_2_9 : _GEN_1889; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2213 = unuse_way == 3'h4 ? ram_2_10 : _GEN_1890; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2214 = unuse_way == 3'h4 ? ram_2_11 : _GEN_1891; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2215 = unuse_way == 3'h4 ? ram_2_12 : _GEN_1892; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2216 = unuse_way == 3'h4 ? ram_2_13 : _GEN_1893; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2217 = unuse_way == 3'h4 ? ram_2_14 : _GEN_1894; // @[d_cache.scala 162:40 21:24]
  wire [127:0] _GEN_2218 = unuse_way == 3'h4 ? ram_2_15 : _GEN_1895; // @[d_cache.scala 162:40 21:24]
  wire [31:0] _GEN_2219 = unuse_way == 3'h4 ? tag_2_0 : _GEN_1896; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2220 = unuse_way == 3'h4 ? tag_2_1 : _GEN_1897; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2221 = unuse_way == 3'h4 ? tag_2_2 : _GEN_1898; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2222 = unuse_way == 3'h4 ? tag_2_3 : _GEN_1899; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2223 = unuse_way == 3'h4 ? tag_2_4 : _GEN_1900; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2224 = unuse_way == 3'h4 ? tag_2_5 : _GEN_1901; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2225 = unuse_way == 3'h4 ? tag_2_6 : _GEN_1902; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2226 = unuse_way == 3'h4 ? tag_2_7 : _GEN_1903; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2227 = unuse_way == 3'h4 ? tag_2_8 : _GEN_1904; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2228 = unuse_way == 3'h4 ? tag_2_9 : _GEN_1905; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2229 = unuse_way == 3'h4 ? tag_2_10 : _GEN_1906; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2230 = unuse_way == 3'h4 ? tag_2_11 : _GEN_1907; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2231 = unuse_way == 3'h4 ? tag_2_12 : _GEN_1908; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2232 = unuse_way == 3'h4 ? tag_2_13 : _GEN_1909; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2233 = unuse_way == 3'h4 ? tag_2_14 : _GEN_1910; // @[d_cache.scala 162:40 26:24]
  wire [31:0] _GEN_2234 = unuse_way == 3'h4 ? tag_2_15 : _GEN_1911; // @[d_cache.scala 162:40 26:24]
  wire  _GEN_2235 = unuse_way == 3'h4 ? valid_2_0 : _GEN_1912; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2236 = unuse_way == 3'h4 ? valid_2_1 : _GEN_1913; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2237 = unuse_way == 3'h4 ? valid_2_2 : _GEN_1914; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2238 = unuse_way == 3'h4 ? valid_2_3 : _GEN_1915; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2239 = unuse_way == 3'h4 ? valid_2_4 : _GEN_1916; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2240 = unuse_way == 3'h4 ? valid_2_5 : _GEN_1917; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2241 = unuse_way == 3'h4 ? valid_2_6 : _GEN_1918; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2242 = unuse_way == 3'h4 ? valid_2_7 : _GEN_1919; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2243 = unuse_way == 3'h4 ? valid_2_8 : _GEN_1920; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2244 = unuse_way == 3'h4 ? valid_2_9 : _GEN_1921; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2245 = unuse_way == 3'h4 ? valid_2_10 : _GEN_1922; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2246 = unuse_way == 3'h4 ? valid_2_11 : _GEN_1923; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2247 = unuse_way == 3'h4 ? valid_2_12 : _GEN_1924; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2248 = unuse_way == 3'h4 ? valid_2_13 : _GEN_1925; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2249 = unuse_way == 3'h4 ? valid_2_14 : _GEN_1926; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2250 = unuse_way == 3'h4 ? valid_2_15 : _GEN_1927; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_2251 = unuse_way == 3'h4 ? dirty_3_0 : _GEN_1928; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2252 = unuse_way == 3'h4 ? dirty_3_1 : _GEN_1929; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2253 = unuse_way == 3'h4 ? dirty_3_2 : _GEN_1930; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2254 = unuse_way == 3'h4 ? dirty_3_3 : _GEN_1931; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2255 = unuse_way == 3'h4 ? dirty_3_4 : _GEN_1932; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2256 = unuse_way == 3'h4 ? dirty_3_5 : _GEN_1933; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2257 = unuse_way == 3'h4 ? dirty_3_6 : _GEN_1934; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2258 = unuse_way == 3'h4 ? dirty_3_7 : _GEN_1935; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2259 = unuse_way == 3'h4 ? dirty_3_8 : _GEN_1936; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2260 = unuse_way == 3'h4 ? dirty_3_9 : _GEN_1937; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2261 = unuse_way == 3'h4 ? dirty_3_10 : _GEN_1938; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2262 = unuse_way == 3'h4 ? dirty_3_11 : _GEN_1939; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2263 = unuse_way == 3'h4 ? dirty_3_12 : _GEN_1940; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2264 = unuse_way == 3'h4 ? dirty_3_13 : _GEN_1941; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2265 = unuse_way == 3'h4 ? dirty_3_14 : _GEN_1942; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_2266 = unuse_way == 3'h4 ? dirty_3_15 : _GEN_1943; // @[d_cache.scala 162:40 35:26]
  wire [3:0] _GEN_2267 = unuse_way == 3'h3 ? 4'h1 : _GEN_1992; // @[d_cache.scala 156:40 157:23]
  wire [127:0] _GEN_2268 = unuse_way == 3'h3 ? _GEN_803 : _GEN_2203; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2269 = unuse_way == 3'h3 ? _GEN_804 : _GEN_2204; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2270 = unuse_way == 3'h3 ? _GEN_805 : _GEN_2205; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2271 = unuse_way == 3'h3 ? _GEN_806 : _GEN_2206; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2272 = unuse_way == 3'h3 ? _GEN_807 : _GEN_2207; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2273 = unuse_way == 3'h3 ? _GEN_808 : _GEN_2208; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2274 = unuse_way == 3'h3 ? _GEN_809 : _GEN_2209; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2275 = unuse_way == 3'h3 ? _GEN_810 : _GEN_2210; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2276 = unuse_way == 3'h3 ? _GEN_811 : _GEN_2211; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2277 = unuse_way == 3'h3 ? _GEN_812 : _GEN_2212; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2278 = unuse_way == 3'h3 ? _GEN_813 : _GEN_2213; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2279 = unuse_way == 3'h3 ? _GEN_814 : _GEN_2214; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2280 = unuse_way == 3'h3 ? _GEN_815 : _GEN_2215; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2281 = unuse_way == 3'h3 ? _GEN_816 : _GEN_2216; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2282 = unuse_way == 3'h3 ? _GEN_817 : _GEN_2217; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2283 = unuse_way == 3'h3 ? _GEN_818 : _GEN_2218; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2284 = unuse_way == 3'h3 ? _GEN_819 : _GEN_2219; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2285 = unuse_way == 3'h3 ? _GEN_820 : _GEN_2220; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2286 = unuse_way == 3'h3 ? _GEN_821 : _GEN_2221; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2287 = unuse_way == 3'h3 ? _GEN_822 : _GEN_2222; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2288 = unuse_way == 3'h3 ? _GEN_823 : _GEN_2223; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2289 = unuse_way == 3'h3 ? _GEN_824 : _GEN_2224; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2290 = unuse_way == 3'h3 ? _GEN_825 : _GEN_2225; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2291 = unuse_way == 3'h3 ? _GEN_826 : _GEN_2226; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2292 = unuse_way == 3'h3 ? _GEN_827 : _GEN_2227; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2293 = unuse_way == 3'h3 ? _GEN_828 : _GEN_2228; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2294 = unuse_way == 3'h3 ? _GEN_829 : _GEN_2229; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2295 = unuse_way == 3'h3 ? _GEN_830 : _GEN_2230; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2296 = unuse_way == 3'h3 ? _GEN_831 : _GEN_2231; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2297 = unuse_way == 3'h3 ? _GEN_832 : _GEN_2232; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2298 = unuse_way == 3'h3 ? _GEN_833 : _GEN_2233; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_2299 = unuse_way == 3'h3 ? _GEN_834 : _GEN_2234; // @[d_cache.scala 156:40]
  wire  _GEN_2300 = unuse_way == 3'h3 ? _GEN_835 : _GEN_2235; // @[d_cache.scala 156:40]
  wire  _GEN_2301 = unuse_way == 3'h3 ? _GEN_836 : _GEN_2236; // @[d_cache.scala 156:40]
  wire  _GEN_2302 = unuse_way == 3'h3 ? _GEN_837 : _GEN_2237; // @[d_cache.scala 156:40]
  wire  _GEN_2303 = unuse_way == 3'h3 ? _GEN_838 : _GEN_2238; // @[d_cache.scala 156:40]
  wire  _GEN_2304 = unuse_way == 3'h3 ? _GEN_839 : _GEN_2239; // @[d_cache.scala 156:40]
  wire  _GEN_2305 = unuse_way == 3'h3 ? _GEN_840 : _GEN_2240; // @[d_cache.scala 156:40]
  wire  _GEN_2306 = unuse_way == 3'h3 ? _GEN_841 : _GEN_2241; // @[d_cache.scala 156:40]
  wire  _GEN_2307 = unuse_way == 3'h3 ? _GEN_842 : _GEN_2242; // @[d_cache.scala 156:40]
  wire  _GEN_2308 = unuse_way == 3'h3 ? _GEN_843 : _GEN_2243; // @[d_cache.scala 156:40]
  wire  _GEN_2309 = unuse_way == 3'h3 ? _GEN_844 : _GEN_2244; // @[d_cache.scala 156:40]
  wire  _GEN_2310 = unuse_way == 3'h3 ? _GEN_845 : _GEN_2245; // @[d_cache.scala 156:40]
  wire  _GEN_2311 = unuse_way == 3'h3 ? _GEN_846 : _GEN_2246; // @[d_cache.scala 156:40]
  wire  _GEN_2312 = unuse_way == 3'h3 ? _GEN_847 : _GEN_2247; // @[d_cache.scala 156:40]
  wire  _GEN_2313 = unuse_way == 3'h3 ? _GEN_848 : _GEN_2248; // @[d_cache.scala 156:40]
  wire  _GEN_2314 = unuse_way == 3'h3 ? _GEN_849 : _GEN_2249; // @[d_cache.scala 156:40]
  wire  _GEN_2315 = unuse_way == 3'h3 ? _GEN_850 : _GEN_2250; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2316 = unuse_way == 3'h3 ? _GEN_851 : _GEN_2041; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2317 = unuse_way == 3'h3 ? _GEN_852 : _GEN_2042; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2318 = unuse_way == 3'h3 ? _GEN_853 : _GEN_2043; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2319 = unuse_way == 3'h3 ? _GEN_854 : _GEN_2044; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2320 = unuse_way == 3'h3 ? _GEN_855 : _GEN_2045; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2321 = unuse_way == 3'h3 ? _GEN_856 : _GEN_2046; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2322 = unuse_way == 3'h3 ? _GEN_857 : _GEN_2047; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2323 = unuse_way == 3'h3 ? _GEN_858 : _GEN_2048; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2324 = unuse_way == 3'h3 ? _GEN_859 : _GEN_2049; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2325 = unuse_way == 3'h3 ? _GEN_860 : _GEN_2050; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2326 = unuse_way == 3'h3 ? _GEN_861 : _GEN_2051; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2327 = unuse_way == 3'h3 ? _GEN_862 : _GEN_2052; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2328 = unuse_way == 3'h3 ? _GEN_863 : _GEN_2053; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2329 = unuse_way == 3'h3 ? _GEN_864 : _GEN_2054; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2330 = unuse_way == 3'h3 ? _GEN_865 : _GEN_2055; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_2331 = unuse_way == 3'h3 ? _GEN_866 : _GEN_2056; // @[d_cache.scala 156:40]
  wire [127:0] _GEN_2332 = unuse_way == 3'h3 ? ram_3_0 : _GEN_1993; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2333 = unuse_way == 3'h3 ? ram_3_1 : _GEN_1994; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2334 = unuse_way == 3'h3 ? ram_3_2 : _GEN_1995; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2335 = unuse_way == 3'h3 ? ram_3_3 : _GEN_1996; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2336 = unuse_way == 3'h3 ? ram_3_4 : _GEN_1997; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2337 = unuse_way == 3'h3 ? ram_3_5 : _GEN_1998; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2338 = unuse_way == 3'h3 ? ram_3_6 : _GEN_1999; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2339 = unuse_way == 3'h3 ? ram_3_7 : _GEN_2000; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2340 = unuse_way == 3'h3 ? ram_3_8 : _GEN_2001; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2341 = unuse_way == 3'h3 ? ram_3_9 : _GEN_2002; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2342 = unuse_way == 3'h3 ? ram_3_10 : _GEN_2003; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2343 = unuse_way == 3'h3 ? ram_3_11 : _GEN_2004; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2344 = unuse_way == 3'h3 ? ram_3_12 : _GEN_2005; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2345 = unuse_way == 3'h3 ? ram_3_13 : _GEN_2006; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2346 = unuse_way == 3'h3 ? ram_3_14 : _GEN_2007; // @[d_cache.scala 156:40 22:24]
  wire [127:0] _GEN_2347 = unuse_way == 3'h3 ? ram_3_15 : _GEN_2008; // @[d_cache.scala 156:40 22:24]
  wire [31:0] _GEN_2348 = unuse_way == 3'h3 ? tag_3_0 : _GEN_2009; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2349 = unuse_way == 3'h3 ? tag_3_1 : _GEN_2010; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2350 = unuse_way == 3'h3 ? tag_3_2 : _GEN_2011; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2351 = unuse_way == 3'h3 ? tag_3_3 : _GEN_2012; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2352 = unuse_way == 3'h3 ? tag_3_4 : _GEN_2013; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2353 = unuse_way == 3'h3 ? tag_3_5 : _GEN_2014; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2354 = unuse_way == 3'h3 ? tag_3_6 : _GEN_2015; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2355 = unuse_way == 3'h3 ? tag_3_7 : _GEN_2016; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2356 = unuse_way == 3'h3 ? tag_3_8 : _GEN_2017; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2357 = unuse_way == 3'h3 ? tag_3_9 : _GEN_2018; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2358 = unuse_way == 3'h3 ? tag_3_10 : _GEN_2019; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2359 = unuse_way == 3'h3 ? tag_3_11 : _GEN_2020; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2360 = unuse_way == 3'h3 ? tag_3_12 : _GEN_2021; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2361 = unuse_way == 3'h3 ? tag_3_13 : _GEN_2022; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2362 = unuse_way == 3'h3 ? tag_3_14 : _GEN_2023; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_2363 = unuse_way == 3'h3 ? tag_3_15 : _GEN_2024; // @[d_cache.scala 156:40 27:24]
  wire  _GEN_2364 = unuse_way == 3'h3 ? valid_3_0 : _GEN_2025; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2365 = unuse_way == 3'h3 ? valid_3_1 : _GEN_2026; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2366 = unuse_way == 3'h3 ? valid_3_2 : _GEN_2027; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2367 = unuse_way == 3'h3 ? valid_3_3 : _GEN_2028; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2368 = unuse_way == 3'h3 ? valid_3_4 : _GEN_2029; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2369 = unuse_way == 3'h3 ? valid_3_5 : _GEN_2030; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2370 = unuse_way == 3'h3 ? valid_3_6 : _GEN_2031; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2371 = unuse_way == 3'h3 ? valid_3_7 : _GEN_2032; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2372 = unuse_way == 3'h3 ? valid_3_8 : _GEN_2033; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2373 = unuse_way == 3'h3 ? valid_3_9 : _GEN_2034; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2374 = unuse_way == 3'h3 ? valid_3_10 : _GEN_2035; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2375 = unuse_way == 3'h3 ? valid_3_11 : _GEN_2036; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2376 = unuse_way == 3'h3 ? valid_3_12 : _GEN_2037; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2377 = unuse_way == 3'h3 ? valid_3_13 : _GEN_2038; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2378 = unuse_way == 3'h3 ? valid_3_14 : _GEN_2039; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_2379 = unuse_way == 3'h3 ? valid_3_15 : _GEN_2040; // @[d_cache.scala 156:40 31:26]
  wire [127:0] _GEN_2380 = unuse_way == 3'h3 ? write_back_data : _GEN_2057; // @[d_cache.scala 156:40 41:34]
  wire [39:0] _GEN_2381 = unuse_way == 3'h3 ? {{8'd0}, write_back_addr} : _GEN_2058; // @[d_cache.scala 156:40 42:34]
  wire  _GEN_2382 = unuse_way == 3'h3 ? dirty_0_0 : _GEN_2059; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2383 = unuse_way == 3'h3 ? dirty_0_1 : _GEN_2060; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2384 = unuse_way == 3'h3 ? dirty_0_2 : _GEN_2061; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2385 = unuse_way == 3'h3 ? dirty_0_3 : _GEN_2062; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2386 = unuse_way == 3'h3 ? dirty_0_4 : _GEN_2063; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2387 = unuse_way == 3'h3 ? dirty_0_5 : _GEN_2064; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2388 = unuse_way == 3'h3 ? dirty_0_6 : _GEN_2065; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2389 = unuse_way == 3'h3 ? dirty_0_7 : _GEN_2066; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2390 = unuse_way == 3'h3 ? dirty_0_8 : _GEN_2067; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2391 = unuse_way == 3'h3 ? dirty_0_9 : _GEN_2068; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2392 = unuse_way == 3'h3 ? dirty_0_10 : _GEN_2069; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2393 = unuse_way == 3'h3 ? dirty_0_11 : _GEN_2070; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2394 = unuse_way == 3'h3 ? dirty_0_12 : _GEN_2071; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2395 = unuse_way == 3'h3 ? dirty_0_13 : _GEN_2072; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2396 = unuse_way == 3'h3 ? dirty_0_14 : _GEN_2073; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_2397 = unuse_way == 3'h3 ? dirty_0_15 : _GEN_2074; // @[d_cache.scala 156:40 32:26]
  wire [127:0] _GEN_2398 = unuse_way == 3'h3 ? ram_0_0 : _GEN_2075; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2399 = unuse_way == 3'h3 ? ram_0_1 : _GEN_2076; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2400 = unuse_way == 3'h3 ? ram_0_2 : _GEN_2077; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2401 = unuse_way == 3'h3 ? ram_0_3 : _GEN_2078; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2402 = unuse_way == 3'h3 ? ram_0_4 : _GEN_2079; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2403 = unuse_way == 3'h3 ? ram_0_5 : _GEN_2080; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2404 = unuse_way == 3'h3 ? ram_0_6 : _GEN_2081; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2405 = unuse_way == 3'h3 ? ram_0_7 : _GEN_2082; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2406 = unuse_way == 3'h3 ? ram_0_8 : _GEN_2083; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2407 = unuse_way == 3'h3 ? ram_0_9 : _GEN_2084; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2408 = unuse_way == 3'h3 ? ram_0_10 : _GEN_2085; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2409 = unuse_way == 3'h3 ? ram_0_11 : _GEN_2086; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2410 = unuse_way == 3'h3 ? ram_0_12 : _GEN_2087; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2411 = unuse_way == 3'h3 ? ram_0_13 : _GEN_2088; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2412 = unuse_way == 3'h3 ? ram_0_14 : _GEN_2089; // @[d_cache.scala 156:40 19:24]
  wire [127:0] _GEN_2413 = unuse_way == 3'h3 ? ram_0_15 : _GEN_2090; // @[d_cache.scala 156:40 19:24]
  wire [31:0] _GEN_2414 = unuse_way == 3'h3 ? tag_0_0 : _GEN_2091; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2415 = unuse_way == 3'h3 ? tag_0_1 : _GEN_2092; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2416 = unuse_way == 3'h3 ? tag_0_2 : _GEN_2093; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2417 = unuse_way == 3'h3 ? tag_0_3 : _GEN_2094; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2418 = unuse_way == 3'h3 ? tag_0_4 : _GEN_2095; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2419 = unuse_way == 3'h3 ? tag_0_5 : _GEN_2096; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2420 = unuse_way == 3'h3 ? tag_0_6 : _GEN_2097; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2421 = unuse_way == 3'h3 ? tag_0_7 : _GEN_2098; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2422 = unuse_way == 3'h3 ? tag_0_8 : _GEN_2099; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2423 = unuse_way == 3'h3 ? tag_0_9 : _GEN_2100; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2424 = unuse_way == 3'h3 ? tag_0_10 : _GEN_2101; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2425 = unuse_way == 3'h3 ? tag_0_11 : _GEN_2102; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2426 = unuse_way == 3'h3 ? tag_0_12 : _GEN_2103; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2427 = unuse_way == 3'h3 ? tag_0_13 : _GEN_2104; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2428 = unuse_way == 3'h3 ? tag_0_14 : _GEN_2105; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_2429 = unuse_way == 3'h3 ? tag_0_15 : _GEN_2106; // @[d_cache.scala 156:40 24:24]
  wire  _GEN_2430 = unuse_way == 3'h3 ? valid_0_0 : _GEN_2107; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2431 = unuse_way == 3'h3 ? valid_0_1 : _GEN_2108; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2432 = unuse_way == 3'h3 ? valid_0_2 : _GEN_2109; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2433 = unuse_way == 3'h3 ? valid_0_3 : _GEN_2110; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2434 = unuse_way == 3'h3 ? valid_0_4 : _GEN_2111; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2435 = unuse_way == 3'h3 ? valid_0_5 : _GEN_2112; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2436 = unuse_way == 3'h3 ? valid_0_6 : _GEN_2113; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2437 = unuse_way == 3'h3 ? valid_0_7 : _GEN_2114; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2438 = unuse_way == 3'h3 ? valid_0_8 : _GEN_2115; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2439 = unuse_way == 3'h3 ? valid_0_9 : _GEN_2116; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2440 = unuse_way == 3'h3 ? valid_0_10 : _GEN_2117; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2441 = unuse_way == 3'h3 ? valid_0_11 : _GEN_2118; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2442 = unuse_way == 3'h3 ? valid_0_12 : _GEN_2119; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2443 = unuse_way == 3'h3 ? valid_0_13 : _GEN_2120; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2444 = unuse_way == 3'h3 ? valid_0_14 : _GEN_2121; // @[d_cache.scala 156:40 28:26]
  wire  _GEN_2445 = unuse_way == 3'h3 ? valid_0_15 : _GEN_2122; // @[d_cache.scala 156:40 28:26]
  wire [127:0] _GEN_2462 = unuse_way == 3'h3 ? ram_1_0 : _GEN_2139; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2463 = unuse_way == 3'h3 ? ram_1_1 : _GEN_2140; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2464 = unuse_way == 3'h3 ? ram_1_2 : _GEN_2141; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2465 = unuse_way == 3'h3 ? ram_1_3 : _GEN_2142; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2466 = unuse_way == 3'h3 ? ram_1_4 : _GEN_2143; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2467 = unuse_way == 3'h3 ? ram_1_5 : _GEN_2144; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2468 = unuse_way == 3'h3 ? ram_1_6 : _GEN_2145; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2469 = unuse_way == 3'h3 ? ram_1_7 : _GEN_2146; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2470 = unuse_way == 3'h3 ? ram_1_8 : _GEN_2147; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2471 = unuse_way == 3'h3 ? ram_1_9 : _GEN_2148; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2472 = unuse_way == 3'h3 ? ram_1_10 : _GEN_2149; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2473 = unuse_way == 3'h3 ? ram_1_11 : _GEN_2150; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2474 = unuse_way == 3'h3 ? ram_1_12 : _GEN_2151; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2475 = unuse_way == 3'h3 ? ram_1_13 : _GEN_2152; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2476 = unuse_way == 3'h3 ? ram_1_14 : _GEN_2153; // @[d_cache.scala 156:40 20:24]
  wire [127:0] _GEN_2477 = unuse_way == 3'h3 ? ram_1_15 : _GEN_2154; // @[d_cache.scala 156:40 20:24]
  wire [31:0] _GEN_2478 = unuse_way == 3'h3 ? tag_1_0 : _GEN_2155; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2479 = unuse_way == 3'h3 ? tag_1_1 : _GEN_2156; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2480 = unuse_way == 3'h3 ? tag_1_2 : _GEN_2157; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2481 = unuse_way == 3'h3 ? tag_1_3 : _GEN_2158; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2482 = unuse_way == 3'h3 ? tag_1_4 : _GEN_2159; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2483 = unuse_way == 3'h3 ? tag_1_5 : _GEN_2160; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2484 = unuse_way == 3'h3 ? tag_1_6 : _GEN_2161; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2485 = unuse_way == 3'h3 ? tag_1_7 : _GEN_2162; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2486 = unuse_way == 3'h3 ? tag_1_8 : _GEN_2163; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2487 = unuse_way == 3'h3 ? tag_1_9 : _GEN_2164; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2488 = unuse_way == 3'h3 ? tag_1_10 : _GEN_2165; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2489 = unuse_way == 3'h3 ? tag_1_11 : _GEN_2166; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2490 = unuse_way == 3'h3 ? tag_1_12 : _GEN_2167; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2491 = unuse_way == 3'h3 ? tag_1_13 : _GEN_2168; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2492 = unuse_way == 3'h3 ? tag_1_14 : _GEN_2169; // @[d_cache.scala 156:40 25:24]
  wire [31:0] _GEN_2493 = unuse_way == 3'h3 ? tag_1_15 : _GEN_2170; // @[d_cache.scala 156:40 25:24]
  wire  _GEN_2494 = unuse_way == 3'h3 ? valid_1_0 : _GEN_2171; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2495 = unuse_way == 3'h3 ? valid_1_1 : _GEN_2172; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2496 = unuse_way == 3'h3 ? valid_1_2 : _GEN_2173; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2497 = unuse_way == 3'h3 ? valid_1_3 : _GEN_2174; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2498 = unuse_way == 3'h3 ? valid_1_4 : _GEN_2175; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2499 = unuse_way == 3'h3 ? valid_1_5 : _GEN_2176; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2500 = unuse_way == 3'h3 ? valid_1_6 : _GEN_2177; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2501 = unuse_way == 3'h3 ? valid_1_7 : _GEN_2178; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2502 = unuse_way == 3'h3 ? valid_1_8 : _GEN_2179; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2503 = unuse_way == 3'h3 ? valid_1_9 : _GEN_2180; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2504 = unuse_way == 3'h3 ? valid_1_10 : _GEN_2181; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2505 = unuse_way == 3'h3 ? valid_1_11 : _GEN_2182; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2506 = unuse_way == 3'h3 ? valid_1_12 : _GEN_2183; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2507 = unuse_way == 3'h3 ? valid_1_13 : _GEN_2184; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2508 = unuse_way == 3'h3 ? valid_1_14 : _GEN_2185; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2509 = unuse_way == 3'h3 ? valid_1_15 : _GEN_2186; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_2526 = unuse_way == 3'h3 ? dirty_3_0 : _GEN_2251; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2527 = unuse_way == 3'h3 ? dirty_3_1 : _GEN_2252; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2528 = unuse_way == 3'h3 ? dirty_3_2 : _GEN_2253; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2529 = unuse_way == 3'h3 ? dirty_3_3 : _GEN_2254; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2530 = unuse_way == 3'h3 ? dirty_3_4 : _GEN_2255; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2531 = unuse_way == 3'h3 ? dirty_3_5 : _GEN_2256; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2532 = unuse_way == 3'h3 ? dirty_3_6 : _GEN_2257; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2533 = unuse_way == 3'h3 ? dirty_3_7 : _GEN_2258; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2534 = unuse_way == 3'h3 ? dirty_3_8 : _GEN_2259; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2535 = unuse_way == 3'h3 ? dirty_3_9 : _GEN_2260; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2536 = unuse_way == 3'h3 ? dirty_3_10 : _GEN_2261; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2537 = unuse_way == 3'h3 ? dirty_3_11 : _GEN_2262; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2538 = unuse_way == 3'h3 ? dirty_3_12 : _GEN_2263; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2539 = unuse_way == 3'h3 ? dirty_3_13 : _GEN_2264; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2540 = unuse_way == 3'h3 ? dirty_3_14 : _GEN_2265; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_2541 = unuse_way == 3'h3 ? dirty_3_15 : _GEN_2266; // @[d_cache.scala 156:40 35:26]
  wire [3:0] _GEN_2542 = unuse_way == 3'h2 ? 4'h1 : _GEN_2267; // @[d_cache.scala 150:40 151:23]
  wire [127:0] _GEN_2543 = unuse_way == 3'h2 ? _GEN_739 : _GEN_2462; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2544 = unuse_way == 3'h2 ? _GEN_740 : _GEN_2463; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2545 = unuse_way == 3'h2 ? _GEN_741 : _GEN_2464; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2546 = unuse_way == 3'h2 ? _GEN_742 : _GEN_2465; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2547 = unuse_way == 3'h2 ? _GEN_743 : _GEN_2466; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2548 = unuse_way == 3'h2 ? _GEN_744 : _GEN_2467; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2549 = unuse_way == 3'h2 ? _GEN_745 : _GEN_2468; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2550 = unuse_way == 3'h2 ? _GEN_746 : _GEN_2469; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2551 = unuse_way == 3'h2 ? _GEN_747 : _GEN_2470; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2552 = unuse_way == 3'h2 ? _GEN_748 : _GEN_2471; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2553 = unuse_way == 3'h2 ? _GEN_749 : _GEN_2472; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2554 = unuse_way == 3'h2 ? _GEN_750 : _GEN_2473; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2555 = unuse_way == 3'h2 ? _GEN_751 : _GEN_2474; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2556 = unuse_way == 3'h2 ? _GEN_752 : _GEN_2475; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2557 = unuse_way == 3'h2 ? _GEN_753 : _GEN_2476; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2558 = unuse_way == 3'h2 ? _GEN_754 : _GEN_2477; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2559 = unuse_way == 3'h2 ? _GEN_755 : _GEN_2478; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2560 = unuse_way == 3'h2 ? _GEN_756 : _GEN_2479; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2561 = unuse_way == 3'h2 ? _GEN_757 : _GEN_2480; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2562 = unuse_way == 3'h2 ? _GEN_758 : _GEN_2481; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2563 = unuse_way == 3'h2 ? _GEN_759 : _GEN_2482; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2564 = unuse_way == 3'h2 ? _GEN_760 : _GEN_2483; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2565 = unuse_way == 3'h2 ? _GEN_761 : _GEN_2484; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2566 = unuse_way == 3'h2 ? _GEN_762 : _GEN_2485; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2567 = unuse_way == 3'h2 ? _GEN_763 : _GEN_2486; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2568 = unuse_way == 3'h2 ? _GEN_764 : _GEN_2487; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2569 = unuse_way == 3'h2 ? _GEN_765 : _GEN_2488; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2570 = unuse_way == 3'h2 ? _GEN_766 : _GEN_2489; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2571 = unuse_way == 3'h2 ? _GEN_767 : _GEN_2490; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2572 = unuse_way == 3'h2 ? _GEN_768 : _GEN_2491; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2573 = unuse_way == 3'h2 ? _GEN_769 : _GEN_2492; // @[d_cache.scala 150:40]
  wire [31:0] _GEN_2574 = unuse_way == 3'h2 ? _GEN_770 : _GEN_2493; // @[d_cache.scala 150:40]
  wire  _GEN_2575 = unuse_way == 3'h2 ? _GEN_771 : _GEN_2494; // @[d_cache.scala 150:40]
  wire  _GEN_2576 = unuse_way == 3'h2 ? _GEN_772 : _GEN_2495; // @[d_cache.scala 150:40]
  wire  _GEN_2577 = unuse_way == 3'h2 ? _GEN_773 : _GEN_2496; // @[d_cache.scala 150:40]
  wire  _GEN_2578 = unuse_way == 3'h2 ? _GEN_774 : _GEN_2497; // @[d_cache.scala 150:40]
  wire  _GEN_2579 = unuse_way == 3'h2 ? _GEN_775 : _GEN_2498; // @[d_cache.scala 150:40]
  wire  _GEN_2580 = unuse_way == 3'h2 ? _GEN_776 : _GEN_2499; // @[d_cache.scala 150:40]
  wire  _GEN_2581 = unuse_way == 3'h2 ? _GEN_777 : _GEN_2500; // @[d_cache.scala 150:40]
  wire  _GEN_2582 = unuse_way == 3'h2 ? _GEN_778 : _GEN_2501; // @[d_cache.scala 150:40]
  wire  _GEN_2583 = unuse_way == 3'h2 ? _GEN_779 : _GEN_2502; // @[d_cache.scala 150:40]
  wire  _GEN_2584 = unuse_way == 3'h2 ? _GEN_780 : _GEN_2503; // @[d_cache.scala 150:40]
  wire  _GEN_2585 = unuse_way == 3'h2 ? _GEN_781 : _GEN_2504; // @[d_cache.scala 150:40]
  wire  _GEN_2586 = unuse_way == 3'h2 ? _GEN_782 : _GEN_2505; // @[d_cache.scala 150:40]
  wire  _GEN_2587 = unuse_way == 3'h2 ? _GEN_783 : _GEN_2506; // @[d_cache.scala 150:40]
  wire  _GEN_2588 = unuse_way == 3'h2 ? _GEN_784 : _GEN_2507; // @[d_cache.scala 150:40]
  wire  _GEN_2589 = unuse_way == 3'h2 ? _GEN_785 : _GEN_2508; // @[d_cache.scala 150:40]
  wire  _GEN_2590 = unuse_way == 3'h2 ? _GEN_786 : _GEN_2509; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2591 = unuse_way == 3'h2 ? _GEN_787 : _GEN_2316; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2592 = unuse_way == 3'h2 ? _GEN_788 : _GEN_2317; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2593 = unuse_way == 3'h2 ? _GEN_789 : _GEN_2318; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2594 = unuse_way == 3'h2 ? _GEN_790 : _GEN_2319; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2595 = unuse_way == 3'h2 ? _GEN_791 : _GEN_2320; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2596 = unuse_way == 3'h2 ? _GEN_792 : _GEN_2321; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2597 = unuse_way == 3'h2 ? _GEN_793 : _GEN_2322; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2598 = unuse_way == 3'h2 ? _GEN_794 : _GEN_2323; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2599 = unuse_way == 3'h2 ? _GEN_795 : _GEN_2324; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2600 = unuse_way == 3'h2 ? _GEN_796 : _GEN_2325; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2601 = unuse_way == 3'h2 ? _GEN_797 : _GEN_2326; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2602 = unuse_way == 3'h2 ? _GEN_798 : _GEN_2327; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2603 = unuse_way == 3'h2 ? _GEN_799 : _GEN_2328; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2604 = unuse_way == 3'h2 ? _GEN_800 : _GEN_2329; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2605 = unuse_way == 3'h2 ? _GEN_801 : _GEN_2330; // @[d_cache.scala 150:40]
  wire [7:0] _GEN_2606 = unuse_way == 3'h2 ? _GEN_802 : _GEN_2331; // @[d_cache.scala 150:40]
  wire [127:0] _GEN_2607 = unuse_way == 3'h2 ? ram_2_0 : _GEN_2268; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2608 = unuse_way == 3'h2 ? ram_2_1 : _GEN_2269; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2609 = unuse_way == 3'h2 ? ram_2_2 : _GEN_2270; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2610 = unuse_way == 3'h2 ? ram_2_3 : _GEN_2271; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2611 = unuse_way == 3'h2 ? ram_2_4 : _GEN_2272; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2612 = unuse_way == 3'h2 ? ram_2_5 : _GEN_2273; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2613 = unuse_way == 3'h2 ? ram_2_6 : _GEN_2274; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2614 = unuse_way == 3'h2 ? ram_2_7 : _GEN_2275; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2615 = unuse_way == 3'h2 ? ram_2_8 : _GEN_2276; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2616 = unuse_way == 3'h2 ? ram_2_9 : _GEN_2277; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2617 = unuse_way == 3'h2 ? ram_2_10 : _GEN_2278; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2618 = unuse_way == 3'h2 ? ram_2_11 : _GEN_2279; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2619 = unuse_way == 3'h2 ? ram_2_12 : _GEN_2280; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2620 = unuse_way == 3'h2 ? ram_2_13 : _GEN_2281; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2621 = unuse_way == 3'h2 ? ram_2_14 : _GEN_2282; // @[d_cache.scala 150:40 21:24]
  wire [127:0] _GEN_2622 = unuse_way == 3'h2 ? ram_2_15 : _GEN_2283; // @[d_cache.scala 150:40 21:24]
  wire [31:0] _GEN_2623 = unuse_way == 3'h2 ? tag_2_0 : _GEN_2284; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2624 = unuse_way == 3'h2 ? tag_2_1 : _GEN_2285; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2625 = unuse_way == 3'h2 ? tag_2_2 : _GEN_2286; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2626 = unuse_way == 3'h2 ? tag_2_3 : _GEN_2287; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2627 = unuse_way == 3'h2 ? tag_2_4 : _GEN_2288; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2628 = unuse_way == 3'h2 ? tag_2_5 : _GEN_2289; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2629 = unuse_way == 3'h2 ? tag_2_6 : _GEN_2290; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2630 = unuse_way == 3'h2 ? tag_2_7 : _GEN_2291; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2631 = unuse_way == 3'h2 ? tag_2_8 : _GEN_2292; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2632 = unuse_way == 3'h2 ? tag_2_9 : _GEN_2293; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2633 = unuse_way == 3'h2 ? tag_2_10 : _GEN_2294; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2634 = unuse_way == 3'h2 ? tag_2_11 : _GEN_2295; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2635 = unuse_way == 3'h2 ? tag_2_12 : _GEN_2296; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2636 = unuse_way == 3'h2 ? tag_2_13 : _GEN_2297; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2637 = unuse_way == 3'h2 ? tag_2_14 : _GEN_2298; // @[d_cache.scala 150:40 26:24]
  wire [31:0] _GEN_2638 = unuse_way == 3'h2 ? tag_2_15 : _GEN_2299; // @[d_cache.scala 150:40 26:24]
  wire  _GEN_2639 = unuse_way == 3'h2 ? valid_2_0 : _GEN_2300; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2640 = unuse_way == 3'h2 ? valid_2_1 : _GEN_2301; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2641 = unuse_way == 3'h2 ? valid_2_2 : _GEN_2302; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2642 = unuse_way == 3'h2 ? valid_2_3 : _GEN_2303; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2643 = unuse_way == 3'h2 ? valid_2_4 : _GEN_2304; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2644 = unuse_way == 3'h2 ? valid_2_5 : _GEN_2305; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2645 = unuse_way == 3'h2 ? valid_2_6 : _GEN_2306; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2646 = unuse_way == 3'h2 ? valid_2_7 : _GEN_2307; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2647 = unuse_way == 3'h2 ? valid_2_8 : _GEN_2308; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2648 = unuse_way == 3'h2 ? valid_2_9 : _GEN_2309; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2649 = unuse_way == 3'h2 ? valid_2_10 : _GEN_2310; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2650 = unuse_way == 3'h2 ? valid_2_11 : _GEN_2311; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2651 = unuse_way == 3'h2 ? valid_2_12 : _GEN_2312; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2652 = unuse_way == 3'h2 ? valid_2_13 : _GEN_2313; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2653 = unuse_way == 3'h2 ? valid_2_14 : _GEN_2314; // @[d_cache.scala 150:40 30:26]
  wire  _GEN_2654 = unuse_way == 3'h2 ? valid_2_15 : _GEN_2315; // @[d_cache.scala 150:40 30:26]
  wire [127:0] _GEN_2655 = unuse_way == 3'h2 ? ram_3_0 : _GEN_2332; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2656 = unuse_way == 3'h2 ? ram_3_1 : _GEN_2333; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2657 = unuse_way == 3'h2 ? ram_3_2 : _GEN_2334; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2658 = unuse_way == 3'h2 ? ram_3_3 : _GEN_2335; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2659 = unuse_way == 3'h2 ? ram_3_4 : _GEN_2336; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2660 = unuse_way == 3'h2 ? ram_3_5 : _GEN_2337; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2661 = unuse_way == 3'h2 ? ram_3_6 : _GEN_2338; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2662 = unuse_way == 3'h2 ? ram_3_7 : _GEN_2339; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2663 = unuse_way == 3'h2 ? ram_3_8 : _GEN_2340; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2664 = unuse_way == 3'h2 ? ram_3_9 : _GEN_2341; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2665 = unuse_way == 3'h2 ? ram_3_10 : _GEN_2342; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2666 = unuse_way == 3'h2 ? ram_3_11 : _GEN_2343; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2667 = unuse_way == 3'h2 ? ram_3_12 : _GEN_2344; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2668 = unuse_way == 3'h2 ? ram_3_13 : _GEN_2345; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2669 = unuse_way == 3'h2 ? ram_3_14 : _GEN_2346; // @[d_cache.scala 150:40 22:24]
  wire [127:0] _GEN_2670 = unuse_way == 3'h2 ? ram_3_15 : _GEN_2347; // @[d_cache.scala 150:40 22:24]
  wire [31:0] _GEN_2671 = unuse_way == 3'h2 ? tag_3_0 : _GEN_2348; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2672 = unuse_way == 3'h2 ? tag_3_1 : _GEN_2349; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2673 = unuse_way == 3'h2 ? tag_3_2 : _GEN_2350; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2674 = unuse_way == 3'h2 ? tag_3_3 : _GEN_2351; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2675 = unuse_way == 3'h2 ? tag_3_4 : _GEN_2352; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2676 = unuse_way == 3'h2 ? tag_3_5 : _GEN_2353; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2677 = unuse_way == 3'h2 ? tag_3_6 : _GEN_2354; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2678 = unuse_way == 3'h2 ? tag_3_7 : _GEN_2355; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2679 = unuse_way == 3'h2 ? tag_3_8 : _GEN_2356; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2680 = unuse_way == 3'h2 ? tag_3_9 : _GEN_2357; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2681 = unuse_way == 3'h2 ? tag_3_10 : _GEN_2358; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2682 = unuse_way == 3'h2 ? tag_3_11 : _GEN_2359; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2683 = unuse_way == 3'h2 ? tag_3_12 : _GEN_2360; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2684 = unuse_way == 3'h2 ? tag_3_13 : _GEN_2361; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2685 = unuse_way == 3'h2 ? tag_3_14 : _GEN_2362; // @[d_cache.scala 150:40 27:24]
  wire [31:0] _GEN_2686 = unuse_way == 3'h2 ? tag_3_15 : _GEN_2363; // @[d_cache.scala 150:40 27:24]
  wire  _GEN_2687 = unuse_way == 3'h2 ? valid_3_0 : _GEN_2364; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2688 = unuse_way == 3'h2 ? valid_3_1 : _GEN_2365; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2689 = unuse_way == 3'h2 ? valid_3_2 : _GEN_2366; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2690 = unuse_way == 3'h2 ? valid_3_3 : _GEN_2367; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2691 = unuse_way == 3'h2 ? valid_3_4 : _GEN_2368; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2692 = unuse_way == 3'h2 ? valid_3_5 : _GEN_2369; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2693 = unuse_way == 3'h2 ? valid_3_6 : _GEN_2370; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2694 = unuse_way == 3'h2 ? valid_3_7 : _GEN_2371; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2695 = unuse_way == 3'h2 ? valid_3_8 : _GEN_2372; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2696 = unuse_way == 3'h2 ? valid_3_9 : _GEN_2373; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2697 = unuse_way == 3'h2 ? valid_3_10 : _GEN_2374; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2698 = unuse_way == 3'h2 ? valid_3_11 : _GEN_2375; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2699 = unuse_way == 3'h2 ? valid_3_12 : _GEN_2376; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2700 = unuse_way == 3'h2 ? valid_3_13 : _GEN_2377; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2701 = unuse_way == 3'h2 ? valid_3_14 : _GEN_2378; // @[d_cache.scala 150:40 31:26]
  wire  _GEN_2702 = unuse_way == 3'h2 ? valid_3_15 : _GEN_2379; // @[d_cache.scala 150:40 31:26]
  wire [127:0] _GEN_2703 = unuse_way == 3'h2 ? write_back_data : _GEN_2380; // @[d_cache.scala 150:40 41:34]
  wire [39:0] _GEN_2704 = unuse_way == 3'h2 ? {{8'd0}, write_back_addr} : _GEN_2381; // @[d_cache.scala 150:40 42:34]
  wire  _GEN_2705 = unuse_way == 3'h2 ? dirty_0_0 : _GEN_2382; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2706 = unuse_way == 3'h2 ? dirty_0_1 : _GEN_2383; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2707 = unuse_way == 3'h2 ? dirty_0_2 : _GEN_2384; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2708 = unuse_way == 3'h2 ? dirty_0_3 : _GEN_2385; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2709 = unuse_way == 3'h2 ? dirty_0_4 : _GEN_2386; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2710 = unuse_way == 3'h2 ? dirty_0_5 : _GEN_2387; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2711 = unuse_way == 3'h2 ? dirty_0_6 : _GEN_2388; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2712 = unuse_way == 3'h2 ? dirty_0_7 : _GEN_2389; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2713 = unuse_way == 3'h2 ? dirty_0_8 : _GEN_2390; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2714 = unuse_way == 3'h2 ? dirty_0_9 : _GEN_2391; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2715 = unuse_way == 3'h2 ? dirty_0_10 : _GEN_2392; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2716 = unuse_way == 3'h2 ? dirty_0_11 : _GEN_2393; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2717 = unuse_way == 3'h2 ? dirty_0_12 : _GEN_2394; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2718 = unuse_way == 3'h2 ? dirty_0_13 : _GEN_2395; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2719 = unuse_way == 3'h2 ? dirty_0_14 : _GEN_2396; // @[d_cache.scala 150:40 32:26]
  wire  _GEN_2720 = unuse_way == 3'h2 ? dirty_0_15 : _GEN_2397; // @[d_cache.scala 150:40 32:26]
  wire [127:0] _GEN_2721 = unuse_way == 3'h2 ? ram_0_0 : _GEN_2398; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2722 = unuse_way == 3'h2 ? ram_0_1 : _GEN_2399; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2723 = unuse_way == 3'h2 ? ram_0_2 : _GEN_2400; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2724 = unuse_way == 3'h2 ? ram_0_3 : _GEN_2401; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2725 = unuse_way == 3'h2 ? ram_0_4 : _GEN_2402; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2726 = unuse_way == 3'h2 ? ram_0_5 : _GEN_2403; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2727 = unuse_way == 3'h2 ? ram_0_6 : _GEN_2404; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2728 = unuse_way == 3'h2 ? ram_0_7 : _GEN_2405; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2729 = unuse_way == 3'h2 ? ram_0_8 : _GEN_2406; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2730 = unuse_way == 3'h2 ? ram_0_9 : _GEN_2407; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2731 = unuse_way == 3'h2 ? ram_0_10 : _GEN_2408; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2732 = unuse_way == 3'h2 ? ram_0_11 : _GEN_2409; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2733 = unuse_way == 3'h2 ? ram_0_12 : _GEN_2410; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2734 = unuse_way == 3'h2 ? ram_0_13 : _GEN_2411; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2735 = unuse_way == 3'h2 ? ram_0_14 : _GEN_2412; // @[d_cache.scala 150:40 19:24]
  wire [127:0] _GEN_2736 = unuse_way == 3'h2 ? ram_0_15 : _GEN_2413; // @[d_cache.scala 150:40 19:24]
  wire [31:0] _GEN_2737 = unuse_way == 3'h2 ? tag_0_0 : _GEN_2414; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2738 = unuse_way == 3'h2 ? tag_0_1 : _GEN_2415; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2739 = unuse_way == 3'h2 ? tag_0_2 : _GEN_2416; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2740 = unuse_way == 3'h2 ? tag_0_3 : _GEN_2417; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2741 = unuse_way == 3'h2 ? tag_0_4 : _GEN_2418; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2742 = unuse_way == 3'h2 ? tag_0_5 : _GEN_2419; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2743 = unuse_way == 3'h2 ? tag_0_6 : _GEN_2420; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2744 = unuse_way == 3'h2 ? tag_0_7 : _GEN_2421; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2745 = unuse_way == 3'h2 ? tag_0_8 : _GEN_2422; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2746 = unuse_way == 3'h2 ? tag_0_9 : _GEN_2423; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2747 = unuse_way == 3'h2 ? tag_0_10 : _GEN_2424; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2748 = unuse_way == 3'h2 ? tag_0_11 : _GEN_2425; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2749 = unuse_way == 3'h2 ? tag_0_12 : _GEN_2426; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2750 = unuse_way == 3'h2 ? tag_0_13 : _GEN_2427; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2751 = unuse_way == 3'h2 ? tag_0_14 : _GEN_2428; // @[d_cache.scala 150:40 24:24]
  wire [31:0] _GEN_2752 = unuse_way == 3'h2 ? tag_0_15 : _GEN_2429; // @[d_cache.scala 150:40 24:24]
  wire  _GEN_2753 = unuse_way == 3'h2 ? valid_0_0 : _GEN_2430; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2754 = unuse_way == 3'h2 ? valid_0_1 : _GEN_2431; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2755 = unuse_way == 3'h2 ? valid_0_2 : _GEN_2432; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2756 = unuse_way == 3'h2 ? valid_0_3 : _GEN_2433; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2757 = unuse_way == 3'h2 ? valid_0_4 : _GEN_2434; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2758 = unuse_way == 3'h2 ? valid_0_5 : _GEN_2435; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2759 = unuse_way == 3'h2 ? valid_0_6 : _GEN_2436; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2760 = unuse_way == 3'h2 ? valid_0_7 : _GEN_2437; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2761 = unuse_way == 3'h2 ? valid_0_8 : _GEN_2438; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2762 = unuse_way == 3'h2 ? valid_0_9 : _GEN_2439; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2763 = unuse_way == 3'h2 ? valid_0_10 : _GEN_2440; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2764 = unuse_way == 3'h2 ? valid_0_11 : _GEN_2441; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2765 = unuse_way == 3'h2 ? valid_0_12 : _GEN_2442; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2766 = unuse_way == 3'h2 ? valid_0_13 : _GEN_2443; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2767 = unuse_way == 3'h2 ? valid_0_14 : _GEN_2444; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2768 = unuse_way == 3'h2 ? valid_0_15 : _GEN_2445; // @[d_cache.scala 150:40 28:26]
  wire  _GEN_2801 = unuse_way == 3'h2 ? dirty_3_0 : _GEN_2526; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2802 = unuse_way == 3'h2 ? dirty_3_1 : _GEN_2527; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2803 = unuse_way == 3'h2 ? dirty_3_2 : _GEN_2528; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2804 = unuse_way == 3'h2 ? dirty_3_3 : _GEN_2529; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2805 = unuse_way == 3'h2 ? dirty_3_4 : _GEN_2530; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2806 = unuse_way == 3'h2 ? dirty_3_5 : _GEN_2531; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2807 = unuse_way == 3'h2 ? dirty_3_6 : _GEN_2532; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2808 = unuse_way == 3'h2 ? dirty_3_7 : _GEN_2533; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2809 = unuse_way == 3'h2 ? dirty_3_8 : _GEN_2534; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2810 = unuse_way == 3'h2 ? dirty_3_9 : _GEN_2535; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2811 = unuse_way == 3'h2 ? dirty_3_10 : _GEN_2536; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2812 = unuse_way == 3'h2 ? dirty_3_11 : _GEN_2537; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2813 = unuse_way == 3'h2 ? dirty_3_12 : _GEN_2538; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2814 = unuse_way == 3'h2 ? dirty_3_13 : _GEN_2539; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2815 = unuse_way == 3'h2 ? dirty_3_14 : _GEN_2540; // @[d_cache.scala 150:40 35:26]
  wire  _GEN_2816 = unuse_way == 3'h2 ? dirty_3_15 : _GEN_2541; // @[d_cache.scala 150:40 35:26]
  wire [3:0] _GEN_2817 = unuse_way == 3'h1 ? 4'h1 : _GEN_2542; // @[d_cache.scala 144:34 145:23]
  wire [127:0] _GEN_2818 = unuse_way == 3'h1 ? _GEN_659 : _GEN_2721; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2819 = unuse_way == 3'h1 ? _GEN_660 : _GEN_2722; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2820 = unuse_way == 3'h1 ? _GEN_661 : _GEN_2723; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2821 = unuse_way == 3'h1 ? _GEN_662 : _GEN_2724; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2822 = unuse_way == 3'h1 ? _GEN_663 : _GEN_2725; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2823 = unuse_way == 3'h1 ? _GEN_664 : _GEN_2726; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2824 = unuse_way == 3'h1 ? _GEN_665 : _GEN_2727; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2825 = unuse_way == 3'h1 ? _GEN_666 : _GEN_2728; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2826 = unuse_way == 3'h1 ? _GEN_667 : _GEN_2729; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2827 = unuse_way == 3'h1 ? _GEN_668 : _GEN_2730; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2828 = unuse_way == 3'h1 ? _GEN_669 : _GEN_2731; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2829 = unuse_way == 3'h1 ? _GEN_670 : _GEN_2732; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2830 = unuse_way == 3'h1 ? _GEN_671 : _GEN_2733; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2831 = unuse_way == 3'h1 ? _GEN_672 : _GEN_2734; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2832 = unuse_way == 3'h1 ? _GEN_673 : _GEN_2735; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2833 = unuse_way == 3'h1 ? _GEN_674 : _GEN_2736; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2834 = unuse_way == 3'h1 ? _GEN_675 : _GEN_2737; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2835 = unuse_way == 3'h1 ? _GEN_676 : _GEN_2738; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2836 = unuse_way == 3'h1 ? _GEN_677 : _GEN_2739; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2837 = unuse_way == 3'h1 ? _GEN_678 : _GEN_2740; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2838 = unuse_way == 3'h1 ? _GEN_679 : _GEN_2741; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2839 = unuse_way == 3'h1 ? _GEN_680 : _GEN_2742; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2840 = unuse_way == 3'h1 ? _GEN_681 : _GEN_2743; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2841 = unuse_way == 3'h1 ? _GEN_682 : _GEN_2744; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2842 = unuse_way == 3'h1 ? _GEN_683 : _GEN_2745; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2843 = unuse_way == 3'h1 ? _GEN_684 : _GEN_2746; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2844 = unuse_way == 3'h1 ? _GEN_685 : _GEN_2747; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2845 = unuse_way == 3'h1 ? _GEN_686 : _GEN_2748; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2846 = unuse_way == 3'h1 ? _GEN_687 : _GEN_2749; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2847 = unuse_way == 3'h1 ? _GEN_688 : _GEN_2750; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2848 = unuse_way == 3'h1 ? _GEN_689 : _GEN_2751; // @[d_cache.scala 144:34]
  wire [31:0] _GEN_2849 = unuse_way == 3'h1 ? _GEN_690 : _GEN_2752; // @[d_cache.scala 144:34]
  wire  _GEN_2850 = unuse_way == 3'h1 ? _GEN_691 : _GEN_2753; // @[d_cache.scala 144:34]
  wire  _GEN_2851 = unuse_way == 3'h1 ? _GEN_692 : _GEN_2754; // @[d_cache.scala 144:34]
  wire  _GEN_2852 = unuse_way == 3'h1 ? _GEN_693 : _GEN_2755; // @[d_cache.scala 144:34]
  wire  _GEN_2853 = unuse_way == 3'h1 ? _GEN_694 : _GEN_2756; // @[d_cache.scala 144:34]
  wire  _GEN_2854 = unuse_way == 3'h1 ? _GEN_695 : _GEN_2757; // @[d_cache.scala 144:34]
  wire  _GEN_2855 = unuse_way == 3'h1 ? _GEN_696 : _GEN_2758; // @[d_cache.scala 144:34]
  wire  _GEN_2856 = unuse_way == 3'h1 ? _GEN_697 : _GEN_2759; // @[d_cache.scala 144:34]
  wire  _GEN_2857 = unuse_way == 3'h1 ? _GEN_698 : _GEN_2760; // @[d_cache.scala 144:34]
  wire  _GEN_2858 = unuse_way == 3'h1 ? _GEN_699 : _GEN_2761; // @[d_cache.scala 144:34]
  wire  _GEN_2859 = unuse_way == 3'h1 ? _GEN_700 : _GEN_2762; // @[d_cache.scala 144:34]
  wire  _GEN_2860 = unuse_way == 3'h1 ? _GEN_701 : _GEN_2763; // @[d_cache.scala 144:34]
  wire  _GEN_2861 = unuse_way == 3'h1 ? _GEN_702 : _GEN_2764; // @[d_cache.scala 144:34]
  wire  _GEN_2862 = unuse_way == 3'h1 ? _GEN_703 : _GEN_2765; // @[d_cache.scala 144:34]
  wire  _GEN_2863 = unuse_way == 3'h1 ? _GEN_704 : _GEN_2766; // @[d_cache.scala 144:34]
  wire  _GEN_2864 = unuse_way == 3'h1 ? _GEN_705 : _GEN_2767; // @[d_cache.scala 144:34]
  wire  _GEN_2865 = unuse_way == 3'h1 ? _GEN_706 : _GEN_2768; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2866 = unuse_way == 3'h1 ? _GEN_723 : _GEN_2591; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2867 = unuse_way == 3'h1 ? _GEN_724 : _GEN_2592; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2868 = unuse_way == 3'h1 ? _GEN_725 : _GEN_2593; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2869 = unuse_way == 3'h1 ? _GEN_726 : _GEN_2594; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2870 = unuse_way == 3'h1 ? _GEN_727 : _GEN_2595; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2871 = unuse_way == 3'h1 ? _GEN_728 : _GEN_2596; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2872 = unuse_way == 3'h1 ? _GEN_729 : _GEN_2597; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2873 = unuse_way == 3'h1 ? _GEN_730 : _GEN_2598; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2874 = unuse_way == 3'h1 ? _GEN_731 : _GEN_2599; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2875 = unuse_way == 3'h1 ? _GEN_732 : _GEN_2600; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2876 = unuse_way == 3'h1 ? _GEN_733 : _GEN_2601; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2877 = unuse_way == 3'h1 ? _GEN_734 : _GEN_2602; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2878 = unuse_way == 3'h1 ? _GEN_735 : _GEN_2603; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2879 = unuse_way == 3'h1 ? _GEN_736 : _GEN_2604; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2880 = unuse_way == 3'h1 ? _GEN_737 : _GEN_2605; // @[d_cache.scala 144:34]
  wire [7:0] _GEN_2881 = unuse_way == 3'h1 ? _GEN_738 : _GEN_2606; // @[d_cache.scala 144:34]
  wire [127:0] _GEN_2882 = unuse_way == 3'h1 ? ram_1_0 : _GEN_2543; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2883 = unuse_way == 3'h1 ? ram_1_1 : _GEN_2544; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2884 = unuse_way == 3'h1 ? ram_1_2 : _GEN_2545; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2885 = unuse_way == 3'h1 ? ram_1_3 : _GEN_2546; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2886 = unuse_way == 3'h1 ? ram_1_4 : _GEN_2547; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2887 = unuse_way == 3'h1 ? ram_1_5 : _GEN_2548; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2888 = unuse_way == 3'h1 ? ram_1_6 : _GEN_2549; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2889 = unuse_way == 3'h1 ? ram_1_7 : _GEN_2550; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2890 = unuse_way == 3'h1 ? ram_1_8 : _GEN_2551; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2891 = unuse_way == 3'h1 ? ram_1_9 : _GEN_2552; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2892 = unuse_way == 3'h1 ? ram_1_10 : _GEN_2553; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2893 = unuse_way == 3'h1 ? ram_1_11 : _GEN_2554; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2894 = unuse_way == 3'h1 ? ram_1_12 : _GEN_2555; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2895 = unuse_way == 3'h1 ? ram_1_13 : _GEN_2556; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2896 = unuse_way == 3'h1 ? ram_1_14 : _GEN_2557; // @[d_cache.scala 144:34 20:24]
  wire [127:0] _GEN_2897 = unuse_way == 3'h1 ? ram_1_15 : _GEN_2558; // @[d_cache.scala 144:34 20:24]
  wire [31:0] _GEN_2898 = unuse_way == 3'h1 ? tag_1_0 : _GEN_2559; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2899 = unuse_way == 3'h1 ? tag_1_1 : _GEN_2560; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2900 = unuse_way == 3'h1 ? tag_1_2 : _GEN_2561; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2901 = unuse_way == 3'h1 ? tag_1_3 : _GEN_2562; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2902 = unuse_way == 3'h1 ? tag_1_4 : _GEN_2563; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2903 = unuse_way == 3'h1 ? tag_1_5 : _GEN_2564; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2904 = unuse_way == 3'h1 ? tag_1_6 : _GEN_2565; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2905 = unuse_way == 3'h1 ? tag_1_7 : _GEN_2566; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2906 = unuse_way == 3'h1 ? tag_1_8 : _GEN_2567; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2907 = unuse_way == 3'h1 ? tag_1_9 : _GEN_2568; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2908 = unuse_way == 3'h1 ? tag_1_10 : _GEN_2569; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2909 = unuse_way == 3'h1 ? tag_1_11 : _GEN_2570; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2910 = unuse_way == 3'h1 ? tag_1_12 : _GEN_2571; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2911 = unuse_way == 3'h1 ? tag_1_13 : _GEN_2572; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2912 = unuse_way == 3'h1 ? tag_1_14 : _GEN_2573; // @[d_cache.scala 144:34 25:24]
  wire [31:0] _GEN_2913 = unuse_way == 3'h1 ? tag_1_15 : _GEN_2574; // @[d_cache.scala 144:34 25:24]
  wire  _GEN_2914 = unuse_way == 3'h1 ? valid_1_0 : _GEN_2575; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2915 = unuse_way == 3'h1 ? valid_1_1 : _GEN_2576; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2916 = unuse_way == 3'h1 ? valid_1_2 : _GEN_2577; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2917 = unuse_way == 3'h1 ? valid_1_3 : _GEN_2578; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2918 = unuse_way == 3'h1 ? valid_1_4 : _GEN_2579; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2919 = unuse_way == 3'h1 ? valid_1_5 : _GEN_2580; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2920 = unuse_way == 3'h1 ? valid_1_6 : _GEN_2581; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2921 = unuse_way == 3'h1 ? valid_1_7 : _GEN_2582; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2922 = unuse_way == 3'h1 ? valid_1_8 : _GEN_2583; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2923 = unuse_way == 3'h1 ? valid_1_9 : _GEN_2584; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2924 = unuse_way == 3'h1 ? valid_1_10 : _GEN_2585; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2925 = unuse_way == 3'h1 ? valid_1_11 : _GEN_2586; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2926 = unuse_way == 3'h1 ? valid_1_12 : _GEN_2587; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2927 = unuse_way == 3'h1 ? valid_1_13 : _GEN_2588; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2928 = unuse_way == 3'h1 ? valid_1_14 : _GEN_2589; // @[d_cache.scala 144:34 29:26]
  wire  _GEN_2929 = unuse_way == 3'h1 ? valid_1_15 : _GEN_2590; // @[d_cache.scala 144:34 29:26]
  wire [127:0] _GEN_2930 = unuse_way == 3'h1 ? ram_2_0 : _GEN_2607; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2931 = unuse_way == 3'h1 ? ram_2_1 : _GEN_2608; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2932 = unuse_way == 3'h1 ? ram_2_2 : _GEN_2609; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2933 = unuse_way == 3'h1 ? ram_2_3 : _GEN_2610; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2934 = unuse_way == 3'h1 ? ram_2_4 : _GEN_2611; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2935 = unuse_way == 3'h1 ? ram_2_5 : _GEN_2612; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2936 = unuse_way == 3'h1 ? ram_2_6 : _GEN_2613; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2937 = unuse_way == 3'h1 ? ram_2_7 : _GEN_2614; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2938 = unuse_way == 3'h1 ? ram_2_8 : _GEN_2615; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2939 = unuse_way == 3'h1 ? ram_2_9 : _GEN_2616; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2940 = unuse_way == 3'h1 ? ram_2_10 : _GEN_2617; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2941 = unuse_way == 3'h1 ? ram_2_11 : _GEN_2618; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2942 = unuse_way == 3'h1 ? ram_2_12 : _GEN_2619; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2943 = unuse_way == 3'h1 ? ram_2_13 : _GEN_2620; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2944 = unuse_way == 3'h1 ? ram_2_14 : _GEN_2621; // @[d_cache.scala 144:34 21:24]
  wire [127:0] _GEN_2945 = unuse_way == 3'h1 ? ram_2_15 : _GEN_2622; // @[d_cache.scala 144:34 21:24]
  wire [31:0] _GEN_2946 = unuse_way == 3'h1 ? tag_2_0 : _GEN_2623; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2947 = unuse_way == 3'h1 ? tag_2_1 : _GEN_2624; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2948 = unuse_way == 3'h1 ? tag_2_2 : _GEN_2625; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2949 = unuse_way == 3'h1 ? tag_2_3 : _GEN_2626; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2950 = unuse_way == 3'h1 ? tag_2_4 : _GEN_2627; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2951 = unuse_way == 3'h1 ? tag_2_5 : _GEN_2628; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2952 = unuse_way == 3'h1 ? tag_2_6 : _GEN_2629; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2953 = unuse_way == 3'h1 ? tag_2_7 : _GEN_2630; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2954 = unuse_way == 3'h1 ? tag_2_8 : _GEN_2631; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2955 = unuse_way == 3'h1 ? tag_2_9 : _GEN_2632; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2956 = unuse_way == 3'h1 ? tag_2_10 : _GEN_2633; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2957 = unuse_way == 3'h1 ? tag_2_11 : _GEN_2634; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2958 = unuse_way == 3'h1 ? tag_2_12 : _GEN_2635; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2959 = unuse_way == 3'h1 ? tag_2_13 : _GEN_2636; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2960 = unuse_way == 3'h1 ? tag_2_14 : _GEN_2637; // @[d_cache.scala 144:34 26:24]
  wire [31:0] _GEN_2961 = unuse_way == 3'h1 ? tag_2_15 : _GEN_2638; // @[d_cache.scala 144:34 26:24]
  wire  _GEN_2962 = unuse_way == 3'h1 ? valid_2_0 : _GEN_2639; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2963 = unuse_way == 3'h1 ? valid_2_1 : _GEN_2640; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2964 = unuse_way == 3'h1 ? valid_2_2 : _GEN_2641; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2965 = unuse_way == 3'h1 ? valid_2_3 : _GEN_2642; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2966 = unuse_way == 3'h1 ? valid_2_4 : _GEN_2643; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2967 = unuse_way == 3'h1 ? valid_2_5 : _GEN_2644; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2968 = unuse_way == 3'h1 ? valid_2_6 : _GEN_2645; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2969 = unuse_way == 3'h1 ? valid_2_7 : _GEN_2646; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2970 = unuse_way == 3'h1 ? valid_2_8 : _GEN_2647; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2971 = unuse_way == 3'h1 ? valid_2_9 : _GEN_2648; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2972 = unuse_way == 3'h1 ? valid_2_10 : _GEN_2649; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2973 = unuse_way == 3'h1 ? valid_2_11 : _GEN_2650; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2974 = unuse_way == 3'h1 ? valid_2_12 : _GEN_2651; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2975 = unuse_way == 3'h1 ? valid_2_13 : _GEN_2652; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2976 = unuse_way == 3'h1 ? valid_2_14 : _GEN_2653; // @[d_cache.scala 144:34 30:26]
  wire  _GEN_2977 = unuse_way == 3'h1 ? valid_2_15 : _GEN_2654; // @[d_cache.scala 144:34 30:26]
  wire [127:0] _GEN_2978 = unuse_way == 3'h1 ? ram_3_0 : _GEN_2655; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2979 = unuse_way == 3'h1 ? ram_3_1 : _GEN_2656; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2980 = unuse_way == 3'h1 ? ram_3_2 : _GEN_2657; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2981 = unuse_way == 3'h1 ? ram_3_3 : _GEN_2658; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2982 = unuse_way == 3'h1 ? ram_3_4 : _GEN_2659; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2983 = unuse_way == 3'h1 ? ram_3_5 : _GEN_2660; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2984 = unuse_way == 3'h1 ? ram_3_6 : _GEN_2661; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2985 = unuse_way == 3'h1 ? ram_3_7 : _GEN_2662; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2986 = unuse_way == 3'h1 ? ram_3_8 : _GEN_2663; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2987 = unuse_way == 3'h1 ? ram_3_9 : _GEN_2664; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2988 = unuse_way == 3'h1 ? ram_3_10 : _GEN_2665; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2989 = unuse_way == 3'h1 ? ram_3_11 : _GEN_2666; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2990 = unuse_way == 3'h1 ? ram_3_12 : _GEN_2667; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2991 = unuse_way == 3'h1 ? ram_3_13 : _GEN_2668; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2992 = unuse_way == 3'h1 ? ram_3_14 : _GEN_2669; // @[d_cache.scala 144:34 22:24]
  wire [127:0] _GEN_2993 = unuse_way == 3'h1 ? ram_3_15 : _GEN_2670; // @[d_cache.scala 144:34 22:24]
  wire [31:0] _GEN_2994 = unuse_way == 3'h1 ? tag_3_0 : _GEN_2671; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_2995 = unuse_way == 3'h1 ? tag_3_1 : _GEN_2672; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_2996 = unuse_way == 3'h1 ? tag_3_2 : _GEN_2673; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_2997 = unuse_way == 3'h1 ? tag_3_3 : _GEN_2674; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_2998 = unuse_way == 3'h1 ? tag_3_4 : _GEN_2675; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_2999 = unuse_way == 3'h1 ? tag_3_5 : _GEN_2676; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_3000 = unuse_way == 3'h1 ? tag_3_6 : _GEN_2677; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_3001 = unuse_way == 3'h1 ? tag_3_7 : _GEN_2678; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_3002 = unuse_way == 3'h1 ? tag_3_8 : _GEN_2679; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_3003 = unuse_way == 3'h1 ? tag_3_9 : _GEN_2680; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_3004 = unuse_way == 3'h1 ? tag_3_10 : _GEN_2681; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_3005 = unuse_way == 3'h1 ? tag_3_11 : _GEN_2682; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_3006 = unuse_way == 3'h1 ? tag_3_12 : _GEN_2683; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_3007 = unuse_way == 3'h1 ? tag_3_13 : _GEN_2684; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_3008 = unuse_way == 3'h1 ? tag_3_14 : _GEN_2685; // @[d_cache.scala 144:34 27:24]
  wire [31:0] _GEN_3009 = unuse_way == 3'h1 ? tag_3_15 : _GEN_2686; // @[d_cache.scala 144:34 27:24]
  wire  _GEN_3010 = unuse_way == 3'h1 ? valid_3_0 : _GEN_2687; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3011 = unuse_way == 3'h1 ? valid_3_1 : _GEN_2688; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3012 = unuse_way == 3'h1 ? valid_3_2 : _GEN_2689; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3013 = unuse_way == 3'h1 ? valid_3_3 : _GEN_2690; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3014 = unuse_way == 3'h1 ? valid_3_4 : _GEN_2691; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3015 = unuse_way == 3'h1 ? valid_3_5 : _GEN_2692; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3016 = unuse_way == 3'h1 ? valid_3_6 : _GEN_2693; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3017 = unuse_way == 3'h1 ? valid_3_7 : _GEN_2694; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3018 = unuse_way == 3'h1 ? valid_3_8 : _GEN_2695; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3019 = unuse_way == 3'h1 ? valid_3_9 : _GEN_2696; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3020 = unuse_way == 3'h1 ? valid_3_10 : _GEN_2697; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3021 = unuse_way == 3'h1 ? valid_3_11 : _GEN_2698; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3022 = unuse_way == 3'h1 ? valid_3_12 : _GEN_2699; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3023 = unuse_way == 3'h1 ? valid_3_13 : _GEN_2700; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3024 = unuse_way == 3'h1 ? valid_3_14 : _GEN_2701; // @[d_cache.scala 144:34 31:26]
  wire  _GEN_3025 = unuse_way == 3'h1 ? valid_3_15 : _GEN_2702; // @[d_cache.scala 144:34 31:26]
  wire [127:0] _GEN_3026 = unuse_way == 3'h1 ? write_back_data : _GEN_2703; // @[d_cache.scala 144:34 41:34]
  wire [39:0] _GEN_3027 = unuse_way == 3'h1 ? {{8'd0}, write_back_addr} : _GEN_2704; // @[d_cache.scala 144:34 42:34]
  wire  _GEN_3028 = unuse_way == 3'h1 ? dirty_0_0 : _GEN_2705; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3029 = unuse_way == 3'h1 ? dirty_0_1 : _GEN_2706; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3030 = unuse_way == 3'h1 ? dirty_0_2 : _GEN_2707; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3031 = unuse_way == 3'h1 ? dirty_0_3 : _GEN_2708; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3032 = unuse_way == 3'h1 ? dirty_0_4 : _GEN_2709; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3033 = unuse_way == 3'h1 ? dirty_0_5 : _GEN_2710; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3034 = unuse_way == 3'h1 ? dirty_0_6 : _GEN_2711; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3035 = unuse_way == 3'h1 ? dirty_0_7 : _GEN_2712; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3036 = unuse_way == 3'h1 ? dirty_0_8 : _GEN_2713; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3037 = unuse_way == 3'h1 ? dirty_0_9 : _GEN_2714; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3038 = unuse_way == 3'h1 ? dirty_0_10 : _GEN_2715; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3039 = unuse_way == 3'h1 ? dirty_0_11 : _GEN_2716; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3040 = unuse_way == 3'h1 ? dirty_0_12 : _GEN_2717; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3041 = unuse_way == 3'h1 ? dirty_0_13 : _GEN_2718; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3042 = unuse_way == 3'h1 ? dirty_0_14 : _GEN_2719; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3043 = unuse_way == 3'h1 ? dirty_0_15 : _GEN_2720; // @[d_cache.scala 144:34 32:26]
  wire  _GEN_3076 = unuse_way == 3'h1 ? dirty_3_0 : _GEN_2801; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3077 = unuse_way == 3'h1 ? dirty_3_1 : _GEN_2802; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3078 = unuse_way == 3'h1 ? dirty_3_2 : _GEN_2803; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3079 = unuse_way == 3'h1 ? dirty_3_3 : _GEN_2804; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3080 = unuse_way == 3'h1 ? dirty_3_4 : _GEN_2805; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3081 = unuse_way == 3'h1 ? dirty_3_5 : _GEN_2806; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3082 = unuse_way == 3'h1 ? dirty_3_6 : _GEN_2807; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3083 = unuse_way == 3'h1 ? dirty_3_7 : _GEN_2808; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3084 = unuse_way == 3'h1 ? dirty_3_8 : _GEN_2809; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3085 = unuse_way == 3'h1 ? dirty_3_9 : _GEN_2810; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3086 = unuse_way == 3'h1 ? dirty_3_10 : _GEN_2811; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3087 = unuse_way == 3'h1 ? dirty_3_11 : _GEN_2812; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3088 = unuse_way == 3'h1 ? dirty_3_12 : _GEN_2813; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3089 = unuse_way == 3'h1 ? dirty_3_13 : _GEN_2814; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3090 = unuse_way == 3'h1 ? dirty_3_14 : _GEN_2815; // @[d_cache.scala 144:34 35:26]
  wire  _GEN_3091 = unuse_way == 3'h1 ? dirty_3_15 : _GEN_2816; // @[d_cache.scala 144:34 35:26]
  wire [127:0] _write_back_data_T = {{64'd0}, write_back_data[127:64]}; // @[d_cache.scala 227:52]
  wire [127:0] _GEN_3092 = io_from_axi_wready ? _write_back_data_T : write_back_data; // @[d_cache.scala 226:37 227:33 41:34]
  wire [3:0] _GEN_3093 = io_from_axi_bvalid ? 4'h1 : state; // @[d_cache.scala 229:37 230:23 71:24]
  wire [3:0] _GEN_3094 = io_from_axi_rvalid ? 4'h0 : state; // @[d_cache.scala 234:37 235:23 71:24]
  wire [3:0] _GEN_3096 = 4'h8 == state ? _GEN_658 : state; // @[d_cache.scala 76:18 71:24]
  wire [3:0] _GEN_3097 = 4'h7 == state ? _GEN_3094 : _GEN_3096; // @[d_cache.scala 76:18]
  wire [127:0] _GEN_3098 = 4'h6 == state ? _GEN_3092 : write_back_data; // @[d_cache.scala 76:18 41:34]
  wire [3:0] _GEN_3099 = 4'h6 == state ? _GEN_3093 : _GEN_3097; // @[d_cache.scala 76:18]
  wire [3:0] _GEN_3100 = 4'h5 == state ? _GEN_2817 : _GEN_3099; // @[d_cache.scala 76:18]
  wire [127:0] _GEN_3101 = 4'h5 == state ? _GEN_2818 : ram_0_0; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3102 = 4'h5 == state ? _GEN_2819 : ram_0_1; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3103 = 4'h5 == state ? _GEN_2820 : ram_0_2; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3104 = 4'h5 == state ? _GEN_2821 : ram_0_3; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3105 = 4'h5 == state ? _GEN_2822 : ram_0_4; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3106 = 4'h5 == state ? _GEN_2823 : ram_0_5; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3107 = 4'h5 == state ? _GEN_2824 : ram_0_6; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3108 = 4'h5 == state ? _GEN_2825 : ram_0_7; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3109 = 4'h5 == state ? _GEN_2826 : ram_0_8; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3110 = 4'h5 == state ? _GEN_2827 : ram_0_9; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3111 = 4'h5 == state ? _GEN_2828 : ram_0_10; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3112 = 4'h5 == state ? _GEN_2829 : ram_0_11; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3113 = 4'h5 == state ? _GEN_2830 : ram_0_12; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3114 = 4'h5 == state ? _GEN_2831 : ram_0_13; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3115 = 4'h5 == state ? _GEN_2832 : ram_0_14; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3116 = 4'h5 == state ? _GEN_2833 : ram_0_15; // @[d_cache.scala 76:18 19:24]
  wire [31:0] _GEN_3117 = 4'h5 == state ? _GEN_2834 : tag_0_0; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3118 = 4'h5 == state ? _GEN_2835 : tag_0_1; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3119 = 4'h5 == state ? _GEN_2836 : tag_0_2; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3120 = 4'h5 == state ? _GEN_2837 : tag_0_3; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3121 = 4'h5 == state ? _GEN_2838 : tag_0_4; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3122 = 4'h5 == state ? _GEN_2839 : tag_0_5; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3123 = 4'h5 == state ? _GEN_2840 : tag_0_6; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3124 = 4'h5 == state ? _GEN_2841 : tag_0_7; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3125 = 4'h5 == state ? _GEN_2842 : tag_0_8; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3126 = 4'h5 == state ? _GEN_2843 : tag_0_9; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3127 = 4'h5 == state ? _GEN_2844 : tag_0_10; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3128 = 4'h5 == state ? _GEN_2845 : tag_0_11; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3129 = 4'h5 == state ? _GEN_2846 : tag_0_12; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3130 = 4'h5 == state ? _GEN_2847 : tag_0_13; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3131 = 4'h5 == state ? _GEN_2848 : tag_0_14; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3132 = 4'h5 == state ? _GEN_2849 : tag_0_15; // @[d_cache.scala 76:18 24:24]
  wire  _GEN_3133 = 4'h5 == state ? _GEN_2850 : valid_0_0; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3134 = 4'h5 == state ? _GEN_2851 : valid_0_1; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3135 = 4'h5 == state ? _GEN_2852 : valid_0_2; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3136 = 4'h5 == state ? _GEN_2853 : valid_0_3; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3137 = 4'h5 == state ? _GEN_2854 : valid_0_4; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3138 = 4'h5 == state ? _GEN_2855 : valid_0_5; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3139 = 4'h5 == state ? _GEN_2856 : valid_0_6; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3140 = 4'h5 == state ? _GEN_2857 : valid_0_7; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3141 = 4'h5 == state ? _GEN_2858 : valid_0_8; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3142 = 4'h5 == state ? _GEN_2859 : valid_0_9; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3143 = 4'h5 == state ? _GEN_2860 : valid_0_10; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3144 = 4'h5 == state ? _GEN_2861 : valid_0_11; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3145 = 4'h5 == state ? _GEN_2862 : valid_0_12; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3146 = 4'h5 == state ? _GEN_2863 : valid_0_13; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3147 = 4'h5 == state ? _GEN_2864 : valid_0_14; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3148 = 4'h5 == state ? _GEN_2865 : valid_0_15; // @[d_cache.scala 76:18 28:26]
  wire [7:0] _GEN_3149 = 4'h5 == state ? _GEN_2866 : quene_0; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3150 = 4'h5 == state ? _GEN_2867 : quene_1; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3151 = 4'h5 == state ? _GEN_2868 : quene_2; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3152 = 4'h5 == state ? _GEN_2869 : quene_3; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3153 = 4'h5 == state ? _GEN_2870 : quene_4; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3154 = 4'h5 == state ? _GEN_2871 : quene_5; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3155 = 4'h5 == state ? _GEN_2872 : quene_6; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3156 = 4'h5 == state ? _GEN_2873 : quene_7; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3157 = 4'h5 == state ? _GEN_2874 : quene_8; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3158 = 4'h5 == state ? _GEN_2875 : quene_9; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3159 = 4'h5 == state ? _GEN_2876 : quene_10; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3160 = 4'h5 == state ? _GEN_2877 : quene_11; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3161 = 4'h5 == state ? _GEN_2878 : quene_12; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3162 = 4'h5 == state ? _GEN_2879 : quene_13; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3163 = 4'h5 == state ? _GEN_2880 : quene_14; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3164 = 4'h5 == state ? _GEN_2881 : quene_15; // @[d_cache.scala 76:18 49:24]
  wire [127:0] _GEN_3165 = 4'h5 == state ? _GEN_2882 : ram_1_0; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3166 = 4'h5 == state ? _GEN_2883 : ram_1_1; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3167 = 4'h5 == state ? _GEN_2884 : ram_1_2; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3168 = 4'h5 == state ? _GEN_2885 : ram_1_3; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3169 = 4'h5 == state ? _GEN_2886 : ram_1_4; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3170 = 4'h5 == state ? _GEN_2887 : ram_1_5; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3171 = 4'h5 == state ? _GEN_2888 : ram_1_6; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3172 = 4'h5 == state ? _GEN_2889 : ram_1_7; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3173 = 4'h5 == state ? _GEN_2890 : ram_1_8; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3174 = 4'h5 == state ? _GEN_2891 : ram_1_9; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3175 = 4'h5 == state ? _GEN_2892 : ram_1_10; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3176 = 4'h5 == state ? _GEN_2893 : ram_1_11; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3177 = 4'h5 == state ? _GEN_2894 : ram_1_12; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3178 = 4'h5 == state ? _GEN_2895 : ram_1_13; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3179 = 4'h5 == state ? _GEN_2896 : ram_1_14; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3180 = 4'h5 == state ? _GEN_2897 : ram_1_15; // @[d_cache.scala 76:18 20:24]
  wire [31:0] _GEN_3181 = 4'h5 == state ? _GEN_2898 : tag_1_0; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3182 = 4'h5 == state ? _GEN_2899 : tag_1_1; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3183 = 4'h5 == state ? _GEN_2900 : tag_1_2; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3184 = 4'h5 == state ? _GEN_2901 : tag_1_3; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3185 = 4'h5 == state ? _GEN_2902 : tag_1_4; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3186 = 4'h5 == state ? _GEN_2903 : tag_1_5; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3187 = 4'h5 == state ? _GEN_2904 : tag_1_6; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3188 = 4'h5 == state ? _GEN_2905 : tag_1_7; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3189 = 4'h5 == state ? _GEN_2906 : tag_1_8; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3190 = 4'h5 == state ? _GEN_2907 : tag_1_9; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3191 = 4'h5 == state ? _GEN_2908 : tag_1_10; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3192 = 4'h5 == state ? _GEN_2909 : tag_1_11; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3193 = 4'h5 == state ? _GEN_2910 : tag_1_12; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3194 = 4'h5 == state ? _GEN_2911 : tag_1_13; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3195 = 4'h5 == state ? _GEN_2912 : tag_1_14; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3196 = 4'h5 == state ? _GEN_2913 : tag_1_15; // @[d_cache.scala 76:18 25:24]
  wire  _GEN_3197 = 4'h5 == state ? _GEN_2914 : valid_1_0; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3198 = 4'h5 == state ? _GEN_2915 : valid_1_1; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3199 = 4'h5 == state ? _GEN_2916 : valid_1_2; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3200 = 4'h5 == state ? _GEN_2917 : valid_1_3; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3201 = 4'h5 == state ? _GEN_2918 : valid_1_4; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3202 = 4'h5 == state ? _GEN_2919 : valid_1_5; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3203 = 4'h5 == state ? _GEN_2920 : valid_1_6; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3204 = 4'h5 == state ? _GEN_2921 : valid_1_7; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3205 = 4'h5 == state ? _GEN_2922 : valid_1_8; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3206 = 4'h5 == state ? _GEN_2923 : valid_1_9; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3207 = 4'h5 == state ? _GEN_2924 : valid_1_10; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3208 = 4'h5 == state ? _GEN_2925 : valid_1_11; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3209 = 4'h5 == state ? _GEN_2926 : valid_1_12; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3210 = 4'h5 == state ? _GEN_2927 : valid_1_13; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3211 = 4'h5 == state ? _GEN_2928 : valid_1_14; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3212 = 4'h5 == state ? _GEN_2929 : valid_1_15; // @[d_cache.scala 76:18 29:26]
  wire [127:0] _GEN_3213 = 4'h5 == state ? _GEN_2930 : ram_2_0; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3214 = 4'h5 == state ? _GEN_2931 : ram_2_1; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3215 = 4'h5 == state ? _GEN_2932 : ram_2_2; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3216 = 4'h5 == state ? _GEN_2933 : ram_2_3; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3217 = 4'h5 == state ? _GEN_2934 : ram_2_4; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3218 = 4'h5 == state ? _GEN_2935 : ram_2_5; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3219 = 4'h5 == state ? _GEN_2936 : ram_2_6; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3220 = 4'h5 == state ? _GEN_2937 : ram_2_7; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3221 = 4'h5 == state ? _GEN_2938 : ram_2_8; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3222 = 4'h5 == state ? _GEN_2939 : ram_2_9; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3223 = 4'h5 == state ? _GEN_2940 : ram_2_10; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3224 = 4'h5 == state ? _GEN_2941 : ram_2_11; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3225 = 4'h5 == state ? _GEN_2942 : ram_2_12; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3226 = 4'h5 == state ? _GEN_2943 : ram_2_13; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3227 = 4'h5 == state ? _GEN_2944 : ram_2_14; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3228 = 4'h5 == state ? _GEN_2945 : ram_2_15; // @[d_cache.scala 76:18 21:24]
  wire [31:0] _GEN_3229 = 4'h5 == state ? _GEN_2946 : tag_2_0; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3230 = 4'h5 == state ? _GEN_2947 : tag_2_1; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3231 = 4'h5 == state ? _GEN_2948 : tag_2_2; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3232 = 4'h5 == state ? _GEN_2949 : tag_2_3; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3233 = 4'h5 == state ? _GEN_2950 : tag_2_4; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3234 = 4'h5 == state ? _GEN_2951 : tag_2_5; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3235 = 4'h5 == state ? _GEN_2952 : tag_2_6; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3236 = 4'h5 == state ? _GEN_2953 : tag_2_7; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3237 = 4'h5 == state ? _GEN_2954 : tag_2_8; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3238 = 4'h5 == state ? _GEN_2955 : tag_2_9; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3239 = 4'h5 == state ? _GEN_2956 : tag_2_10; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3240 = 4'h5 == state ? _GEN_2957 : tag_2_11; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3241 = 4'h5 == state ? _GEN_2958 : tag_2_12; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3242 = 4'h5 == state ? _GEN_2959 : tag_2_13; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3243 = 4'h5 == state ? _GEN_2960 : tag_2_14; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3244 = 4'h5 == state ? _GEN_2961 : tag_2_15; // @[d_cache.scala 76:18 26:24]
  wire  _GEN_3245 = 4'h5 == state ? _GEN_2962 : valid_2_0; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3246 = 4'h5 == state ? _GEN_2963 : valid_2_1; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3247 = 4'h5 == state ? _GEN_2964 : valid_2_2; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3248 = 4'h5 == state ? _GEN_2965 : valid_2_3; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3249 = 4'h5 == state ? _GEN_2966 : valid_2_4; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3250 = 4'h5 == state ? _GEN_2967 : valid_2_5; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3251 = 4'h5 == state ? _GEN_2968 : valid_2_6; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3252 = 4'h5 == state ? _GEN_2969 : valid_2_7; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3253 = 4'h5 == state ? _GEN_2970 : valid_2_8; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3254 = 4'h5 == state ? _GEN_2971 : valid_2_9; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3255 = 4'h5 == state ? _GEN_2972 : valid_2_10; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3256 = 4'h5 == state ? _GEN_2973 : valid_2_11; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3257 = 4'h5 == state ? _GEN_2974 : valid_2_12; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3258 = 4'h5 == state ? _GEN_2975 : valid_2_13; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3259 = 4'h5 == state ? _GEN_2976 : valid_2_14; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3260 = 4'h5 == state ? _GEN_2977 : valid_2_15; // @[d_cache.scala 76:18 30:26]
  wire [127:0] _GEN_3261 = 4'h5 == state ? _GEN_2978 : ram_3_0; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3262 = 4'h5 == state ? _GEN_2979 : ram_3_1; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3263 = 4'h5 == state ? _GEN_2980 : ram_3_2; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3264 = 4'h5 == state ? _GEN_2981 : ram_3_3; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3265 = 4'h5 == state ? _GEN_2982 : ram_3_4; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3266 = 4'h5 == state ? _GEN_2983 : ram_3_5; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3267 = 4'h5 == state ? _GEN_2984 : ram_3_6; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3268 = 4'h5 == state ? _GEN_2985 : ram_3_7; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3269 = 4'h5 == state ? _GEN_2986 : ram_3_8; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3270 = 4'h5 == state ? _GEN_2987 : ram_3_9; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3271 = 4'h5 == state ? _GEN_2988 : ram_3_10; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3272 = 4'h5 == state ? _GEN_2989 : ram_3_11; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3273 = 4'h5 == state ? _GEN_2990 : ram_3_12; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3274 = 4'h5 == state ? _GEN_2991 : ram_3_13; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3275 = 4'h5 == state ? _GEN_2992 : ram_3_14; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3276 = 4'h5 == state ? _GEN_2993 : ram_3_15; // @[d_cache.scala 76:18 22:24]
  wire [31:0] _GEN_3277 = 4'h5 == state ? _GEN_2994 : tag_3_0; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3278 = 4'h5 == state ? _GEN_2995 : tag_3_1; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3279 = 4'h5 == state ? _GEN_2996 : tag_3_2; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3280 = 4'h5 == state ? _GEN_2997 : tag_3_3; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3281 = 4'h5 == state ? _GEN_2998 : tag_3_4; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3282 = 4'h5 == state ? _GEN_2999 : tag_3_5; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3283 = 4'h5 == state ? _GEN_3000 : tag_3_6; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3284 = 4'h5 == state ? _GEN_3001 : tag_3_7; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3285 = 4'h5 == state ? _GEN_3002 : tag_3_8; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3286 = 4'h5 == state ? _GEN_3003 : tag_3_9; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3287 = 4'h5 == state ? _GEN_3004 : tag_3_10; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3288 = 4'h5 == state ? _GEN_3005 : tag_3_11; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3289 = 4'h5 == state ? _GEN_3006 : tag_3_12; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3290 = 4'h5 == state ? _GEN_3007 : tag_3_13; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3291 = 4'h5 == state ? _GEN_3008 : tag_3_14; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3292 = 4'h5 == state ? _GEN_3009 : tag_3_15; // @[d_cache.scala 76:18 27:24]
  wire  _GEN_3293 = 4'h5 == state ? _GEN_3010 : valid_3_0; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3294 = 4'h5 == state ? _GEN_3011 : valid_3_1; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3295 = 4'h5 == state ? _GEN_3012 : valid_3_2; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3296 = 4'h5 == state ? _GEN_3013 : valid_3_3; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3297 = 4'h5 == state ? _GEN_3014 : valid_3_4; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3298 = 4'h5 == state ? _GEN_3015 : valid_3_5; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3299 = 4'h5 == state ? _GEN_3016 : valid_3_6; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3300 = 4'h5 == state ? _GEN_3017 : valid_3_7; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3301 = 4'h5 == state ? _GEN_3018 : valid_3_8; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3302 = 4'h5 == state ? _GEN_3019 : valid_3_9; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3303 = 4'h5 == state ? _GEN_3020 : valid_3_10; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3304 = 4'h5 == state ? _GEN_3021 : valid_3_11; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3305 = 4'h5 == state ? _GEN_3022 : valid_3_12; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3306 = 4'h5 == state ? _GEN_3023 : valid_3_13; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3307 = 4'h5 == state ? _GEN_3024 : valid_3_14; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3308 = 4'h5 == state ? _GEN_3025 : valid_3_15; // @[d_cache.scala 76:18 31:26]
  wire [127:0] _GEN_3309 = 4'h5 == state ? _GEN_3026 : _GEN_3098; // @[d_cache.scala 76:18]
  wire [39:0] _GEN_3310 = 4'h5 == state ? _GEN_3027 : {{8'd0}, write_back_addr}; // @[d_cache.scala 76:18 42:34]
  wire  _GEN_3311 = 4'h5 == state ? _GEN_3028 : dirty_0_0; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3312 = 4'h5 == state ? _GEN_3029 : dirty_0_1; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3313 = 4'h5 == state ? _GEN_3030 : dirty_0_2; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3314 = 4'h5 == state ? _GEN_3031 : dirty_0_3; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3315 = 4'h5 == state ? _GEN_3032 : dirty_0_4; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3316 = 4'h5 == state ? _GEN_3033 : dirty_0_5; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3317 = 4'h5 == state ? _GEN_3034 : dirty_0_6; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3318 = 4'h5 == state ? _GEN_3035 : dirty_0_7; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3319 = 4'h5 == state ? _GEN_3036 : dirty_0_8; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3320 = 4'h5 == state ? _GEN_3037 : dirty_0_9; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3321 = 4'h5 == state ? _GEN_3038 : dirty_0_10; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3322 = 4'h5 == state ? _GEN_3039 : dirty_0_11; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3323 = 4'h5 == state ? _GEN_3040 : dirty_0_12; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3324 = 4'h5 == state ? _GEN_3041 : dirty_0_13; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3325 = 4'h5 == state ? _GEN_3042 : dirty_0_14; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3326 = 4'h5 == state ? _GEN_3043 : dirty_0_15; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3359 = 4'h5 == state ? _GEN_3076 : dirty_3_0; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3360 = 4'h5 == state ? _GEN_3077 : dirty_3_1; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3361 = 4'h5 == state ? _GEN_3078 : dirty_3_2; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3362 = 4'h5 == state ? _GEN_3079 : dirty_3_3; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3363 = 4'h5 == state ? _GEN_3080 : dirty_3_4; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3364 = 4'h5 == state ? _GEN_3081 : dirty_3_5; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3365 = 4'h5 == state ? _GEN_3082 : dirty_3_6; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3366 = 4'h5 == state ? _GEN_3083 : dirty_3_7; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3367 = 4'h5 == state ? _GEN_3084 : dirty_3_8; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3368 = 4'h5 == state ? _GEN_3085 : dirty_3_9; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3369 = 4'h5 == state ? _GEN_3086 : dirty_3_10; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3370 = 4'h5 == state ? _GEN_3087 : dirty_3_11; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3371 = 4'h5 == state ? _GEN_3088 : dirty_3_12; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3372 = 4'h5 == state ? _GEN_3089 : dirty_3_13; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3373 = 4'h5 == state ? _GEN_3090 : dirty_3_14; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3374 = 4'h5 == state ? _GEN_3091 : dirty_3_15; // @[d_cache.scala 76:18 35:26]
  wire [3:0] _GEN_3375 = 4'h4 == state ? _GEN_658 : _GEN_3100; // @[d_cache.scala 76:18]
  wire [127:0] _GEN_3376 = 4'h4 == state ? ram_0_0 : _GEN_3101; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3377 = 4'h4 == state ? ram_0_1 : _GEN_3102; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3378 = 4'h4 == state ? ram_0_2 : _GEN_3103; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3379 = 4'h4 == state ? ram_0_3 : _GEN_3104; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3380 = 4'h4 == state ? ram_0_4 : _GEN_3105; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3381 = 4'h4 == state ? ram_0_5 : _GEN_3106; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3382 = 4'h4 == state ? ram_0_6 : _GEN_3107; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3383 = 4'h4 == state ? ram_0_7 : _GEN_3108; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3384 = 4'h4 == state ? ram_0_8 : _GEN_3109; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3385 = 4'h4 == state ? ram_0_9 : _GEN_3110; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3386 = 4'h4 == state ? ram_0_10 : _GEN_3111; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3387 = 4'h4 == state ? ram_0_11 : _GEN_3112; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3388 = 4'h4 == state ? ram_0_12 : _GEN_3113; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3389 = 4'h4 == state ? ram_0_13 : _GEN_3114; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3390 = 4'h4 == state ? ram_0_14 : _GEN_3115; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3391 = 4'h4 == state ? ram_0_15 : _GEN_3116; // @[d_cache.scala 76:18 19:24]
  wire [31:0] _GEN_3392 = 4'h4 == state ? tag_0_0 : _GEN_3117; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3393 = 4'h4 == state ? tag_0_1 : _GEN_3118; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3394 = 4'h4 == state ? tag_0_2 : _GEN_3119; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3395 = 4'h4 == state ? tag_0_3 : _GEN_3120; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3396 = 4'h4 == state ? tag_0_4 : _GEN_3121; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3397 = 4'h4 == state ? tag_0_5 : _GEN_3122; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3398 = 4'h4 == state ? tag_0_6 : _GEN_3123; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3399 = 4'h4 == state ? tag_0_7 : _GEN_3124; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3400 = 4'h4 == state ? tag_0_8 : _GEN_3125; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3401 = 4'h4 == state ? tag_0_9 : _GEN_3126; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3402 = 4'h4 == state ? tag_0_10 : _GEN_3127; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3403 = 4'h4 == state ? tag_0_11 : _GEN_3128; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3404 = 4'h4 == state ? tag_0_12 : _GEN_3129; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3405 = 4'h4 == state ? tag_0_13 : _GEN_3130; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3406 = 4'h4 == state ? tag_0_14 : _GEN_3131; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3407 = 4'h4 == state ? tag_0_15 : _GEN_3132; // @[d_cache.scala 76:18 24:24]
  wire  _GEN_3408 = 4'h4 == state ? valid_0_0 : _GEN_3133; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3409 = 4'h4 == state ? valid_0_1 : _GEN_3134; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3410 = 4'h4 == state ? valid_0_2 : _GEN_3135; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3411 = 4'h4 == state ? valid_0_3 : _GEN_3136; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3412 = 4'h4 == state ? valid_0_4 : _GEN_3137; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3413 = 4'h4 == state ? valid_0_5 : _GEN_3138; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3414 = 4'h4 == state ? valid_0_6 : _GEN_3139; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3415 = 4'h4 == state ? valid_0_7 : _GEN_3140; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3416 = 4'h4 == state ? valid_0_8 : _GEN_3141; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3417 = 4'h4 == state ? valid_0_9 : _GEN_3142; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3418 = 4'h4 == state ? valid_0_10 : _GEN_3143; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3419 = 4'h4 == state ? valid_0_11 : _GEN_3144; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3420 = 4'h4 == state ? valid_0_12 : _GEN_3145; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3421 = 4'h4 == state ? valid_0_13 : _GEN_3146; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3422 = 4'h4 == state ? valid_0_14 : _GEN_3147; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3423 = 4'h4 == state ? valid_0_15 : _GEN_3148; // @[d_cache.scala 76:18 28:26]
  wire [7:0] _GEN_3424 = 4'h4 == state ? quene_0 : _GEN_3149; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3425 = 4'h4 == state ? quene_1 : _GEN_3150; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3426 = 4'h4 == state ? quene_2 : _GEN_3151; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3427 = 4'h4 == state ? quene_3 : _GEN_3152; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3428 = 4'h4 == state ? quene_4 : _GEN_3153; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3429 = 4'h4 == state ? quene_5 : _GEN_3154; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3430 = 4'h4 == state ? quene_6 : _GEN_3155; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3431 = 4'h4 == state ? quene_7 : _GEN_3156; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3432 = 4'h4 == state ? quene_8 : _GEN_3157; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3433 = 4'h4 == state ? quene_9 : _GEN_3158; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3434 = 4'h4 == state ? quene_10 : _GEN_3159; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3435 = 4'h4 == state ? quene_11 : _GEN_3160; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3436 = 4'h4 == state ? quene_12 : _GEN_3161; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3437 = 4'h4 == state ? quene_13 : _GEN_3162; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3438 = 4'h4 == state ? quene_14 : _GEN_3163; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3439 = 4'h4 == state ? quene_15 : _GEN_3164; // @[d_cache.scala 76:18 49:24]
  wire [127:0] _GEN_3440 = 4'h4 == state ? ram_1_0 : _GEN_3165; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3441 = 4'h4 == state ? ram_1_1 : _GEN_3166; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3442 = 4'h4 == state ? ram_1_2 : _GEN_3167; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3443 = 4'h4 == state ? ram_1_3 : _GEN_3168; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3444 = 4'h4 == state ? ram_1_4 : _GEN_3169; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3445 = 4'h4 == state ? ram_1_5 : _GEN_3170; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3446 = 4'h4 == state ? ram_1_6 : _GEN_3171; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3447 = 4'h4 == state ? ram_1_7 : _GEN_3172; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3448 = 4'h4 == state ? ram_1_8 : _GEN_3173; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3449 = 4'h4 == state ? ram_1_9 : _GEN_3174; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3450 = 4'h4 == state ? ram_1_10 : _GEN_3175; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3451 = 4'h4 == state ? ram_1_11 : _GEN_3176; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3452 = 4'h4 == state ? ram_1_12 : _GEN_3177; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3453 = 4'h4 == state ? ram_1_13 : _GEN_3178; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3454 = 4'h4 == state ? ram_1_14 : _GEN_3179; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3455 = 4'h4 == state ? ram_1_15 : _GEN_3180; // @[d_cache.scala 76:18 20:24]
  wire [31:0] _GEN_3456 = 4'h4 == state ? tag_1_0 : _GEN_3181; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3457 = 4'h4 == state ? tag_1_1 : _GEN_3182; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3458 = 4'h4 == state ? tag_1_2 : _GEN_3183; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3459 = 4'h4 == state ? tag_1_3 : _GEN_3184; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3460 = 4'h4 == state ? tag_1_4 : _GEN_3185; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3461 = 4'h4 == state ? tag_1_5 : _GEN_3186; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3462 = 4'h4 == state ? tag_1_6 : _GEN_3187; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3463 = 4'h4 == state ? tag_1_7 : _GEN_3188; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3464 = 4'h4 == state ? tag_1_8 : _GEN_3189; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3465 = 4'h4 == state ? tag_1_9 : _GEN_3190; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3466 = 4'h4 == state ? tag_1_10 : _GEN_3191; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3467 = 4'h4 == state ? tag_1_11 : _GEN_3192; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3468 = 4'h4 == state ? tag_1_12 : _GEN_3193; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3469 = 4'h4 == state ? tag_1_13 : _GEN_3194; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3470 = 4'h4 == state ? tag_1_14 : _GEN_3195; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3471 = 4'h4 == state ? tag_1_15 : _GEN_3196; // @[d_cache.scala 76:18 25:24]
  wire  _GEN_3472 = 4'h4 == state ? valid_1_0 : _GEN_3197; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3473 = 4'h4 == state ? valid_1_1 : _GEN_3198; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3474 = 4'h4 == state ? valid_1_2 : _GEN_3199; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3475 = 4'h4 == state ? valid_1_3 : _GEN_3200; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3476 = 4'h4 == state ? valid_1_4 : _GEN_3201; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3477 = 4'h4 == state ? valid_1_5 : _GEN_3202; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3478 = 4'h4 == state ? valid_1_6 : _GEN_3203; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3479 = 4'h4 == state ? valid_1_7 : _GEN_3204; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3480 = 4'h4 == state ? valid_1_8 : _GEN_3205; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3481 = 4'h4 == state ? valid_1_9 : _GEN_3206; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3482 = 4'h4 == state ? valid_1_10 : _GEN_3207; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3483 = 4'h4 == state ? valid_1_11 : _GEN_3208; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3484 = 4'h4 == state ? valid_1_12 : _GEN_3209; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3485 = 4'h4 == state ? valid_1_13 : _GEN_3210; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3486 = 4'h4 == state ? valid_1_14 : _GEN_3211; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3487 = 4'h4 == state ? valid_1_15 : _GEN_3212; // @[d_cache.scala 76:18 29:26]
  wire [127:0] _GEN_3488 = 4'h4 == state ? ram_2_0 : _GEN_3213; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3489 = 4'h4 == state ? ram_2_1 : _GEN_3214; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3490 = 4'h4 == state ? ram_2_2 : _GEN_3215; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3491 = 4'h4 == state ? ram_2_3 : _GEN_3216; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3492 = 4'h4 == state ? ram_2_4 : _GEN_3217; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3493 = 4'h4 == state ? ram_2_5 : _GEN_3218; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3494 = 4'h4 == state ? ram_2_6 : _GEN_3219; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3495 = 4'h4 == state ? ram_2_7 : _GEN_3220; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3496 = 4'h4 == state ? ram_2_8 : _GEN_3221; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3497 = 4'h4 == state ? ram_2_9 : _GEN_3222; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3498 = 4'h4 == state ? ram_2_10 : _GEN_3223; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3499 = 4'h4 == state ? ram_2_11 : _GEN_3224; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3500 = 4'h4 == state ? ram_2_12 : _GEN_3225; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3501 = 4'h4 == state ? ram_2_13 : _GEN_3226; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3502 = 4'h4 == state ? ram_2_14 : _GEN_3227; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3503 = 4'h4 == state ? ram_2_15 : _GEN_3228; // @[d_cache.scala 76:18 21:24]
  wire [31:0] _GEN_3504 = 4'h4 == state ? tag_2_0 : _GEN_3229; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3505 = 4'h4 == state ? tag_2_1 : _GEN_3230; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3506 = 4'h4 == state ? tag_2_2 : _GEN_3231; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3507 = 4'h4 == state ? tag_2_3 : _GEN_3232; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3508 = 4'h4 == state ? tag_2_4 : _GEN_3233; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3509 = 4'h4 == state ? tag_2_5 : _GEN_3234; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3510 = 4'h4 == state ? tag_2_6 : _GEN_3235; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3511 = 4'h4 == state ? tag_2_7 : _GEN_3236; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3512 = 4'h4 == state ? tag_2_8 : _GEN_3237; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3513 = 4'h4 == state ? tag_2_9 : _GEN_3238; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3514 = 4'h4 == state ? tag_2_10 : _GEN_3239; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3515 = 4'h4 == state ? tag_2_11 : _GEN_3240; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3516 = 4'h4 == state ? tag_2_12 : _GEN_3241; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3517 = 4'h4 == state ? tag_2_13 : _GEN_3242; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3518 = 4'h4 == state ? tag_2_14 : _GEN_3243; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3519 = 4'h4 == state ? tag_2_15 : _GEN_3244; // @[d_cache.scala 76:18 26:24]
  wire  _GEN_3520 = 4'h4 == state ? valid_2_0 : _GEN_3245; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3521 = 4'h4 == state ? valid_2_1 : _GEN_3246; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3522 = 4'h4 == state ? valid_2_2 : _GEN_3247; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3523 = 4'h4 == state ? valid_2_3 : _GEN_3248; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3524 = 4'h4 == state ? valid_2_4 : _GEN_3249; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3525 = 4'h4 == state ? valid_2_5 : _GEN_3250; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3526 = 4'h4 == state ? valid_2_6 : _GEN_3251; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3527 = 4'h4 == state ? valid_2_7 : _GEN_3252; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3528 = 4'h4 == state ? valid_2_8 : _GEN_3253; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3529 = 4'h4 == state ? valid_2_9 : _GEN_3254; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3530 = 4'h4 == state ? valid_2_10 : _GEN_3255; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3531 = 4'h4 == state ? valid_2_11 : _GEN_3256; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3532 = 4'h4 == state ? valid_2_12 : _GEN_3257; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3533 = 4'h4 == state ? valid_2_13 : _GEN_3258; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3534 = 4'h4 == state ? valid_2_14 : _GEN_3259; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3535 = 4'h4 == state ? valid_2_15 : _GEN_3260; // @[d_cache.scala 76:18 30:26]
  wire [127:0] _GEN_3536 = 4'h4 == state ? ram_3_0 : _GEN_3261; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3537 = 4'h4 == state ? ram_3_1 : _GEN_3262; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3538 = 4'h4 == state ? ram_3_2 : _GEN_3263; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3539 = 4'h4 == state ? ram_3_3 : _GEN_3264; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3540 = 4'h4 == state ? ram_3_4 : _GEN_3265; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3541 = 4'h4 == state ? ram_3_5 : _GEN_3266; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3542 = 4'h4 == state ? ram_3_6 : _GEN_3267; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3543 = 4'h4 == state ? ram_3_7 : _GEN_3268; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3544 = 4'h4 == state ? ram_3_8 : _GEN_3269; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3545 = 4'h4 == state ? ram_3_9 : _GEN_3270; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3546 = 4'h4 == state ? ram_3_10 : _GEN_3271; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3547 = 4'h4 == state ? ram_3_11 : _GEN_3272; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3548 = 4'h4 == state ? ram_3_12 : _GEN_3273; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3549 = 4'h4 == state ? ram_3_13 : _GEN_3274; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3550 = 4'h4 == state ? ram_3_14 : _GEN_3275; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3551 = 4'h4 == state ? ram_3_15 : _GEN_3276; // @[d_cache.scala 76:18 22:24]
  wire [31:0] _GEN_3552 = 4'h4 == state ? tag_3_0 : _GEN_3277; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3553 = 4'h4 == state ? tag_3_1 : _GEN_3278; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3554 = 4'h4 == state ? tag_3_2 : _GEN_3279; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3555 = 4'h4 == state ? tag_3_3 : _GEN_3280; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3556 = 4'h4 == state ? tag_3_4 : _GEN_3281; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3557 = 4'h4 == state ? tag_3_5 : _GEN_3282; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3558 = 4'h4 == state ? tag_3_6 : _GEN_3283; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3559 = 4'h4 == state ? tag_3_7 : _GEN_3284; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3560 = 4'h4 == state ? tag_3_8 : _GEN_3285; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3561 = 4'h4 == state ? tag_3_9 : _GEN_3286; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3562 = 4'h4 == state ? tag_3_10 : _GEN_3287; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3563 = 4'h4 == state ? tag_3_11 : _GEN_3288; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3564 = 4'h4 == state ? tag_3_12 : _GEN_3289; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3565 = 4'h4 == state ? tag_3_13 : _GEN_3290; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3566 = 4'h4 == state ? tag_3_14 : _GEN_3291; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3567 = 4'h4 == state ? tag_3_15 : _GEN_3292; // @[d_cache.scala 76:18 27:24]
  wire  _GEN_3568 = 4'h4 == state ? valid_3_0 : _GEN_3293; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3569 = 4'h4 == state ? valid_3_1 : _GEN_3294; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3570 = 4'h4 == state ? valid_3_2 : _GEN_3295; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3571 = 4'h4 == state ? valid_3_3 : _GEN_3296; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3572 = 4'h4 == state ? valid_3_4 : _GEN_3297; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3573 = 4'h4 == state ? valid_3_5 : _GEN_3298; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3574 = 4'h4 == state ? valid_3_6 : _GEN_3299; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3575 = 4'h4 == state ? valid_3_7 : _GEN_3300; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3576 = 4'h4 == state ? valid_3_8 : _GEN_3301; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3577 = 4'h4 == state ? valid_3_9 : _GEN_3302; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3578 = 4'h4 == state ? valid_3_10 : _GEN_3303; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3579 = 4'h4 == state ? valid_3_11 : _GEN_3304; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3580 = 4'h4 == state ? valid_3_12 : _GEN_3305; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3581 = 4'h4 == state ? valid_3_13 : _GEN_3306; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3582 = 4'h4 == state ? valid_3_14 : _GEN_3307; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3583 = 4'h4 == state ? valid_3_15 : _GEN_3308; // @[d_cache.scala 76:18 31:26]
  wire [127:0] _GEN_3584 = 4'h4 == state ? write_back_data : _GEN_3309; // @[d_cache.scala 76:18 41:34]
  wire [39:0] _GEN_3585 = 4'h4 == state ? {{8'd0}, write_back_addr} : _GEN_3310; // @[d_cache.scala 76:18 42:34]
  wire  _GEN_3586 = 4'h4 == state ? dirty_0_0 : _GEN_3311; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3587 = 4'h4 == state ? dirty_0_1 : _GEN_3312; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3588 = 4'h4 == state ? dirty_0_2 : _GEN_3313; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3589 = 4'h4 == state ? dirty_0_3 : _GEN_3314; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3590 = 4'h4 == state ? dirty_0_4 : _GEN_3315; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3591 = 4'h4 == state ? dirty_0_5 : _GEN_3316; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3592 = 4'h4 == state ? dirty_0_6 : _GEN_3317; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3593 = 4'h4 == state ? dirty_0_7 : _GEN_3318; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3594 = 4'h4 == state ? dirty_0_8 : _GEN_3319; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3595 = 4'h4 == state ? dirty_0_9 : _GEN_3320; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3596 = 4'h4 == state ? dirty_0_10 : _GEN_3321; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3597 = 4'h4 == state ? dirty_0_11 : _GEN_3322; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3598 = 4'h4 == state ? dirty_0_12 : _GEN_3323; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3599 = 4'h4 == state ? dirty_0_13 : _GEN_3324; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3600 = 4'h4 == state ? dirty_0_14 : _GEN_3325; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3601 = 4'h4 == state ? dirty_0_15 : _GEN_3326; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3634 = 4'h4 == state ? dirty_3_0 : _GEN_3359; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3635 = 4'h4 == state ? dirty_3_1 : _GEN_3360; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3636 = 4'h4 == state ? dirty_3_2 : _GEN_3361; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3637 = 4'h4 == state ? dirty_3_3 : _GEN_3362; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3638 = 4'h4 == state ? dirty_3_4 : _GEN_3363; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3639 = 4'h4 == state ? dirty_3_5 : _GEN_3364; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3640 = 4'h4 == state ? dirty_3_6 : _GEN_3365; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3641 = 4'h4 == state ? dirty_3_7 : _GEN_3366; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3642 = 4'h4 == state ? dirty_3_8 : _GEN_3367; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3643 = 4'h4 == state ? dirty_3_9 : _GEN_3368; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3644 = 4'h4 == state ? dirty_3_10 : _GEN_3369; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3645 = 4'h4 == state ? dirty_3_11 : _GEN_3370; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3646 = 4'h4 == state ? dirty_3_12 : _GEN_3371; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3647 = 4'h4 == state ? dirty_3_13 : _GEN_3372; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3648 = 4'h4 == state ? dirty_3_14 : _GEN_3373; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3649 = 4'h4 == state ? dirty_3_15 : _GEN_3374; // @[d_cache.scala 76:18 35:26]
  wire [63:0] _GEN_3650 = 4'h3 == state ? _GEN_654 : receive_data_0; // @[d_cache.scala 76:18 47:31]
  wire [63:0] _GEN_3651 = 4'h3 == state ? _GEN_655 : receive_data_1; // @[d_cache.scala 76:18 47:31]
  wire [2:0] _GEN_3652 = 4'h3 == state ? _GEN_656 : receive_num; // @[d_cache.scala 76:18 48:30]
  wire [3:0] _GEN_3653 = 4'h3 == state ? _GEN_657 : _GEN_3375; // @[d_cache.scala 76:18]
  wire [127:0] _GEN_3654 = 4'h3 == state ? ram_0_0 : _GEN_3376; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3655 = 4'h3 == state ? ram_0_1 : _GEN_3377; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3656 = 4'h3 == state ? ram_0_2 : _GEN_3378; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3657 = 4'h3 == state ? ram_0_3 : _GEN_3379; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3658 = 4'h3 == state ? ram_0_4 : _GEN_3380; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3659 = 4'h3 == state ? ram_0_5 : _GEN_3381; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3660 = 4'h3 == state ? ram_0_6 : _GEN_3382; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3661 = 4'h3 == state ? ram_0_7 : _GEN_3383; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3662 = 4'h3 == state ? ram_0_8 : _GEN_3384; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3663 = 4'h3 == state ? ram_0_9 : _GEN_3385; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3664 = 4'h3 == state ? ram_0_10 : _GEN_3386; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3665 = 4'h3 == state ? ram_0_11 : _GEN_3387; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3666 = 4'h3 == state ? ram_0_12 : _GEN_3388; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3667 = 4'h3 == state ? ram_0_13 : _GEN_3389; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3668 = 4'h3 == state ? ram_0_14 : _GEN_3390; // @[d_cache.scala 76:18 19:24]
  wire [127:0] _GEN_3669 = 4'h3 == state ? ram_0_15 : _GEN_3391; // @[d_cache.scala 76:18 19:24]
  wire [31:0] _GEN_3670 = 4'h3 == state ? tag_0_0 : _GEN_3392; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3671 = 4'h3 == state ? tag_0_1 : _GEN_3393; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3672 = 4'h3 == state ? tag_0_2 : _GEN_3394; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3673 = 4'h3 == state ? tag_0_3 : _GEN_3395; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3674 = 4'h3 == state ? tag_0_4 : _GEN_3396; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3675 = 4'h3 == state ? tag_0_5 : _GEN_3397; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3676 = 4'h3 == state ? tag_0_6 : _GEN_3398; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3677 = 4'h3 == state ? tag_0_7 : _GEN_3399; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3678 = 4'h3 == state ? tag_0_8 : _GEN_3400; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3679 = 4'h3 == state ? tag_0_9 : _GEN_3401; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3680 = 4'h3 == state ? tag_0_10 : _GEN_3402; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3681 = 4'h3 == state ? tag_0_11 : _GEN_3403; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3682 = 4'h3 == state ? tag_0_12 : _GEN_3404; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3683 = 4'h3 == state ? tag_0_13 : _GEN_3405; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3684 = 4'h3 == state ? tag_0_14 : _GEN_3406; // @[d_cache.scala 76:18 24:24]
  wire [31:0] _GEN_3685 = 4'h3 == state ? tag_0_15 : _GEN_3407; // @[d_cache.scala 76:18 24:24]
  wire  _GEN_3686 = 4'h3 == state ? valid_0_0 : _GEN_3408; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3687 = 4'h3 == state ? valid_0_1 : _GEN_3409; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3688 = 4'h3 == state ? valid_0_2 : _GEN_3410; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3689 = 4'h3 == state ? valid_0_3 : _GEN_3411; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3690 = 4'h3 == state ? valid_0_4 : _GEN_3412; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3691 = 4'h3 == state ? valid_0_5 : _GEN_3413; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3692 = 4'h3 == state ? valid_0_6 : _GEN_3414; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3693 = 4'h3 == state ? valid_0_7 : _GEN_3415; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3694 = 4'h3 == state ? valid_0_8 : _GEN_3416; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3695 = 4'h3 == state ? valid_0_9 : _GEN_3417; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3696 = 4'h3 == state ? valid_0_10 : _GEN_3418; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3697 = 4'h3 == state ? valid_0_11 : _GEN_3419; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3698 = 4'h3 == state ? valid_0_12 : _GEN_3420; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3699 = 4'h3 == state ? valid_0_13 : _GEN_3421; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3700 = 4'h3 == state ? valid_0_14 : _GEN_3422; // @[d_cache.scala 76:18 28:26]
  wire  _GEN_3701 = 4'h3 == state ? valid_0_15 : _GEN_3423; // @[d_cache.scala 76:18 28:26]
  wire [7:0] _GEN_3702 = 4'h3 == state ? quene_0 : _GEN_3424; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3703 = 4'h3 == state ? quene_1 : _GEN_3425; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3704 = 4'h3 == state ? quene_2 : _GEN_3426; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3705 = 4'h3 == state ? quene_3 : _GEN_3427; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3706 = 4'h3 == state ? quene_4 : _GEN_3428; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3707 = 4'h3 == state ? quene_5 : _GEN_3429; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3708 = 4'h3 == state ? quene_6 : _GEN_3430; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3709 = 4'h3 == state ? quene_7 : _GEN_3431; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3710 = 4'h3 == state ? quene_8 : _GEN_3432; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3711 = 4'h3 == state ? quene_9 : _GEN_3433; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3712 = 4'h3 == state ? quene_10 : _GEN_3434; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3713 = 4'h3 == state ? quene_11 : _GEN_3435; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3714 = 4'h3 == state ? quene_12 : _GEN_3436; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3715 = 4'h3 == state ? quene_13 : _GEN_3437; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3716 = 4'h3 == state ? quene_14 : _GEN_3438; // @[d_cache.scala 76:18 49:24]
  wire [7:0] _GEN_3717 = 4'h3 == state ? quene_15 : _GEN_3439; // @[d_cache.scala 76:18 49:24]
  wire [127:0] _GEN_3718 = 4'h3 == state ? ram_1_0 : _GEN_3440; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3719 = 4'h3 == state ? ram_1_1 : _GEN_3441; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3720 = 4'h3 == state ? ram_1_2 : _GEN_3442; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3721 = 4'h3 == state ? ram_1_3 : _GEN_3443; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3722 = 4'h3 == state ? ram_1_4 : _GEN_3444; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3723 = 4'h3 == state ? ram_1_5 : _GEN_3445; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3724 = 4'h3 == state ? ram_1_6 : _GEN_3446; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3725 = 4'h3 == state ? ram_1_7 : _GEN_3447; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3726 = 4'h3 == state ? ram_1_8 : _GEN_3448; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3727 = 4'h3 == state ? ram_1_9 : _GEN_3449; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3728 = 4'h3 == state ? ram_1_10 : _GEN_3450; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3729 = 4'h3 == state ? ram_1_11 : _GEN_3451; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3730 = 4'h3 == state ? ram_1_12 : _GEN_3452; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3731 = 4'h3 == state ? ram_1_13 : _GEN_3453; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3732 = 4'h3 == state ? ram_1_14 : _GEN_3454; // @[d_cache.scala 76:18 20:24]
  wire [127:0] _GEN_3733 = 4'h3 == state ? ram_1_15 : _GEN_3455; // @[d_cache.scala 76:18 20:24]
  wire [31:0] _GEN_3734 = 4'h3 == state ? tag_1_0 : _GEN_3456; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3735 = 4'h3 == state ? tag_1_1 : _GEN_3457; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3736 = 4'h3 == state ? tag_1_2 : _GEN_3458; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3737 = 4'h3 == state ? tag_1_3 : _GEN_3459; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3738 = 4'h3 == state ? tag_1_4 : _GEN_3460; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3739 = 4'h3 == state ? tag_1_5 : _GEN_3461; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3740 = 4'h3 == state ? tag_1_6 : _GEN_3462; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3741 = 4'h3 == state ? tag_1_7 : _GEN_3463; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3742 = 4'h3 == state ? tag_1_8 : _GEN_3464; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3743 = 4'h3 == state ? tag_1_9 : _GEN_3465; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3744 = 4'h3 == state ? tag_1_10 : _GEN_3466; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3745 = 4'h3 == state ? tag_1_11 : _GEN_3467; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3746 = 4'h3 == state ? tag_1_12 : _GEN_3468; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3747 = 4'h3 == state ? tag_1_13 : _GEN_3469; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3748 = 4'h3 == state ? tag_1_14 : _GEN_3470; // @[d_cache.scala 76:18 25:24]
  wire [31:0] _GEN_3749 = 4'h3 == state ? tag_1_15 : _GEN_3471; // @[d_cache.scala 76:18 25:24]
  wire  _GEN_3750 = 4'h3 == state ? valid_1_0 : _GEN_3472; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3751 = 4'h3 == state ? valid_1_1 : _GEN_3473; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3752 = 4'h3 == state ? valid_1_2 : _GEN_3474; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3753 = 4'h3 == state ? valid_1_3 : _GEN_3475; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3754 = 4'h3 == state ? valid_1_4 : _GEN_3476; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3755 = 4'h3 == state ? valid_1_5 : _GEN_3477; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3756 = 4'h3 == state ? valid_1_6 : _GEN_3478; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3757 = 4'h3 == state ? valid_1_7 : _GEN_3479; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3758 = 4'h3 == state ? valid_1_8 : _GEN_3480; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3759 = 4'h3 == state ? valid_1_9 : _GEN_3481; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3760 = 4'h3 == state ? valid_1_10 : _GEN_3482; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3761 = 4'h3 == state ? valid_1_11 : _GEN_3483; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3762 = 4'h3 == state ? valid_1_12 : _GEN_3484; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3763 = 4'h3 == state ? valid_1_13 : _GEN_3485; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3764 = 4'h3 == state ? valid_1_14 : _GEN_3486; // @[d_cache.scala 76:18 29:26]
  wire  _GEN_3765 = 4'h3 == state ? valid_1_15 : _GEN_3487; // @[d_cache.scala 76:18 29:26]
  wire [127:0] _GEN_3766 = 4'h3 == state ? ram_2_0 : _GEN_3488; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3767 = 4'h3 == state ? ram_2_1 : _GEN_3489; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3768 = 4'h3 == state ? ram_2_2 : _GEN_3490; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3769 = 4'h3 == state ? ram_2_3 : _GEN_3491; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3770 = 4'h3 == state ? ram_2_4 : _GEN_3492; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3771 = 4'h3 == state ? ram_2_5 : _GEN_3493; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3772 = 4'h3 == state ? ram_2_6 : _GEN_3494; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3773 = 4'h3 == state ? ram_2_7 : _GEN_3495; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3774 = 4'h3 == state ? ram_2_8 : _GEN_3496; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3775 = 4'h3 == state ? ram_2_9 : _GEN_3497; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3776 = 4'h3 == state ? ram_2_10 : _GEN_3498; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3777 = 4'h3 == state ? ram_2_11 : _GEN_3499; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3778 = 4'h3 == state ? ram_2_12 : _GEN_3500; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3779 = 4'h3 == state ? ram_2_13 : _GEN_3501; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3780 = 4'h3 == state ? ram_2_14 : _GEN_3502; // @[d_cache.scala 76:18 21:24]
  wire [127:0] _GEN_3781 = 4'h3 == state ? ram_2_15 : _GEN_3503; // @[d_cache.scala 76:18 21:24]
  wire [31:0] _GEN_3782 = 4'h3 == state ? tag_2_0 : _GEN_3504; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3783 = 4'h3 == state ? tag_2_1 : _GEN_3505; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3784 = 4'h3 == state ? tag_2_2 : _GEN_3506; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3785 = 4'h3 == state ? tag_2_3 : _GEN_3507; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3786 = 4'h3 == state ? tag_2_4 : _GEN_3508; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3787 = 4'h3 == state ? tag_2_5 : _GEN_3509; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3788 = 4'h3 == state ? tag_2_6 : _GEN_3510; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3789 = 4'h3 == state ? tag_2_7 : _GEN_3511; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3790 = 4'h3 == state ? tag_2_8 : _GEN_3512; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3791 = 4'h3 == state ? tag_2_9 : _GEN_3513; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3792 = 4'h3 == state ? tag_2_10 : _GEN_3514; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3793 = 4'h3 == state ? tag_2_11 : _GEN_3515; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3794 = 4'h3 == state ? tag_2_12 : _GEN_3516; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3795 = 4'h3 == state ? tag_2_13 : _GEN_3517; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3796 = 4'h3 == state ? tag_2_14 : _GEN_3518; // @[d_cache.scala 76:18 26:24]
  wire [31:0] _GEN_3797 = 4'h3 == state ? tag_2_15 : _GEN_3519; // @[d_cache.scala 76:18 26:24]
  wire  _GEN_3798 = 4'h3 == state ? valid_2_0 : _GEN_3520; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3799 = 4'h3 == state ? valid_2_1 : _GEN_3521; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3800 = 4'h3 == state ? valid_2_2 : _GEN_3522; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3801 = 4'h3 == state ? valid_2_3 : _GEN_3523; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3802 = 4'h3 == state ? valid_2_4 : _GEN_3524; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3803 = 4'h3 == state ? valid_2_5 : _GEN_3525; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3804 = 4'h3 == state ? valid_2_6 : _GEN_3526; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3805 = 4'h3 == state ? valid_2_7 : _GEN_3527; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3806 = 4'h3 == state ? valid_2_8 : _GEN_3528; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3807 = 4'h3 == state ? valid_2_9 : _GEN_3529; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3808 = 4'h3 == state ? valid_2_10 : _GEN_3530; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3809 = 4'h3 == state ? valid_2_11 : _GEN_3531; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3810 = 4'h3 == state ? valid_2_12 : _GEN_3532; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3811 = 4'h3 == state ? valid_2_13 : _GEN_3533; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3812 = 4'h3 == state ? valid_2_14 : _GEN_3534; // @[d_cache.scala 76:18 30:26]
  wire  _GEN_3813 = 4'h3 == state ? valid_2_15 : _GEN_3535; // @[d_cache.scala 76:18 30:26]
  wire [127:0] _GEN_3814 = 4'h3 == state ? ram_3_0 : _GEN_3536; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3815 = 4'h3 == state ? ram_3_1 : _GEN_3537; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3816 = 4'h3 == state ? ram_3_2 : _GEN_3538; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3817 = 4'h3 == state ? ram_3_3 : _GEN_3539; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3818 = 4'h3 == state ? ram_3_4 : _GEN_3540; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3819 = 4'h3 == state ? ram_3_5 : _GEN_3541; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3820 = 4'h3 == state ? ram_3_6 : _GEN_3542; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3821 = 4'h3 == state ? ram_3_7 : _GEN_3543; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3822 = 4'h3 == state ? ram_3_8 : _GEN_3544; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3823 = 4'h3 == state ? ram_3_9 : _GEN_3545; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3824 = 4'h3 == state ? ram_3_10 : _GEN_3546; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3825 = 4'h3 == state ? ram_3_11 : _GEN_3547; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3826 = 4'h3 == state ? ram_3_12 : _GEN_3548; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3827 = 4'h3 == state ? ram_3_13 : _GEN_3549; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3828 = 4'h3 == state ? ram_3_14 : _GEN_3550; // @[d_cache.scala 76:18 22:24]
  wire [127:0] _GEN_3829 = 4'h3 == state ? ram_3_15 : _GEN_3551; // @[d_cache.scala 76:18 22:24]
  wire [31:0] _GEN_3830 = 4'h3 == state ? tag_3_0 : _GEN_3552; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3831 = 4'h3 == state ? tag_3_1 : _GEN_3553; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3832 = 4'h3 == state ? tag_3_2 : _GEN_3554; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3833 = 4'h3 == state ? tag_3_3 : _GEN_3555; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3834 = 4'h3 == state ? tag_3_4 : _GEN_3556; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3835 = 4'h3 == state ? tag_3_5 : _GEN_3557; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3836 = 4'h3 == state ? tag_3_6 : _GEN_3558; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3837 = 4'h3 == state ? tag_3_7 : _GEN_3559; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3838 = 4'h3 == state ? tag_3_8 : _GEN_3560; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3839 = 4'h3 == state ? tag_3_9 : _GEN_3561; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3840 = 4'h3 == state ? tag_3_10 : _GEN_3562; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3841 = 4'h3 == state ? tag_3_11 : _GEN_3563; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3842 = 4'h3 == state ? tag_3_12 : _GEN_3564; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3843 = 4'h3 == state ? tag_3_13 : _GEN_3565; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3844 = 4'h3 == state ? tag_3_14 : _GEN_3566; // @[d_cache.scala 76:18 27:24]
  wire [31:0] _GEN_3845 = 4'h3 == state ? tag_3_15 : _GEN_3567; // @[d_cache.scala 76:18 27:24]
  wire  _GEN_3846 = 4'h3 == state ? valid_3_0 : _GEN_3568; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3847 = 4'h3 == state ? valid_3_1 : _GEN_3569; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3848 = 4'h3 == state ? valid_3_2 : _GEN_3570; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3849 = 4'h3 == state ? valid_3_3 : _GEN_3571; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3850 = 4'h3 == state ? valid_3_4 : _GEN_3572; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3851 = 4'h3 == state ? valid_3_5 : _GEN_3573; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3852 = 4'h3 == state ? valid_3_6 : _GEN_3574; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3853 = 4'h3 == state ? valid_3_7 : _GEN_3575; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3854 = 4'h3 == state ? valid_3_8 : _GEN_3576; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3855 = 4'h3 == state ? valid_3_9 : _GEN_3577; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3856 = 4'h3 == state ? valid_3_10 : _GEN_3578; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3857 = 4'h3 == state ? valid_3_11 : _GEN_3579; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3858 = 4'h3 == state ? valid_3_12 : _GEN_3580; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3859 = 4'h3 == state ? valid_3_13 : _GEN_3581; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3860 = 4'h3 == state ? valid_3_14 : _GEN_3582; // @[d_cache.scala 76:18 31:26]
  wire  _GEN_3861 = 4'h3 == state ? valid_3_15 : _GEN_3583; // @[d_cache.scala 76:18 31:26]
  wire [127:0] _GEN_3862 = 4'h3 == state ? write_back_data : _GEN_3584; // @[d_cache.scala 76:18 41:34]
  wire [39:0] _GEN_3863 = 4'h3 == state ? {{8'd0}, write_back_addr} : _GEN_3585; // @[d_cache.scala 76:18 42:34]
  wire  _GEN_3864 = 4'h3 == state ? dirty_0_0 : _GEN_3586; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3865 = 4'h3 == state ? dirty_0_1 : _GEN_3587; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3866 = 4'h3 == state ? dirty_0_2 : _GEN_3588; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3867 = 4'h3 == state ? dirty_0_3 : _GEN_3589; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3868 = 4'h3 == state ? dirty_0_4 : _GEN_3590; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3869 = 4'h3 == state ? dirty_0_5 : _GEN_3591; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3870 = 4'h3 == state ? dirty_0_6 : _GEN_3592; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3871 = 4'h3 == state ? dirty_0_7 : _GEN_3593; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3872 = 4'h3 == state ? dirty_0_8 : _GEN_3594; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3873 = 4'h3 == state ? dirty_0_9 : _GEN_3595; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3874 = 4'h3 == state ? dirty_0_10 : _GEN_3596; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3875 = 4'h3 == state ? dirty_0_11 : _GEN_3597; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3876 = 4'h3 == state ? dirty_0_12 : _GEN_3598; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3877 = 4'h3 == state ? dirty_0_13 : _GEN_3599; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3878 = 4'h3 == state ? dirty_0_14 : _GEN_3600; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3879 = 4'h3 == state ? dirty_0_15 : _GEN_3601; // @[d_cache.scala 76:18 32:26]
  wire  _GEN_3912 = 4'h3 == state ? dirty_3_0 : _GEN_3634; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3913 = 4'h3 == state ? dirty_3_1 : _GEN_3635; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3914 = 4'h3 == state ? dirty_3_2 : _GEN_3636; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3915 = 4'h3 == state ? dirty_3_3 : _GEN_3637; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3916 = 4'h3 == state ? dirty_3_4 : _GEN_3638; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3917 = 4'h3 == state ? dirty_3_5 : _GEN_3639; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3918 = 4'h3 == state ? dirty_3_6 : _GEN_3640; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3919 = 4'h3 == state ? dirty_3_7 : _GEN_3641; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3920 = 4'h3 == state ? dirty_3_8 : _GEN_3642; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3921 = 4'h3 == state ? dirty_3_9 : _GEN_3643; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3922 = 4'h3 == state ? dirty_3_10 : _GEN_3644; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3923 = 4'h3 == state ? dirty_3_11 : _GEN_3645; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3924 = 4'h3 == state ? dirty_3_12 : _GEN_3646; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3925 = 4'h3 == state ? dirty_3_13 : _GEN_3647; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3926 = 4'h3 == state ? dirty_3_14 : _GEN_3648; // @[d_cache.scala 76:18 35:26]
  wire  _GEN_3927 = 4'h3 == state ? dirty_3_15 : _GEN_3649; // @[d_cache.scala 76:18 35:26]
  wire [39:0] _GEN_4205 = 4'h2 == state ? {{8'd0}, write_back_addr} : _GEN_3863; // @[d_cache.scala 76:18 42:34]
  wire [39:0] _GEN_4483 = 4'h1 == state ? {{8'd0}, write_back_addr} : _GEN_4205; // @[d_cache.scala 76:18 42:34]
  wire [39:0] _GEN_4761 = 4'h0 == state ? {{8'd0}, write_back_addr} : _GEN_4483; // @[d_cache.scala 76:18 42:34]
  wire [127:0] _io_to_lsu_rdata_T = _GEN_150 >> shift_bit; // @[d_cache.scala 262:54]
  wire [127:0] _io_to_lsu_rdata_T_1 = _GEN_198 >> shift_bit; // @[d_cache.scala 262:94]
  wire [127:0] _io_to_lsu_rdata_T_2 = _GEN_246 >> shift_bit; // @[d_cache.scala 262:134]
  wire [127:0] _io_to_lsu_rdata_T_3 = _GEN_294 >> shift_bit; // @[d_cache.scala 262:161]
  wire [127:0] _io_to_lsu_rdata_T_4 = way2_hit ? _io_to_lsu_rdata_T_2 : _io_to_lsu_rdata_T_3; // @[d_cache.scala 262:111]
  wire [127:0] _io_to_lsu_rdata_T_5 = way1_hit ? _io_to_lsu_rdata_T_1 : _io_to_lsu_rdata_T_4; // @[d_cache.scala 262:71]
  wire [127:0] _io_to_lsu_rdata_T_6 = way0_hit ? _io_to_lsu_rdata_T : _io_to_lsu_rdata_T_5; // @[d_cache.scala 262:31]
  wire [63:0] _GEN_1362 = {{32'd0}, io_from_lsu_araddr}; // @[d_cache.scala 303:49]
  wire [63:0] _io_to_axi_araddr_T = _GEN_1362 & 64'hfffffffffffffff0; // @[d_cache.scala 303:49]
  wire  _T_45 = state == 4'h0 & _T_5; // @[d_cache.scala 371:27]
  wire [63:0] _GEN_4763 = state == 4'h0 & _T_5 ? io_from_axi_rdata : 64'h0; // @[d_cache.scala 371:117 372:23 375:29]
  wire  _GEN_4765 = state == 4'h0 & _T_5 & io_from_axi_rvalid; // @[d_cache.scala 371:117 372:23 377:30]
  wire  _GEN_4768 = state == 4'h0 & _T_5 & io_from_axi_bvalid; // @[d_cache.scala 371:117 372:23 380:30]
  wire  _GEN_4773 = state == 4'h0 & _T_5 & io_from_lsu_arvalid; // @[d_cache.scala 371:117 373:23 382:31]
  wire [31:0] _GEN_4775 = state == 4'h0 & _T_5 ? io_from_lsu_awaddr : 32'h0; // @[d_cache.scala 371:117 373:23 388:30]
  wire  _GEN_4779 = state == 4'h0 & _T_5 & io_from_lsu_awvalid; // @[d_cache.scala 371:117 373:23 389:31]
  wire [63:0] _GEN_4780 = state == 4'h0 & _T_5 ? io_from_lsu_wdata : 64'h0; // @[d_cache.scala 371:117 373:23 393:29]
  wire [7:0] _GEN_4781 = state == 4'h0 & _T_5 ? io_from_lsu_wstrb : 8'h0; // @[d_cache.scala 371:117 373:23 394:29]
  wire  _GEN_4783 = state == 4'h0 & _T_5 & io_from_lsu_wvalid; // @[d_cache.scala 371:117 373:23 396:30]
  wire [63:0] _GEN_4786 = state == 4'h7 ? io_from_axi_rdata : _GEN_4763; // @[d_cache.scala 367:30 368:19]
  wire  _GEN_4788 = state == 4'h7 ? io_from_axi_rvalid : _GEN_4765; // @[d_cache.scala 367:30 368:19]
  wire  _GEN_4791 = state == 4'h7 ? io_from_axi_bvalid : _GEN_4768; // @[d_cache.scala 367:30 368:19]
  wire  _GEN_4796 = state == 4'h7 ? io_from_lsu_arvalid : _GEN_4773; // @[d_cache.scala 367:30 369:19]
  wire [31:0] _GEN_4798 = state == 4'h7 ? io_from_lsu_awaddr : _GEN_4775; // @[d_cache.scala 367:30 369:19]
  wire  _GEN_4802 = state == 4'h7 ? io_from_lsu_awvalid : _GEN_4779; // @[d_cache.scala 367:30 369:19]
  wire [63:0] _GEN_4803 = state == 4'h7 ? io_from_lsu_wdata : _GEN_4780; // @[d_cache.scala 367:30 369:19]
  wire [7:0] _GEN_4804 = state == 4'h7 ? io_from_lsu_wstrb : _GEN_4781; // @[d_cache.scala 367:30 369:19]
  wire  _GEN_4806 = state == 4'h7 ? io_from_lsu_wvalid : _GEN_4783; // @[d_cache.scala 367:30 369:19]
  wire  _GEN_4807 = state == 4'h7 | _T_45; // @[d_cache.scala 367:30 369:19]
  wire [63:0] _GEN_4808 = state == 4'h6 ? 64'h0 : _GEN_4786; // @[d_cache.scala 343:35 344:25]
  wire  _GEN_4810 = state == 4'h6 ? 1'h0 : _GEN_4788; // @[d_cache.scala 343:35 346:26]
  wire  _GEN_4813 = state == 4'h6 ? 1'h0 : _GEN_4791; // @[d_cache.scala 343:35 349:26]
  wire  _GEN_4815 = state == 4'h6 ? 1'h0 : _GEN_4796; // @[d_cache.scala 343:35 351:27]
  wire [31:0] _GEN_4816 = state == 4'h6 ? 32'h0 : io_from_lsu_araddr; // @[d_cache.scala 343:35 352:26]
  wire [7:0] _GEN_4817 = state == 4'h6 ? 8'h1 : 8'h0; // @[d_cache.scala 343:35 353:25]
  wire  _GEN_4820 = state == 4'h6 ? 1'h0 : 1'h1; // @[d_cache.scala 343:35 356:26]
  wire [31:0] _GEN_4821 = state == 4'h6 ? write_back_addr : _GEN_4798; // @[d_cache.scala 343:35 357:26]
  wire  _GEN_4822 = state == 4'h6 | _GEN_4802; // @[d_cache.scala 343:35 358:27]
  wire [63:0] _GEN_4826 = state == 4'h6 ? write_back_data[63:0] : _GEN_4803; // @[d_cache.scala 343:35 362:25]
  wire [7:0] _GEN_4827 = state == 4'h6 ? 8'hff : _GEN_4804; // @[d_cache.scala 343:35 363:25]
  wire  _GEN_4829 = state == 4'h6 | _GEN_4806; // @[d_cache.scala 343:35 365:26]
  wire  _GEN_4830 = state == 4'h6 | _GEN_4807; // @[d_cache.scala 343:35 366:26]
  wire [63:0] _GEN_4831 = state == 4'h4 | state == 4'h8 ? 64'h0 : _GEN_4808; // @[d_cache.scala 318:50 319:25]
  wire  _GEN_4833 = state == 4'h4 | state == 4'h8 ? 1'h0 : _GEN_4810; // @[d_cache.scala 318:50 321:26]
  wire  _GEN_4836 = state == 4'h4 | state == 4'h8 ? io_from_axi_bvalid : _GEN_4813; // @[d_cache.scala 318:50 324:26]
  wire  _GEN_4838 = state == 4'h4 | state == 4'h8 ? 1'h0 : _GEN_4815; // @[d_cache.scala 318:50 326:27]
  wire [31:0] _GEN_4839 = state == 4'h4 | state == 4'h8 ? 32'h0 : _GEN_4816; // @[d_cache.scala 318:50 327:26]
  wire [7:0] _GEN_4840 = state == 4'h4 | state == 4'h8 ? 8'h0 : _GEN_4817; // @[d_cache.scala 318:50 328:25]
  wire  _GEN_4843 = state == 4'h4 | state == 4'h8 | _GEN_4820; // @[d_cache.scala 318:50 331:26]
  wire [31:0] _GEN_4844 = state == 4'h4 | state == 4'h8 ? io_from_lsu_awaddr : _GEN_4821; // @[d_cache.scala 318:50 332:26]
  wire  _GEN_4845 = state == 4'h4 | state == 4'h8 ? io_from_lsu_awvalid : _GEN_4822; // @[d_cache.scala 318:50 333:27]
  wire [63:0] _GEN_4849 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wdata : _GEN_4826; // @[d_cache.scala 318:50 337:25]
  wire [7:0] _GEN_4850 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wstrb : _GEN_4827; // @[d_cache.scala 318:50 338:25]
  wire  _GEN_4852 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wvalid : _GEN_4829; // @[d_cache.scala 318:50 340:26]
  wire  _GEN_4853 = state == 4'h4 | state == 4'h8 | _GEN_4830; // @[d_cache.scala 318:50 341:26]
  wire [63:0] _GEN_4854 = state == 4'h3 ? 64'h0 : _GEN_4831; // @[d_cache.scala 294:31 295:25]
  wire  _GEN_4856 = state == 4'h3 ? 1'h0 : _GEN_4833; // @[d_cache.scala 294:31 297:26]
  wire  _GEN_4859 = state == 4'h3 ? 1'h0 : _GEN_4836; // @[d_cache.scala 294:31 300:26]
  wire  _GEN_4861 = state == 4'h3 | _GEN_4838; // @[d_cache.scala 294:31 302:27]
  wire [63:0] _GEN_4862 = state == 4'h3 ? _io_to_axi_araddr_T : {{32'd0}, _GEN_4839}; // @[d_cache.scala 294:31 303:26]
  wire [7:0] _GEN_4863 = state == 4'h3 ? 8'h1 : _GEN_4840; // @[d_cache.scala 294:31 304:25]
  wire  _GEN_4866 = state == 4'h3 | _GEN_4843; // @[d_cache.scala 294:31 307:26]
  wire [31:0] _GEN_4867 = state == 4'h3 ? 32'h0 : _GEN_4844; // @[d_cache.scala 294:31 308:26]
  wire  _GEN_4868 = state == 4'h3 ? 1'h0 : _GEN_4845; // @[d_cache.scala 294:31 309:27]
  wire [7:0] _GEN_4869 = state == 4'h3 ? 8'h0 : _GEN_4840; // @[d_cache.scala 294:31 310:25]
  wire [63:0] _GEN_4872 = state == 4'h3 ? 64'h0 : _GEN_4849; // @[d_cache.scala 294:31 313:25]
  wire [7:0] _GEN_4873 = state == 4'h3 ? 8'h0 : _GEN_4850; // @[d_cache.scala 294:31 314:25]
  wire  _GEN_4875 = state == 4'h3 ? 1'h0 : _GEN_4852; // @[d_cache.scala 294:31 316:26]
  wire  _GEN_4876 = state == 4'h3 ? 1'h0 : _GEN_4853; // @[d_cache.scala 294:31 317:26]
  wire  _GEN_4877 = state == 4'h2 ? 1'h0 : _GEN_4861; // @[d_cache.scala 270:33 271:27]
  wire [63:0] _GEN_4878 = state == 4'h2 ? {{32'd0}, io_from_lsu_araddr} : _GEN_4862; // @[d_cache.scala 270:33 272:26]
  wire [7:0] _GEN_4879 = state == 4'h2 ? 8'h0 : _GEN_4863; // @[d_cache.scala 270:33 273:25]
  wire  _GEN_4882 = state == 4'h2 ? 1'h0 : _GEN_4866; // @[d_cache.scala 270:33 276:26]
  wire [31:0] _GEN_4883 = state == 4'h2 ? 32'h0 : _GEN_4867; // @[d_cache.scala 270:33 277:26]
  wire  _GEN_4884 = state == 4'h2 ? 1'h0 : _GEN_4868; // @[d_cache.scala 270:33 278:27]
  wire [7:0] _GEN_4885 = state == 4'h2 ? 8'h0 : _GEN_4869; // @[d_cache.scala 270:33 279:25]
  wire [63:0] _GEN_4888 = state == 4'h2 ? 64'h0 : _GEN_4872; // @[d_cache.scala 270:33 282:25]
  wire [7:0] _GEN_4889 = state == 4'h2 ? 8'h0 : _GEN_4873; // @[d_cache.scala 270:33 283:25]
  wire  _GEN_4891 = state == 4'h2 ? 1'h0 : _GEN_4875; // @[d_cache.scala 270:33 285:26]
  wire  _GEN_4892 = state == 4'h2 ? 1'h0 : _GEN_4876; // @[d_cache.scala 270:33 286:26]
  wire [63:0] _GEN_4893 = state == 4'h2 ? 64'h0 : _GEN_4854; // @[d_cache.scala 270:33 287:25]
  wire  _GEN_4895 = state == 4'h2 ? 1'h0 : _GEN_4856; // @[d_cache.scala 270:33 289:26]
  wire  _GEN_4899 = state == 4'h2 ? _T_9 : _GEN_4859; // @[d_cache.scala 270:33 293:26]
  wire [63:0] _GEN_4901 = state == 4'h1 ? {{32'd0}, io_from_lsu_araddr} : _GEN_4878; // @[d_cache.scala 245:27 247:26]
  wire [127:0] _GEN_4916 = state == 4'h1 ? _io_to_lsu_rdata_T_6 : {{64'd0}, _GEN_4893}; // @[d_cache.scala 245:27 262:25]
  wire [39:0] _GEN_1363 = reset ? 40'h0 : _GEN_4761; // @[d_cache.scala 42:{34,34}]
  assign io_to_lsu_rdata = _GEN_4916[63:0];
  assign io_to_lsu_rvalid = state == 4'h1 ? _T_9 : _GEN_4895; // @[d_cache.scala 245:27 264:26]
  assign io_to_lsu_bvalid = state == 4'h1 ? 1'h0 : _GEN_4899; // @[d_cache.scala 245:27 268:26]
  assign io_to_axi_araddr = _GEN_4901[31:0];
  assign io_to_axi_arlen = state == 4'h1 ? 8'h0 : _GEN_4879; // @[d_cache.scala 245:27 248:25]
  assign io_to_axi_arvalid = state == 4'h1 ? 1'h0 : _GEN_4877; // @[d_cache.scala 245:27 246:27]
  assign io_to_axi_rready = state == 4'h1 ? 1'h0 : _GEN_4882; // @[d_cache.scala 245:27 251:26]
  assign io_to_axi_awaddr = state == 4'h1 ? 32'h0 : _GEN_4883; // @[d_cache.scala 245:27 252:26]
  assign io_to_axi_awlen = state == 4'h1 ? 8'h0 : _GEN_4885; // @[d_cache.scala 245:27 254:25]
  assign io_to_axi_awvalid = state == 4'h1 ? 1'h0 : _GEN_4884; // @[d_cache.scala 245:27 253:27]
  assign io_to_axi_wdata = state == 4'h1 ? 64'h0 : _GEN_4888; // @[d_cache.scala 245:27 257:25]
  assign io_to_axi_wstrb = state == 4'h1 ? 8'h0 : _GEN_4889; // @[d_cache.scala 245:27 258:25]
  assign io_to_axi_wvalid = state == 4'h1 ? 1'h0 : _GEN_4891; // @[d_cache.scala 245:27 260:26]
  assign io_to_axi_bready = state == 4'h1 ? 1'h0 : _GEN_4892; // @[d_cache.scala 245:27 261:26]
  always @(posedge clock) begin
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_0 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_0 <= _GEN_523;
        end else begin
          ram_0_0 <= _GEN_3654;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_1 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_1 <= _GEN_524;
        end else begin
          ram_0_1 <= _GEN_3655;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_2 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_2 <= _GEN_525;
        end else begin
          ram_0_2 <= _GEN_3656;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_3 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_3 <= _GEN_526;
        end else begin
          ram_0_3 <= _GEN_3657;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_4 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_4 <= _GEN_527;
        end else begin
          ram_0_4 <= _GEN_3658;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_5 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_5 <= _GEN_528;
        end else begin
          ram_0_5 <= _GEN_3659;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_6 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_6 <= _GEN_529;
        end else begin
          ram_0_6 <= _GEN_3660;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_7 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_7 <= _GEN_530;
        end else begin
          ram_0_7 <= _GEN_3661;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_8 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_8 <= _GEN_531;
        end else begin
          ram_0_8 <= _GEN_3662;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_9 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_9 <= _GEN_532;
        end else begin
          ram_0_9 <= _GEN_3663;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_10 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_10 <= _GEN_533;
        end else begin
          ram_0_10 <= _GEN_3664;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_11 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_11 <= _GEN_534;
        end else begin
          ram_0_11 <= _GEN_3665;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_12 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_12 <= _GEN_535;
        end else begin
          ram_0_12 <= _GEN_3666;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_13 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_13 <= _GEN_536;
        end else begin
          ram_0_13 <= _GEN_3667;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_14 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_14 <= _GEN_537;
        end else begin
          ram_0_14 <= _GEN_3668;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_15 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_0_15 <= _GEN_538;
        end else begin
          ram_0_15 <= _GEN_3669;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_0 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_0 <= _GEN_555;
        end else begin
          ram_1_0 <= _GEN_3718;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_1 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_1 <= _GEN_556;
        end else begin
          ram_1_1 <= _GEN_3719;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_2 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_2 <= _GEN_557;
        end else begin
          ram_1_2 <= _GEN_3720;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_3 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_3 <= _GEN_558;
        end else begin
          ram_1_3 <= _GEN_3721;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_4 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_4 <= _GEN_559;
        end else begin
          ram_1_4 <= _GEN_3722;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_5 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_5 <= _GEN_560;
        end else begin
          ram_1_5 <= _GEN_3723;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_6 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_6 <= _GEN_561;
        end else begin
          ram_1_6 <= _GEN_3724;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_7 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_7 <= _GEN_562;
        end else begin
          ram_1_7 <= _GEN_3725;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_8 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_8 <= _GEN_563;
        end else begin
          ram_1_8 <= _GEN_3726;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_9 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_9 <= _GEN_564;
        end else begin
          ram_1_9 <= _GEN_3727;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_10 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_10 <= _GEN_565;
        end else begin
          ram_1_10 <= _GEN_3728;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_11 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_11 <= _GEN_566;
        end else begin
          ram_1_11 <= _GEN_3729;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_12 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_12 <= _GEN_567;
        end else begin
          ram_1_12 <= _GEN_3730;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_13 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_13 <= _GEN_568;
        end else begin
          ram_1_13 <= _GEN_3731;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_14 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_14 <= _GEN_569;
        end else begin
          ram_1_14 <= _GEN_3732;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_15 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_1_15 <= _GEN_570;
        end else begin
          ram_1_15 <= _GEN_3733;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_0 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_0 <= _GEN_587;
        end else begin
          ram_2_0 <= _GEN_3766;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_1 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_1 <= _GEN_588;
        end else begin
          ram_2_1 <= _GEN_3767;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_2 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_2 <= _GEN_589;
        end else begin
          ram_2_2 <= _GEN_3768;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_3 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_3 <= _GEN_590;
        end else begin
          ram_2_3 <= _GEN_3769;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_4 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_4 <= _GEN_591;
        end else begin
          ram_2_4 <= _GEN_3770;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_5 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_5 <= _GEN_592;
        end else begin
          ram_2_5 <= _GEN_3771;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_6 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_6 <= _GEN_593;
        end else begin
          ram_2_6 <= _GEN_3772;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_7 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_7 <= _GEN_594;
        end else begin
          ram_2_7 <= _GEN_3773;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_8 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_8 <= _GEN_595;
        end else begin
          ram_2_8 <= _GEN_3774;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_9 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_9 <= _GEN_596;
        end else begin
          ram_2_9 <= _GEN_3775;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_10 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_10 <= _GEN_597;
        end else begin
          ram_2_10 <= _GEN_3776;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_11 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_11 <= _GEN_598;
        end else begin
          ram_2_11 <= _GEN_3777;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_12 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_12 <= _GEN_599;
        end else begin
          ram_2_12 <= _GEN_3778;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_13 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_13 <= _GEN_600;
        end else begin
          ram_2_13 <= _GEN_3779;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_14 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_14 <= _GEN_601;
        end else begin
          ram_2_14 <= _GEN_3780;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_15 <= 128'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_2_15 <= _GEN_602;
        end else begin
          ram_2_15 <= _GEN_3781;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_0 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_0 <= _GEN_619;
        end else begin
          ram_3_0 <= _GEN_3814;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_1 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_1 <= _GEN_620;
        end else begin
          ram_3_1 <= _GEN_3815;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_2 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_2 <= _GEN_621;
        end else begin
          ram_3_2 <= _GEN_3816;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_3 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_3 <= _GEN_622;
        end else begin
          ram_3_3 <= _GEN_3817;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_4 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_4 <= _GEN_623;
        end else begin
          ram_3_4 <= _GEN_3818;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_5 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_5 <= _GEN_624;
        end else begin
          ram_3_5 <= _GEN_3819;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_6 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_6 <= _GEN_625;
        end else begin
          ram_3_6 <= _GEN_3820;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_7 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_7 <= _GEN_626;
        end else begin
          ram_3_7 <= _GEN_3821;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_8 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_8 <= _GEN_627;
        end else begin
          ram_3_8 <= _GEN_3822;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_9 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_9 <= _GEN_628;
        end else begin
          ram_3_9 <= _GEN_3823;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_10 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_10 <= _GEN_629;
        end else begin
          ram_3_10 <= _GEN_3824;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_11 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_11 <= _GEN_630;
        end else begin
          ram_3_11 <= _GEN_3825;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_12 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_12 <= _GEN_631;
        end else begin
          ram_3_12 <= _GEN_3826;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_13 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_13 <= _GEN_632;
        end else begin
          ram_3_13 <= _GEN_3827;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_14 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_14 <= _GEN_633;
        end else begin
          ram_3_14 <= _GEN_3828;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_15 <= 128'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          ram_3_15 <= _GEN_634;
        end else begin
          ram_3_15 <= _GEN_3829;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_0 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_0 <= _GEN_3670;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_1 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_1 <= _GEN_3671;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_2 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_2 <= _GEN_3672;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_3 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_3 <= _GEN_3673;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_4 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_4 <= _GEN_3674;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_5 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_5 <= _GEN_3675;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_6 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_6 <= _GEN_3676;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_7 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_7 <= _GEN_3677;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_8 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_8 <= _GEN_3678;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_9 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_9 <= _GEN_3679;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_10 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_10 <= _GEN_3680;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_11 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_11 <= _GEN_3681;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_12 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_12 <= _GEN_3682;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_13 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_13 <= _GEN_3683;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_14 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_14 <= _GEN_3684;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_15 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_0_15 <= _GEN_3685;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_0 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_0 <= _GEN_3734;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_1 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_1 <= _GEN_3735;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_2 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_2 <= _GEN_3736;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_3 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_3 <= _GEN_3737;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_4 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_4 <= _GEN_3738;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_5 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_5 <= _GEN_3739;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_6 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_6 <= _GEN_3740;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_7 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_7 <= _GEN_3741;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_8 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_8 <= _GEN_3742;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_9 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_9 <= _GEN_3743;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_10 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_10 <= _GEN_3744;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_11 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_11 <= _GEN_3745;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_12 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_12 <= _GEN_3746;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_13 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_13 <= _GEN_3747;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_14 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_14 <= _GEN_3748;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_15 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_1_15 <= _GEN_3749;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_0 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_0 <= _GEN_3782;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_1 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_1 <= _GEN_3783;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_2 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_2 <= _GEN_3784;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_3 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_3 <= _GEN_3785;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_4 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_4 <= _GEN_3786;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_5 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_5 <= _GEN_3787;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_6 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_6 <= _GEN_3788;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_7 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_7 <= _GEN_3789;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_8 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_8 <= _GEN_3790;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_9 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_9 <= _GEN_3791;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_10 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_10 <= _GEN_3792;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_11 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_11 <= _GEN_3793;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_12 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_12 <= _GEN_3794;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_13 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_13 <= _GEN_3795;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_14 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_14 <= _GEN_3796;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_15 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_2_15 <= _GEN_3797;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_0 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_0 <= _GEN_3830;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_1 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_1 <= _GEN_3831;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_2 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_2 <= _GEN_3832;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_3 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_3 <= _GEN_3833;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_4 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_4 <= _GEN_3834;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_5 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_5 <= _GEN_3835;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_6 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_6 <= _GEN_3836;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_7 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_7 <= _GEN_3837;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_8 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_8 <= _GEN_3838;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_9 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_9 <= _GEN_3839;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_10 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_10 <= _GEN_3840;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_11 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_11 <= _GEN_3841;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_12 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_12 <= _GEN_3842;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_13 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_13 <= _GEN_3843;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_14 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_14 <= _GEN_3844;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_15 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          tag_3_15 <= _GEN_3845;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_0 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_0 <= _GEN_3686;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_1 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_1 <= _GEN_3687;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_2 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_2 <= _GEN_3688;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_3 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_3 <= _GEN_3689;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_4 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_4 <= _GEN_3690;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_5 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_5 <= _GEN_3691;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_6 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_6 <= _GEN_3692;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_7 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_7 <= _GEN_3693;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_8 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_8 <= _GEN_3694;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_9 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_9 <= _GEN_3695;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_10 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_10 <= _GEN_3696;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_11 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_11 <= _GEN_3697;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_12 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_12 <= _GEN_3698;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_13 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_13 <= _GEN_3699;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_14 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_14 <= _GEN_3700;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:26]
      valid_0_15 <= 1'h0; // @[d_cache.scala 28:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_0_15 <= _GEN_3701;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_0 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_0 <= _GEN_3750;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_1 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_1 <= _GEN_3751;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_2 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_2 <= _GEN_3752;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_3 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_3 <= _GEN_3753;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_4 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_4 <= _GEN_3754;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_5 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_5 <= _GEN_3755;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_6 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_6 <= _GEN_3756;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_7 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_7 <= _GEN_3757;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_8 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_8 <= _GEN_3758;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_9 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_9 <= _GEN_3759;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_10 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_10 <= _GEN_3760;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_11 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_11 <= _GEN_3761;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_12 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_12 <= _GEN_3762;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_13 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_13 <= _GEN_3763;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_14 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_14 <= _GEN_3764;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_1_15 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_1_15 <= _GEN_3765;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_0 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_0 <= _GEN_3798;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_1 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_1 <= _GEN_3799;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_2 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_2 <= _GEN_3800;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_3 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_3 <= _GEN_3801;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_4 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_4 <= _GEN_3802;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_5 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_5 <= _GEN_3803;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_6 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_6 <= _GEN_3804;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_7 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_7 <= _GEN_3805;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_8 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_8 <= _GEN_3806;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_9 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_9 <= _GEN_3807;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_10 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_10 <= _GEN_3808;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_11 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_11 <= _GEN_3809;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_12 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_12 <= _GEN_3810;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_13 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_13 <= _GEN_3811;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_14 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_14 <= _GEN_3812;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_2_15 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_2_15 <= _GEN_3813;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_0 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_0 <= _GEN_3846;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_1 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_1 <= _GEN_3847;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_2 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_2 <= _GEN_3848;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_3 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_3 <= _GEN_3849;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_4 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_4 <= _GEN_3850;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_5 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_5 <= _GEN_3851;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_6 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_6 <= _GEN_3852;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_7 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_7 <= _GEN_3853;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_8 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_8 <= _GEN_3854;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_9 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_9 <= _GEN_3855;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_10 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_10 <= _GEN_3856;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_11 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_11 <= _GEN_3857;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_12 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_12 <= _GEN_3858;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_13 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_13 <= _GEN_3859;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_14 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_14 <= _GEN_3860;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_3_15 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          valid_3_15 <= _GEN_3861;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_0 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_0 <= _GEN_539;
        end else begin
          dirty_0_0 <= _GEN_3864;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_1 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_1 <= _GEN_540;
        end else begin
          dirty_0_1 <= _GEN_3865;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_2 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_2 <= _GEN_541;
        end else begin
          dirty_0_2 <= _GEN_3866;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_3 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_3 <= _GEN_542;
        end else begin
          dirty_0_3 <= _GEN_3867;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_4 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_4 <= _GEN_543;
        end else begin
          dirty_0_4 <= _GEN_3868;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_5 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_5 <= _GEN_544;
        end else begin
          dirty_0_5 <= _GEN_3869;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_6 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_6 <= _GEN_545;
        end else begin
          dirty_0_6 <= _GEN_3870;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_7 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_7 <= _GEN_546;
        end else begin
          dirty_0_7 <= _GEN_3871;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_8 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_8 <= _GEN_547;
        end else begin
          dirty_0_8 <= _GEN_3872;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_9 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_9 <= _GEN_548;
        end else begin
          dirty_0_9 <= _GEN_3873;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_10 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_10 <= _GEN_549;
        end else begin
          dirty_0_10 <= _GEN_3874;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_11 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_11 <= _GEN_550;
        end else begin
          dirty_0_11 <= _GEN_3875;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_12 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_12 <= _GEN_551;
        end else begin
          dirty_0_12 <= _GEN_3876;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_13 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_13 <= _GEN_552;
        end else begin
          dirty_0_13 <= _GEN_3877;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_14 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_14 <= _GEN_553;
        end else begin
          dirty_0_14 <= _GEN_3878;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_15 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_0_15 <= _GEN_554;
        end else begin
          dirty_0_15 <= _GEN_3879;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_0 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_0 <= _GEN_635;
        end else begin
          dirty_3_0 <= _GEN_3912;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_1 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_1 <= _GEN_636;
        end else begin
          dirty_3_1 <= _GEN_3913;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_2 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_2 <= _GEN_637;
        end else begin
          dirty_3_2 <= _GEN_3914;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_3 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_3 <= _GEN_638;
        end else begin
          dirty_3_3 <= _GEN_3915;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_4 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_4 <= _GEN_639;
        end else begin
          dirty_3_4 <= _GEN_3916;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_5 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_5 <= _GEN_640;
        end else begin
          dirty_3_5 <= _GEN_3917;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_6 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_6 <= _GEN_641;
        end else begin
          dirty_3_6 <= _GEN_3918;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_7 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_7 <= _GEN_642;
        end else begin
          dirty_3_7 <= _GEN_3919;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_8 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_8 <= _GEN_643;
        end else begin
          dirty_3_8 <= _GEN_3920;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_9 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_9 <= _GEN_644;
        end else begin
          dirty_3_9 <= _GEN_3921;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_10 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_10 <= _GEN_645;
        end else begin
          dirty_3_10 <= _GEN_3922;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_11 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_11 <= _GEN_646;
        end else begin
          dirty_3_11 <= _GEN_3923;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_12 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_12 <= _GEN_647;
        end else begin
          dirty_3_12 <= _GEN_3924;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_13 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_13 <= _GEN_648;
        end else begin
          dirty_3_13 <= _GEN_3925;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_14 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_14 <= _GEN_649;
        end else begin
          dirty_3_14 <= _GEN_3926;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_3_15 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (4'h2 == state) begin // @[d_cache.scala 76:18]
          dirty_3_15 <= _GEN_650;
        end else begin
          dirty_3_15 <= _GEN_3927;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 41:34]
      write_back_data <= 128'h0; // @[d_cache.scala 41:34]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          write_back_data <= _GEN_3862;
        end
      end
    end
    write_back_addr <= _GEN_1363[31:0]; // @[d_cache.scala 42:{34,34}]
    if (reset) begin // @[d_cache.scala 47:31]
      receive_data_0 <= 64'h0; // @[d_cache.scala 47:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          receive_data_0 <= _GEN_3650;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 47:31]
      receive_data_1 <= 64'h0; // @[d_cache.scala 47:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          receive_data_1 <= _GEN_3651;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 48:30]
      receive_num <= 3'h0; // @[d_cache.scala 48:30]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (4'h1 == state) begin // @[d_cache.scala 76:18]
        if (!(way0_hit | way1_hit | way2_hit | way3_hit)) begin // @[d_cache.scala 87:57]
          receive_num <= 3'h0; // @[d_cache.scala 93:29]
        end
      end else if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
        receive_num <= _GEN_3652;
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_0 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_0 <= _GEN_3702;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_1 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_1 <= _GEN_3703;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_2 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_2 <= _GEN_3704;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_3 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_3 <= _GEN_3705;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_4 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_4 <= _GEN_3706;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_5 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_5 <= _GEN_3707;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_6 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_6 <= _GEN_3708;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_7 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_7 <= _GEN_3709;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_8 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_8 <= _GEN_3710;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_9 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_9 <= _GEN_3711;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_10 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_10 <= _GEN_3712;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_11 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_11 <= _GEN_3713;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_12 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_12 <= _GEN_3714;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_13 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_13 <= _GEN_3715;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_14 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_14 <= _GEN_3716;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 49:24]
      quene_15 <= 8'h0; // @[d_cache.scala 49:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 76:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 76:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 76:18]
          quene_15 <= _GEN_3717;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 71:24]
      state <= 4'h0; // @[d_cache.scala 71:24]
    end else if (4'h0 == state) begin // @[d_cache.scala 76:18]
      if ((io_from_lsu_arvalid | io_from_lsu_awvalid) & io_from_lsu_araddr >= 32'ha0000000) begin // @[d_cache.scala 78:99]
        state <= 4'h0; // @[d_cache.scala 79:23]
      end else if (io_from_lsu_arvalid) begin // @[d_cache.scala 80:44]
        state <= 4'h1; // @[d_cache.scala 81:23]
      end else begin
        state <= _GEN_128;
      end
    end else if (4'h1 == state) begin // @[d_cache.scala 76:18]
      if (way0_hit | way1_hit | way2_hit | way3_hit) begin // @[d_cache.scala 87:57]
        state <= 4'h0;
      end else begin
        state <= 4'h3; // @[d_cache.scala 92:23]
      end
    end else if (4'h2 == state) begin // @[d_cache.scala 76:18]
      state <= _GEN_522;
    end else begin
      state <= _GEN_3653;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"d_cache state:%d\n",state); // @[d_cache.scala 72:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  ram_0_0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  ram_0_1 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  ram_0_2 = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  ram_0_3 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  ram_0_4 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  ram_0_5 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  ram_0_6 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  ram_0_7 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  ram_0_8 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  ram_0_9 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  ram_0_10 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  ram_0_11 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  ram_0_12 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  ram_0_13 = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  ram_0_14 = _RAND_14[127:0];
  _RAND_15 = {4{`RANDOM}};
  ram_0_15 = _RAND_15[127:0];
  _RAND_16 = {4{`RANDOM}};
  ram_1_0 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  ram_1_1 = _RAND_17[127:0];
  _RAND_18 = {4{`RANDOM}};
  ram_1_2 = _RAND_18[127:0];
  _RAND_19 = {4{`RANDOM}};
  ram_1_3 = _RAND_19[127:0];
  _RAND_20 = {4{`RANDOM}};
  ram_1_4 = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  ram_1_5 = _RAND_21[127:0];
  _RAND_22 = {4{`RANDOM}};
  ram_1_6 = _RAND_22[127:0];
  _RAND_23 = {4{`RANDOM}};
  ram_1_7 = _RAND_23[127:0];
  _RAND_24 = {4{`RANDOM}};
  ram_1_8 = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  ram_1_9 = _RAND_25[127:0];
  _RAND_26 = {4{`RANDOM}};
  ram_1_10 = _RAND_26[127:0];
  _RAND_27 = {4{`RANDOM}};
  ram_1_11 = _RAND_27[127:0];
  _RAND_28 = {4{`RANDOM}};
  ram_1_12 = _RAND_28[127:0];
  _RAND_29 = {4{`RANDOM}};
  ram_1_13 = _RAND_29[127:0];
  _RAND_30 = {4{`RANDOM}};
  ram_1_14 = _RAND_30[127:0];
  _RAND_31 = {4{`RANDOM}};
  ram_1_15 = _RAND_31[127:0];
  _RAND_32 = {4{`RANDOM}};
  ram_2_0 = _RAND_32[127:0];
  _RAND_33 = {4{`RANDOM}};
  ram_2_1 = _RAND_33[127:0];
  _RAND_34 = {4{`RANDOM}};
  ram_2_2 = _RAND_34[127:0];
  _RAND_35 = {4{`RANDOM}};
  ram_2_3 = _RAND_35[127:0];
  _RAND_36 = {4{`RANDOM}};
  ram_2_4 = _RAND_36[127:0];
  _RAND_37 = {4{`RANDOM}};
  ram_2_5 = _RAND_37[127:0];
  _RAND_38 = {4{`RANDOM}};
  ram_2_6 = _RAND_38[127:0];
  _RAND_39 = {4{`RANDOM}};
  ram_2_7 = _RAND_39[127:0];
  _RAND_40 = {4{`RANDOM}};
  ram_2_8 = _RAND_40[127:0];
  _RAND_41 = {4{`RANDOM}};
  ram_2_9 = _RAND_41[127:0];
  _RAND_42 = {4{`RANDOM}};
  ram_2_10 = _RAND_42[127:0];
  _RAND_43 = {4{`RANDOM}};
  ram_2_11 = _RAND_43[127:0];
  _RAND_44 = {4{`RANDOM}};
  ram_2_12 = _RAND_44[127:0];
  _RAND_45 = {4{`RANDOM}};
  ram_2_13 = _RAND_45[127:0];
  _RAND_46 = {4{`RANDOM}};
  ram_2_14 = _RAND_46[127:0];
  _RAND_47 = {4{`RANDOM}};
  ram_2_15 = _RAND_47[127:0];
  _RAND_48 = {4{`RANDOM}};
  ram_3_0 = _RAND_48[127:0];
  _RAND_49 = {4{`RANDOM}};
  ram_3_1 = _RAND_49[127:0];
  _RAND_50 = {4{`RANDOM}};
  ram_3_2 = _RAND_50[127:0];
  _RAND_51 = {4{`RANDOM}};
  ram_3_3 = _RAND_51[127:0];
  _RAND_52 = {4{`RANDOM}};
  ram_3_4 = _RAND_52[127:0];
  _RAND_53 = {4{`RANDOM}};
  ram_3_5 = _RAND_53[127:0];
  _RAND_54 = {4{`RANDOM}};
  ram_3_6 = _RAND_54[127:0];
  _RAND_55 = {4{`RANDOM}};
  ram_3_7 = _RAND_55[127:0];
  _RAND_56 = {4{`RANDOM}};
  ram_3_8 = _RAND_56[127:0];
  _RAND_57 = {4{`RANDOM}};
  ram_3_9 = _RAND_57[127:0];
  _RAND_58 = {4{`RANDOM}};
  ram_3_10 = _RAND_58[127:0];
  _RAND_59 = {4{`RANDOM}};
  ram_3_11 = _RAND_59[127:0];
  _RAND_60 = {4{`RANDOM}};
  ram_3_12 = _RAND_60[127:0];
  _RAND_61 = {4{`RANDOM}};
  ram_3_13 = _RAND_61[127:0];
  _RAND_62 = {4{`RANDOM}};
  ram_3_14 = _RAND_62[127:0];
  _RAND_63 = {4{`RANDOM}};
  ram_3_15 = _RAND_63[127:0];
  _RAND_64 = {1{`RANDOM}};
  tag_0_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  tag_0_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  tag_0_2 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  tag_0_3 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  tag_0_4 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  tag_0_5 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  tag_0_6 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  tag_0_7 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  tag_0_8 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  tag_0_9 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  tag_0_10 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  tag_0_11 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  tag_0_12 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  tag_0_13 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  tag_0_14 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  tag_0_15 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  tag_1_0 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  tag_1_1 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  tag_1_2 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  tag_1_3 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  tag_1_4 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  tag_1_5 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  tag_1_6 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  tag_1_7 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  tag_1_8 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  tag_1_9 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  tag_1_10 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  tag_1_11 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  tag_1_12 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  tag_1_13 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  tag_1_14 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  tag_1_15 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  tag_2_0 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  tag_2_1 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  tag_2_2 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  tag_2_3 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  tag_2_4 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  tag_2_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  tag_2_6 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  tag_2_7 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  tag_2_8 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  tag_2_9 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  tag_2_10 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  tag_2_11 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  tag_2_12 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  tag_2_13 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  tag_2_14 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  tag_2_15 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  tag_3_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  tag_3_1 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  tag_3_2 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  tag_3_3 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  tag_3_4 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  tag_3_5 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  tag_3_6 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  tag_3_7 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  tag_3_8 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  tag_3_9 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  tag_3_10 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  tag_3_11 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  tag_3_12 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  tag_3_13 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  tag_3_14 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  tag_3_15 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  valid_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_0_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_0_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_0_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_0_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_0_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_0_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_0_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_0_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_0_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_0_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_0_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_0_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_0_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_0_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_1_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_1_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_1_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_1_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_1_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_1_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_1_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_1_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_1_8 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_1_9 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_1_10 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_1_11 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_1_12 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_1_13 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_1_14 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_1_15 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_2_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_2_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_2_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_2_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_2_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_2_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_2_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_2_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_2_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_2_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_2_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_2_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_2_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_2_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_2_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_2_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_3_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_3_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_3_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_3_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_3_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_3_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_3_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_3_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_3_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_3_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_3_10 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_3_11 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_3_12 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_3_13 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_3_14 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_3_15 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  dirty_0_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  dirty_0_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  dirty_0_2 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  dirty_0_3 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  dirty_0_4 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  dirty_0_5 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  dirty_0_6 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  dirty_0_7 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  dirty_0_8 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  dirty_0_9 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  dirty_0_10 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  dirty_0_11 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  dirty_0_12 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  dirty_0_13 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  dirty_0_14 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  dirty_0_15 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  dirty_3_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  dirty_3_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  dirty_3_2 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  dirty_3_3 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  dirty_3_4 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  dirty_3_5 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  dirty_3_6 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  dirty_3_7 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  dirty_3_8 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  dirty_3_9 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  dirty_3_10 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  dirty_3_11 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  dirty_3_12 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  dirty_3_13 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  dirty_3_14 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  dirty_3_15 = _RAND_223[0:0];
  _RAND_224 = {4{`RANDOM}};
  write_back_data = _RAND_224[127:0];
  _RAND_225 = {1{`RANDOM}};
  write_back_addr = _RAND_225[31:0];
  _RAND_226 = {2{`RANDOM}};
  receive_data_0 = _RAND_226[63:0];
  _RAND_227 = {2{`RANDOM}};
  receive_data_1 = _RAND_227[63:0];
  _RAND_228 = {1{`RANDOM}};
  receive_num = _RAND_228[2:0];
  _RAND_229 = {1{`RANDOM}};
  quene_0 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  quene_1 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  quene_2 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  quene_3 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  quene_4 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  quene_5 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  quene_6 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  quene_7 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  quene_8 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  quene_9 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  quene_10 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  quene_11 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  quene_12 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  quene_13 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  quene_14 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  quene_15 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  state = _RAND_245[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
