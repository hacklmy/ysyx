module AXI(
  input         clock,
  input         reset,
  input  [31:0] io_axi_in_araddr,
  input         io_axi_in_arvalid,
  input         io_axi_in_rready,
  input  [31:0] io_axi_in_awaddr,
  input         io_axi_in_awvalid,
  input  [63:0] io_axi_in_wdata,
  input  [7:0]  io_axi_in_wstrb,
  input         io_axi_in_wvalid,
  input         io_axi_in_bready,
  output        io_axi_out_arready,
  output [63:0] io_axi_out_rdata,
  output        io_axi_out_rvalid,
  output        io_axi_out_awready,
  output        io_axi_out_wready,
  output        io_axi_out_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] Mem_modle_Raddr; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Rdata; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Waddr; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Wdata; // @[AXI.scala 26:27]
  wire [7:0] Mem_modle_Wmask; // @[AXI.scala 26:27]
  wire  Mem_modle_Write_en; // @[AXI.scala 26:27]
  wire  Mem_modle_Read_en; // @[AXI.scala 26:27]
  reg  axi_awready; // @[AXI.scala 13:30]
  reg  axi_wready; // @[AXI.scala 14:29]
  reg  axi_bvalid; // @[AXI.scala 17:29]
  reg  axi_arready; // @[AXI.scala 19:30]
  reg  axi_rvalid; // @[AXI.scala 21:29]
  reg [2:0] state; // @[AXI.scala 24:24]
  wire  _GEN_1 = io_axi_in_arvalid ? 1'h0 : axi_arready; // @[AXI.scala 49:42 51:29 19:30]
  wire  _GEN_2 = io_axi_in_arvalid | axi_rvalid; // @[AXI.scala 49:42 52:28 21:29]
  wire  _GEN_4 = io_axi_in_awvalid & io_axi_in_wvalid ? 1'h0 : axi_awready; // @[AXI.scala 39:56 41:29 13:30]
  wire  _GEN_5 = io_axi_in_awvalid & io_axi_in_wvalid ? 1'h0 : axi_wready; // @[AXI.scala 39:56 42:28 14:29]
  wire  _GEN_6 = io_axi_in_awvalid & io_axi_in_wvalid | axi_bvalid; // @[AXI.scala 39:56 43:28 17:29]
  wire  _GEN_7 = io_axi_in_awvalid & io_axi_in_wvalid ? axi_arready : _GEN_1; // @[AXI.scala 19:30 39:56]
  wire  _GEN_11 = io_axi_in_bready | axi_awready; // @[AXI.scala 56:35 59:29 13:30]
  wire  _GEN_12 = io_axi_in_bready | axi_wready; // @[AXI.scala 56:35 60:28 14:29]
  wire [2:0] _GEN_13 = io_axi_in_rready ? 3'h0 : state; // @[AXI.scala 64:35 65:23 24:24]
  wire  _GEN_14 = io_axi_in_rready | axi_arready; // @[AXI.scala 64:35 66:29 19:30]
  wire  _GEN_15 = io_axi_in_rready ? 1'h0 : axi_rvalid; // @[AXI.scala 64:35 67:28 21:29]
  wire  _GEN_17 = 3'h4 == state ? _GEN_14 : axi_arready; // @[AXI.scala 37:18 19:30]
  wire  _GEN_21 = 3'h3 == state ? _GEN_11 : axi_awready; // @[AXI.scala 37:18 13:30]
  wire  _GEN_22 = 3'h3 == state ? _GEN_12 : axi_wready; // @[AXI.scala 37:18 14:29]
  wire  _GEN_23 = 3'h3 == state ? axi_arready : _GEN_17; // @[AXI.scala 37:18 19:30]
  wire  _GEN_26 = 3'h0 == state ? _GEN_4 : _GEN_21; // @[AXI.scala 37:18]
  wire  _GEN_27 = 3'h0 == state ? _GEN_5 : _GEN_22; // @[AXI.scala 37:18]
  wire  _GEN_29 = 3'h0 == state ? _GEN_7 : _GEN_23; // @[AXI.scala 37:18]
  MEM Mem_modle ( // @[AXI.scala 26:27]
    .Raddr(Mem_modle_Raddr),
    .Rdata(Mem_modle_Rdata),
    .Waddr(Mem_modle_Waddr),
    .Wdata(Mem_modle_Wdata),
    .Wmask(Mem_modle_Wmask),
    .Write_en(Mem_modle_Write_en),
    .Read_en(Mem_modle_Read_en)
  );
  assign io_axi_out_arready = axi_arready; // @[AXI.scala 71:24]
  assign io_axi_out_rdata = Mem_modle_Rdata; // @[AXI.scala 72:22]
  assign io_axi_out_rvalid = axi_rvalid; // @[AXI.scala 73:23]
  assign io_axi_out_awready = axi_awready; // @[AXI.scala 74:24]
  assign io_axi_out_wready = axi_wready; // @[AXI.scala 75:23]
  assign io_axi_out_bvalid = axi_bvalid; // @[AXI.scala 76:23]
  assign Mem_modle_Raddr = {32'h0,io_axi_in_araddr}; // @[Cat.scala 31:58]
  assign Mem_modle_Waddr = {{32'd0}, io_axi_in_awaddr}; // @[AXI.scala 28:24]
  assign Mem_modle_Wdata = io_axi_in_wdata; // @[AXI.scala 29:24]
  assign Mem_modle_Wmask = io_axi_in_wstrb; // @[AXI.scala 30:24]
  assign Mem_modle_Write_en = axi_wready & io_axi_in_wvalid; // @[AXI.scala 31:48]
  assign Mem_modle_Read_en = axi_arready & io_axi_in_arvalid; // @[AXI.scala 32:48]
  always @(posedge clock) begin
    axi_awready <= reset | _GEN_26; // @[AXI.scala 13:{30,30}]
    axi_wready <= reset | _GEN_27; // @[AXI.scala 14:{29,29}]
    if (reset) begin // @[AXI.scala 17:29]
      axi_bvalid <= 1'h0; // @[AXI.scala 17:29]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      axi_bvalid <= _GEN_6;
    end else if (3'h3 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_bready) begin // @[AXI.scala 56:35]
        axi_bvalid <= 1'h0; // @[AXI.scala 58:28]
      end
    end
    axi_arready <= reset | _GEN_29; // @[AXI.scala 19:{30,30}]
    if (reset) begin // @[AXI.scala 21:29]
      axi_rvalid <= 1'h0; // @[AXI.scala 21:29]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      if (!(io_axi_in_awvalid & io_axi_in_wvalid)) begin // @[AXI.scala 39:56]
        axi_rvalid <= _GEN_2;
      end
    end else if (!(3'h3 == state)) begin // @[AXI.scala 37:18]
      if (3'h4 == state) begin // @[AXI.scala 37:18]
        axi_rvalid <= _GEN_15;
      end
    end
    if (reset) begin // @[AXI.scala 24:24]
      state <= 3'h0; // @[AXI.scala 24:24]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_awvalid & io_axi_in_wvalid) begin // @[AXI.scala 39:56]
        state <= 3'h3; // @[AXI.scala 40:23]
      end else if (io_axi_in_arvalid) begin // @[AXI.scala 49:42]
        state <= 3'h4; // @[AXI.scala 50:23]
      end
    end else if (3'h3 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_bready) begin // @[AXI.scala 56:35]
        state <= 3'h0; // @[AXI.scala 57:23]
      end
    end else if (3'h4 == state) begin // @[AXI.scala 37:18]
      state <= _GEN_13;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_awready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  axi_wready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  axi_bvalid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  axi_arready = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  axi_rvalid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSU(
  input         clock,
  input         reset,
  input         io_inst_store,
  input         io_inst_load,
  input  [31:0] io_mem_addr,
  input  [63:0] io_mem_wdata,
  input  [7:0]  io_mem_wstrb,
  output [63:0] io_mem_rdata,
  input         io_axi_in_arready,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  input         io_axi_in_awready,
  input         io_axi_in_wready,
  input         io_axi_in_bvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  output [31:0] io_axi_out_awaddr,
  output        io_axi_out_awvalid,
  output [63:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid,
  output        io_axi_out_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  axi_arvalid; // @[LSU.scala 19:30]
  reg  axi_rready; // @[LSU.scala 22:29]
  reg  axi_awvalid; // @[LSU.scala 23:30]
  reg  axi_wvalid; // @[LSU.scala 24:29]
  reg  axi_bready; // @[LSU.scala 25:29]
  reg [1:0] state; // @[LSU.scala 28:24]
  wire  _GEN_1 = io_inst_store | axi_awvalid; // @[LSU.scala 36:38 38:29 23:30]
  wire  _GEN_2 = io_inst_store | axi_wvalid; // @[LSU.scala 36:38 39:28 24:29]
  wire  _GEN_3 = io_inst_store | axi_bready; // @[LSU.scala 36:38 40:28 25:29]
  wire  _GEN_5 = io_inst_load | axi_arvalid; // @[LSU.scala 32:31 34:29 19:30]
  wire  _GEN_6 = io_inst_load | axi_rready; // @[LSU.scala 32:31 35:28 22:29]
  wire  _GEN_9 = io_inst_load ? axi_bready : _GEN_3; // @[LSU.scala 25:29 32:31]
  wire  _GEN_11 = io_axi_in_bvalid ? 1'h0 : axi_bready; // @[LSU.scala 44:35 46:28 25:29]
  wire  _GEN_14 = io_axi_in_arready ? 1'h0 : axi_arvalid; // @[LSU.scala 56:36 57:29 19:30]
  wire [1:0] _GEN_15 = io_axi_in_rvalid ? 2'h0 : state; // @[LSU.scala 59:35 60:23 28:24]
  wire  _GEN_16 = io_axi_in_rvalid ? 1'h0 : axi_rready; // @[LSU.scala 59:35 61:28 22:29]
  wire  _GEN_19 = 2'h2 == state ? _GEN_16 : axi_rready; // @[LSU.scala 30:18 22:29]
  wire  _GEN_21 = 2'h1 == state ? _GEN_11 : axi_bready; // @[LSU.scala 30:18 25:29]
  wire  _GEN_25 = 2'h1 == state ? axi_rready : _GEN_19; // @[LSU.scala 30:18 22:29]
  wire  _GEN_28 = 2'h0 == state ? _GEN_6 : _GEN_25; // @[LSU.scala 30:18]
  wire  _GEN_31 = 2'h0 == state ? _GEN_9 : _GEN_21; // @[LSU.scala 30:18]
  assign io_mem_rdata = io_axi_in_rdata; // @[LSU.scala 72:18]
  assign io_axi_out_araddr = io_mem_addr; // @[LSU.scala 73:23]
  assign io_axi_out_arvalid = axi_arvalid; // @[LSU.scala 74:24]
  assign io_axi_out_rready = axi_rready; // @[LSU.scala 75:23]
  assign io_axi_out_awaddr = io_mem_addr; // @[LSU.scala 76:23]
  assign io_axi_out_awvalid = axi_awvalid; // @[LSU.scala 77:24]
  assign io_axi_out_wdata = io_mem_wdata; // @[LSU.scala 78:22]
  assign io_axi_out_wstrb = io_mem_wstrb; // @[LSU.scala 79:22]
  assign io_axi_out_wvalid = axi_wvalid; // @[LSU.scala 80:23]
  assign io_axi_out_bready = axi_bready; // @[LSU.scala 81:23]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 19:30]
      axi_arvalid <= 1'h0; // @[LSU.scala 19:30]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      axi_arvalid <= _GEN_5;
    end else if (!(2'h1 == state)) begin // @[LSU.scala 30:18]
      if (2'h2 == state) begin // @[LSU.scala 30:18]
        axi_arvalid <= _GEN_14;
      end
    end
    axi_rready <= reset | _GEN_28; // @[LSU.scala 22:{29,29}]
    if (reset) begin // @[LSU.scala 23:30]
      axi_awvalid <= 1'h0; // @[LSU.scala 23:30]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (!(io_inst_load)) begin // @[LSU.scala 32:31]
        axi_awvalid <= _GEN_1;
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_awready) begin // @[LSU.scala 51:36]
        axi_awvalid <= 1'h0; // @[LSU.scala 52:29]
      end
    end
    if (reset) begin // @[LSU.scala 24:29]
      axi_wvalid <= 1'h0; // @[LSU.scala 24:29]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (!(io_inst_load)) begin // @[LSU.scala 32:31]
        axi_wvalid <= _GEN_2;
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_wready) begin // @[LSU.scala 48:35]
        axi_wvalid <= 1'h0; // @[LSU.scala 49:28]
      end
    end
    axi_bready <= reset | _GEN_31; // @[LSU.scala 25:{29,29}]
    if (reset) begin // @[LSU.scala 28:24]
      state <= 2'h0; // @[LSU.scala 28:24]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (io_inst_load) begin // @[LSU.scala 32:31]
        state <= 2'h2; // @[LSU.scala 33:23]
      end else if (io_inst_store) begin // @[LSU.scala 36:38]
        state <= 2'h1; // @[LSU.scala 37:23]
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_bvalid) begin // @[LSU.scala 44:35]
        state <= 2'h0; // @[LSU.scala 45:23]
      end
    end else if (2'h2 == state) begin // @[LSU.scala 30:18]
      state <= _GEN_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_arvalid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  axi_rready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  axi_awvalid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  axi_wvalid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  axi_bready = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI_ARBITER(
  input         clock,
  input         reset,
  input  [31:0] io_ifu_axi_in_araddr,
  input         io_ifu_axi_in_arvalid,
  input         io_ifu_axi_in_rready,
  output [63:0] io_ifu_axi_out_rdata,
  output        io_ifu_axi_out_rvalid,
  input  [31:0] io_lsu_axi_in_araddr,
  input         io_lsu_axi_in_arvalid,
  input         io_lsu_axi_in_rready,
  input  [31:0] io_lsu_axi_in_awaddr,
  input         io_lsu_axi_in_awvalid,
  input  [63:0] io_lsu_axi_in_wdata,
  input  [7:0]  io_lsu_axi_in_wstrb,
  input         io_lsu_axi_in_wvalid,
  input         io_lsu_axi_in_bready,
  output        io_lsu_axi_out_arready,
  output [63:0] io_lsu_axi_out_rdata,
  output        io_lsu_axi_out_rvalid,
  output        io_lsu_axi_out_awready,
  output        io_lsu_axi_out_wready,
  output        io_lsu_axi_out_bvalid,
  input         io_axi_in_arready,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  input         io_axi_in_awready,
  input         io_axi_in_wready,
  input         io_axi_in_bvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  output [31:0] io_axi_out_awaddr,
  output        io_axi_out_awvalid,
  output [63:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid,
  output        io_axi_out_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[axi_arbiter.scala 18:24]
  wire [1:0] _GEN_0 = io_ifu_axi_in_arvalid ? 2'h1 : state; // @[axi_arbiter.scala 51:46 52:23 18:24]
  wire [31:0] _GEN_1 = io_ifu_axi_in_arvalid ? io_ifu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 51:46 53:28 57:28]
  wire  _GEN_3 = io_ifu_axi_in_arvalid & io_ifu_axi_in_rready; // @[axi_arbiter.scala 51:46 53:28 57:28]
  wire [63:0] _GEN_11 = io_ifu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 51:46 54:32 59:32]
  wire  _GEN_12 = io_ifu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 51:46 54:32 59:32]
  wire [31:0] _GEN_23 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_araddr : _GEN_1; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_24 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_arvalid : io_ifu_axi_in_arvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_25 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_rready : _GEN_3; // @[axi_arbiter.scala 46:46 48:28]
  wire [31:0] _GEN_26 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_27 = io_lsu_axi_in_arvalid & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire [63:0] _GEN_28 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wdata : 64'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire [7:0] _GEN_29 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_30 = io_lsu_axi_in_arvalid & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_31 = io_lsu_axi_in_arvalid & io_lsu_axi_in_bready; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_32 = io_lsu_axi_in_arvalid & io_axi_in_arready; // @[axi_arbiter.scala 46:46 49:32]
  wire [63:0] _GEN_33 = io_lsu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_34 = io_lsu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_35 = io_lsu_axi_in_arvalid & io_axi_in_awready; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_36 = io_lsu_axi_in_arvalid & io_axi_in_wready; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_37 = io_lsu_axi_in_arvalid & io_axi_in_bvalid; // @[axi_arbiter.scala 46:46 49:32]
  wire [63:0] _GEN_39 = io_lsu_axi_in_arvalid ? 64'h0 : _GEN_11; // @[axi_arbiter.scala 46:46 50:32]
  wire  _GEN_40 = io_lsu_axi_in_arvalid ? 1'h0 : _GEN_12; // @[axi_arbiter.scala 46:46 50:32]
  wire [31:0] _GEN_45 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_araddr : _GEN_23; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_46 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_arvalid : _GEN_24; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_47 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_rready : _GEN_25; // @[axi_arbiter.scala 41:40 43:28]
  wire [31:0] _GEN_48 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awaddr : _GEN_26; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_49 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awvalid : _GEN_27; // @[axi_arbiter.scala 41:40 43:28]
  wire [63:0] _GEN_50 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wdata : _GEN_28; // @[axi_arbiter.scala 41:40 43:28]
  wire [7:0] _GEN_51 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wstrb : _GEN_29; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_52 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wvalid : _GEN_30; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_53 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_bready : _GEN_31; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_54 = io_lsu_axi_in_awvalid ? io_axi_in_arready : _GEN_32; // @[axi_arbiter.scala 41:40 44:32]
  wire [63:0] _GEN_55 = io_lsu_axi_in_awvalid ? io_axi_in_rdata : _GEN_33; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_56 = io_lsu_axi_in_awvalid ? io_axi_in_rvalid : _GEN_34; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_57 = io_lsu_axi_in_awvalid ? io_axi_in_awready : _GEN_35; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_58 = io_lsu_axi_in_awvalid ? io_axi_in_wready : _GEN_36; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_59 = io_lsu_axi_in_awvalid ? io_axi_in_bvalid : _GEN_37; // @[axi_arbiter.scala 41:40 44:32]
  wire [63:0] _GEN_61 = io_lsu_axi_in_awvalid ? 64'h0 : _GEN_39; // @[axi_arbiter.scala 41:40 45:32]
  wire  _GEN_62 = io_lsu_axi_in_awvalid ? 1'h0 : _GEN_40; // @[axi_arbiter.scala 41:40 45:32]
  wire [1:0] _GEN_67 = io_lsu_axi_out_rvalid & io_lsu_axi_in_rready ? 2'h0 : state; // @[axi_arbiter.scala 74:64 75:23 18:24]
  wire [1:0] _GEN_68 = io_lsu_axi_out_bvalid & io_lsu_axi_in_bready ? 2'h0 : state; // @[axi_arbiter.scala 82:64 83:23 18:24]
  wire [31:0] _GEN_69 = state == 2'h3 ? io_lsu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_70 = state == 2'h3 & io_lsu_axi_in_arvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_71 = state == 2'h3 & io_lsu_axi_in_rready; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [31:0] _GEN_72 = state == 2'h3 ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_73 = state == 2'h3 & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [63:0] _GEN_74 = state == 2'h3 ? io_lsu_axi_in_wdata : 64'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [7:0] _GEN_75 = state == 2'h3 ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_76 = state == 2'h3 & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_77 = state == 2'h3 & io_lsu_axi_in_bready; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_78 = state == 2'h3 & io_axi_in_arready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire [63:0] _GEN_79 = state == 2'h3 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_80 = state == 2'h3 & io_axi_in_rvalid; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_81 = state == 2'h3 & io_axi_in_awready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_82 = state == 2'h3 & io_axi_in_wready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_83 = state == 2'h3 & io_axi_in_bvalid; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire [1:0] _GEN_90 = state == 2'h3 ? _GEN_68 : state; // @[axi_arbiter.scala 18:24 78:39]
  wire [31:0] _GEN_91 = state == 2'h2 ? io_lsu_axi_in_araddr : _GEN_69; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_92 = state == 2'h2 ? io_lsu_axi_in_arvalid : _GEN_70; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_93 = state == 2'h2 ? io_lsu_axi_in_rready : _GEN_71; // @[axi_arbiter.scala 70:39 71:24]
  wire [31:0] _GEN_94 = state == 2'h2 ? io_lsu_axi_in_awaddr : _GEN_72; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_95 = state == 2'h2 ? io_lsu_axi_in_awvalid : _GEN_73; // @[axi_arbiter.scala 70:39 71:24]
  wire [63:0] _GEN_96 = state == 2'h2 ? io_lsu_axi_in_wdata : _GEN_74; // @[axi_arbiter.scala 70:39 71:24]
  wire [7:0] _GEN_97 = state == 2'h2 ? io_lsu_axi_in_wstrb : _GEN_75; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_98 = state == 2'h2 ? io_lsu_axi_in_wvalid : _GEN_76; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_99 = state == 2'h2 ? io_lsu_axi_in_bready : _GEN_77; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_100 = state == 2'h2 ? io_axi_in_arready : _GEN_78; // @[axi_arbiter.scala 70:39 72:28]
  wire [63:0] _GEN_101 = state == 2'h2 ? io_axi_in_rdata : _GEN_79; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_102 = state == 2'h2 ? io_axi_in_rvalid : _GEN_80; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_103 = state == 2'h2 ? io_axi_in_awready : _GEN_81; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_104 = state == 2'h2 ? io_axi_in_wready : _GEN_82; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_105 = state == 2'h2 ? io_axi_in_bvalid : _GEN_83; // @[axi_arbiter.scala 70:39 72:28]
  wire [31:0] _GEN_113 = state == 2'h1 ? io_ifu_axi_in_araddr : _GEN_91; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_114 = state == 2'h1 ? io_ifu_axi_in_arvalid : _GEN_92; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_115 = state == 2'h1 ? io_ifu_axi_in_rready : _GEN_93; // @[axi_arbiter.scala 62:39 63:24]
  wire [31:0] _GEN_116 = state == 2'h1 ? 32'h0 : _GEN_94; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_117 = state == 2'h1 ? 1'h0 : _GEN_95; // @[axi_arbiter.scala 62:39 63:24]
  wire [63:0] _GEN_118 = state == 2'h1 ? 64'h0 : _GEN_96; // @[axi_arbiter.scala 62:39 63:24]
  wire [7:0] _GEN_119 = state == 2'h1 ? 8'h0 : _GEN_97; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_120 = state == 2'h1 ? 1'h0 : _GEN_98; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_121 = state == 2'h1 ? 1'h0 : _GEN_99; // @[axi_arbiter.scala 62:39 63:24]
  wire [63:0] _GEN_123 = state == 2'h1 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 62:39 64:28]
  wire  _GEN_124 = state == 2'h1 & io_axi_in_rvalid; // @[axi_arbiter.scala 62:39 64:28]
  wire  _GEN_128 = state == 2'h1 ? 1'h0 : _GEN_100; // @[axi_arbiter.scala 62:39 65:28]
  wire [63:0] _GEN_129 = state == 2'h1 ? 64'h0 : _GEN_101; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_130 = state == 2'h1 ? 1'h0 : _GEN_102; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_131 = state == 2'h1 ? 1'h0 : _GEN_103; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_132 = state == 2'h1 ? 1'h0 : _GEN_104; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_133 = state == 2'h1 ? 1'h0 : _GEN_105; // @[axi_arbiter.scala 62:39 65:28]
  assign io_ifu_axi_out_rdata = state == 2'h0 ? _GEN_61 : _GEN_123; // @[axi_arbiter.scala 40:27]
  assign io_ifu_axi_out_rvalid = state == 2'h0 ? _GEN_62 : _GEN_124; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_arready = state == 2'h0 ? _GEN_54 : _GEN_128; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_rdata = state == 2'h0 ? _GEN_55 : _GEN_129; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_rvalid = state == 2'h0 ? _GEN_56 : _GEN_130; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_awready = state == 2'h0 ? _GEN_57 : _GEN_131; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_wready = state == 2'h0 ? _GEN_58 : _GEN_132; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_bvalid = state == 2'h0 ? _GEN_59 : _GEN_133; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_araddr = state == 2'h0 ? _GEN_45 : _GEN_113; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_arvalid = state == 2'h0 ? _GEN_46 : _GEN_114; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_rready = state == 2'h0 ? _GEN_47 : _GEN_115; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_awaddr = state == 2'h0 ? _GEN_48 : _GEN_116; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_awvalid = state == 2'h0 ? _GEN_49 : _GEN_117; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wdata = state == 2'h0 ? _GEN_50 : _GEN_118; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wstrb = state == 2'h0 ? _GEN_51 : _GEN_119; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wvalid = state == 2'h0 ? _GEN_52 : _GEN_120; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_bready = state == 2'h0 ? _GEN_53 : _GEN_121; // @[axi_arbiter.scala 40:27]
  always @(posedge clock) begin
    if (reset) begin // @[axi_arbiter.scala 18:24]
      state <= 2'h0; // @[axi_arbiter.scala 18:24]
    end else if (state == 2'h0) begin // @[axi_arbiter.scala 40:27]
      if (io_lsu_axi_in_awvalid) begin // @[axi_arbiter.scala 41:40]
        state <= 2'h3; // @[axi_arbiter.scala 42:23]
      end else if (io_lsu_axi_in_arvalid) begin // @[axi_arbiter.scala 46:46]
        state <= 2'h2; // @[axi_arbiter.scala 47:23]
      end else begin
        state <= _GEN_0;
      end
    end else if (state == 2'h1) begin // @[axi_arbiter.scala 62:39]
      if (io_ifu_axi_out_rvalid & io_ifu_axi_in_rready) begin // @[axi_arbiter.scala 66:64]
        state <= 2'h0; // @[axi_arbiter.scala 67:23]
      end
    end else if (state == 2'h2) begin // @[axi_arbiter.scala 70:39]
      state <= _GEN_67;
    end else begin
      state <= _GEN_90;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU_AXI(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_pc_valid,
  output        io_inst_valid,
  output [31:0] io_inst,
  output [31:0] io_inst_reg,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  inst_ready; // @[IFU_AXI.scala 19:29]
  wire  _GEN_0 = io_axi_in_rvalid & inst_ready ? 1'h0 : 1'h1; // @[IFU_AXI.scala 20:41 21:20 23:20]
  reg [31:0] inst_reg; // @[IFU_AXI.scala 25:27]
  assign io_inst_valid = io_axi_in_rvalid; // @[IFU_AXI.scala 43:19]
  assign io_inst = io_axi_in_rdata[31:0]; // @[IFU_AXI.scala 41:31]
  assign io_inst_reg = inst_reg; // @[IFU_AXI.scala 42:17]
  assign io_axi_out_araddr = io_pc[31:0]; // @[IFU_AXI.scala 31:31]
  assign io_axi_out_arvalid = io_pc_valid; // @[IFU_AXI.scala 32:24]
  assign io_axi_out_rready = inst_ready; // @[IFU_AXI.scala 33:23]
  always @(posedge clock) begin
    inst_ready <= reset | _GEN_0; // @[IFU_AXI.scala 19:{29,29}]
    if (reset) begin // @[IFU_AXI.scala 25:27]
      inst_reg <= 32'h0; // @[IFU_AXI.scala 25:27]
    end else if (io_axi_in_rvalid) begin // @[IFU_AXI.scala 26:27]
      inst_reg <= io_axi_in_rdata[31:0]; // @[IFU_AXI.scala 27:18]
    end else if (io_pc_valid) begin // @[IFU_AXI.scala 28:28]
      inst_reg <= 32'h0; // @[IFU_AXI.scala 29:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst_ready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  inst_reg = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module I_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_ifu_araddr,
  input         io_from_ifu_arvalid,
  input         io_from_ifu_rready,
  output [63:0] io_to_ifu_rdata,
  output        io_to_ifu_rvalid,
  output [31:0] io_to_axi_araddr,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [63:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_0_0; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_1; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_2; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_3; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_4; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_5; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_6; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_7; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_8; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_9; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_10; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_11; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_12; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_13; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_14; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_15; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_16; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_17; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_18; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_19; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_20; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_21; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_22; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_23; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_24; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_25; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_26; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_27; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_28; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_29; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_30; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_31; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_32; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_33; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_34; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_35; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_36; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_37; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_38; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_39; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_40; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_41; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_42; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_43; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_44; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_45; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_46; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_47; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_48; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_49; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_50; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_51; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_52; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_53; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_54; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_55; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_56; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_57; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_58; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_59; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_60; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_61; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_62; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_63; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_64; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_65; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_66; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_67; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_68; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_69; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_70; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_71; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_72; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_73; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_74; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_75; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_76; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_77; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_78; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_79; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_80; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_81; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_82; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_83; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_84; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_85; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_86; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_87; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_88; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_89; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_90; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_91; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_92; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_93; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_94; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_95; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_96; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_97; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_98; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_99; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_100; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_101; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_102; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_103; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_104; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_105; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_106; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_107; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_108; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_109; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_110; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_111; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_112; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_113; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_114; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_115; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_116; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_117; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_118; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_119; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_120; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_121; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_122; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_123; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_124; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_125; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_126; // @[i_cache.scala 17:24]
  reg [63:0] ram_0_127; // @[i_cache.scala 17:24]
  reg [63:0] ram_1_0; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_1; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_2; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_3; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_4; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_5; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_6; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_7; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_8; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_9; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_10; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_11; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_12; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_13; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_14; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_15; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_16; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_17; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_18; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_19; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_20; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_21; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_22; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_23; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_24; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_25; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_26; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_27; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_28; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_29; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_30; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_31; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_32; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_33; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_34; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_35; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_36; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_37; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_38; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_39; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_40; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_41; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_42; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_43; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_44; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_45; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_46; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_47; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_48; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_49; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_50; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_51; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_52; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_53; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_54; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_55; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_56; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_57; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_58; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_59; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_60; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_61; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_62; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_63; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_64; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_65; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_66; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_67; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_68; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_69; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_70; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_71; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_72; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_73; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_74; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_75; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_76; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_77; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_78; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_79; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_80; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_81; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_82; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_83; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_84; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_85; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_86; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_87; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_88; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_89; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_90; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_91; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_92; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_93; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_94; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_95; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_96; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_97; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_98; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_99; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_100; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_101; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_102; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_103; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_104; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_105; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_106; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_107; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_108; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_109; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_110; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_111; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_112; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_113; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_114; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_115; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_116; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_117; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_118; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_119; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_120; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_121; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_122; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_123; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_124; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_125; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_126; // @[i_cache.scala 18:24]
  reg [63:0] ram_1_127; // @[i_cache.scala 18:24]
  reg [31:0] tag_0_0; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_1; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_2; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_3; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_4; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_5; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_6; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_7; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_8; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_9; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_10; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_11; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_12; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_13; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_14; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_15; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_16; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_17; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_18; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_19; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_20; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_21; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_22; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_23; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_24; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_25; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_26; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_27; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_28; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_29; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_30; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_31; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_32; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_33; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_34; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_35; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_36; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_37; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_38; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_39; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_40; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_41; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_42; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_43; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_44; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_45; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_46; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_47; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_48; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_49; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_50; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_51; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_52; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_53; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_54; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_55; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_56; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_57; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_58; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_59; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_60; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_61; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_62; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_63; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_64; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_65; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_66; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_67; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_68; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_69; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_70; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_71; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_72; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_73; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_74; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_75; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_76; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_77; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_78; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_79; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_80; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_81; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_82; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_83; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_84; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_85; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_86; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_87; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_88; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_89; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_90; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_91; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_92; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_93; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_94; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_95; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_96; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_97; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_98; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_99; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_100; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_101; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_102; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_103; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_104; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_105; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_106; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_107; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_108; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_109; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_110; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_111; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_112; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_113; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_114; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_115; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_116; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_117; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_118; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_119; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_120; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_121; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_122; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_123; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_124; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_125; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_126; // @[i_cache.scala 19:24]
  reg [31:0] tag_0_127; // @[i_cache.scala 19:24]
  reg [31:0] tag_1_0; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_1; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_2; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_3; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_4; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_5; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_6; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_7; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_8; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_9; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_10; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_11; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_12; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_13; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_14; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_15; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_16; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_17; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_18; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_19; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_20; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_21; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_22; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_23; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_24; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_25; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_26; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_27; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_28; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_29; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_30; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_31; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_32; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_33; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_34; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_35; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_36; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_37; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_38; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_39; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_40; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_41; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_42; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_43; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_44; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_45; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_46; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_47; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_48; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_49; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_50; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_51; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_52; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_53; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_54; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_55; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_56; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_57; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_58; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_59; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_60; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_61; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_62; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_63; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_64; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_65; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_66; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_67; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_68; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_69; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_70; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_71; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_72; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_73; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_74; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_75; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_76; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_77; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_78; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_79; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_80; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_81; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_82; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_83; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_84; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_85; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_86; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_87; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_88; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_89; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_90; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_91; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_92; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_93; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_94; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_95; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_96; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_97; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_98; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_99; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_100; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_101; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_102; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_103; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_104; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_105; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_106; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_107; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_108; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_109; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_110; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_111; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_112; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_113; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_114; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_115; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_116; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_117; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_118; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_119; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_120; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_121; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_122; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_123; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_124; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_125; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_126; // @[i_cache.scala 20:24]
  reg [31:0] tag_1_127; // @[i_cache.scala 20:24]
  reg  valid_0_0; // @[i_cache.scala 21:26]
  reg  valid_0_1; // @[i_cache.scala 21:26]
  reg  valid_0_2; // @[i_cache.scala 21:26]
  reg  valid_0_3; // @[i_cache.scala 21:26]
  reg  valid_0_4; // @[i_cache.scala 21:26]
  reg  valid_0_5; // @[i_cache.scala 21:26]
  reg  valid_0_6; // @[i_cache.scala 21:26]
  reg  valid_0_7; // @[i_cache.scala 21:26]
  reg  valid_0_8; // @[i_cache.scala 21:26]
  reg  valid_0_9; // @[i_cache.scala 21:26]
  reg  valid_0_10; // @[i_cache.scala 21:26]
  reg  valid_0_11; // @[i_cache.scala 21:26]
  reg  valid_0_12; // @[i_cache.scala 21:26]
  reg  valid_0_13; // @[i_cache.scala 21:26]
  reg  valid_0_14; // @[i_cache.scala 21:26]
  reg  valid_0_15; // @[i_cache.scala 21:26]
  reg  valid_0_16; // @[i_cache.scala 21:26]
  reg  valid_0_17; // @[i_cache.scala 21:26]
  reg  valid_0_18; // @[i_cache.scala 21:26]
  reg  valid_0_19; // @[i_cache.scala 21:26]
  reg  valid_0_20; // @[i_cache.scala 21:26]
  reg  valid_0_21; // @[i_cache.scala 21:26]
  reg  valid_0_22; // @[i_cache.scala 21:26]
  reg  valid_0_23; // @[i_cache.scala 21:26]
  reg  valid_0_24; // @[i_cache.scala 21:26]
  reg  valid_0_25; // @[i_cache.scala 21:26]
  reg  valid_0_26; // @[i_cache.scala 21:26]
  reg  valid_0_27; // @[i_cache.scala 21:26]
  reg  valid_0_28; // @[i_cache.scala 21:26]
  reg  valid_0_29; // @[i_cache.scala 21:26]
  reg  valid_0_30; // @[i_cache.scala 21:26]
  reg  valid_0_31; // @[i_cache.scala 21:26]
  reg  valid_0_32; // @[i_cache.scala 21:26]
  reg  valid_0_33; // @[i_cache.scala 21:26]
  reg  valid_0_34; // @[i_cache.scala 21:26]
  reg  valid_0_35; // @[i_cache.scala 21:26]
  reg  valid_0_36; // @[i_cache.scala 21:26]
  reg  valid_0_37; // @[i_cache.scala 21:26]
  reg  valid_0_38; // @[i_cache.scala 21:26]
  reg  valid_0_39; // @[i_cache.scala 21:26]
  reg  valid_0_40; // @[i_cache.scala 21:26]
  reg  valid_0_41; // @[i_cache.scala 21:26]
  reg  valid_0_42; // @[i_cache.scala 21:26]
  reg  valid_0_43; // @[i_cache.scala 21:26]
  reg  valid_0_44; // @[i_cache.scala 21:26]
  reg  valid_0_45; // @[i_cache.scala 21:26]
  reg  valid_0_46; // @[i_cache.scala 21:26]
  reg  valid_0_47; // @[i_cache.scala 21:26]
  reg  valid_0_48; // @[i_cache.scala 21:26]
  reg  valid_0_49; // @[i_cache.scala 21:26]
  reg  valid_0_50; // @[i_cache.scala 21:26]
  reg  valid_0_51; // @[i_cache.scala 21:26]
  reg  valid_0_52; // @[i_cache.scala 21:26]
  reg  valid_0_53; // @[i_cache.scala 21:26]
  reg  valid_0_54; // @[i_cache.scala 21:26]
  reg  valid_0_55; // @[i_cache.scala 21:26]
  reg  valid_0_56; // @[i_cache.scala 21:26]
  reg  valid_0_57; // @[i_cache.scala 21:26]
  reg  valid_0_58; // @[i_cache.scala 21:26]
  reg  valid_0_59; // @[i_cache.scala 21:26]
  reg  valid_0_60; // @[i_cache.scala 21:26]
  reg  valid_0_61; // @[i_cache.scala 21:26]
  reg  valid_0_62; // @[i_cache.scala 21:26]
  reg  valid_0_63; // @[i_cache.scala 21:26]
  reg  valid_0_64; // @[i_cache.scala 21:26]
  reg  valid_0_65; // @[i_cache.scala 21:26]
  reg  valid_0_66; // @[i_cache.scala 21:26]
  reg  valid_0_67; // @[i_cache.scala 21:26]
  reg  valid_0_68; // @[i_cache.scala 21:26]
  reg  valid_0_69; // @[i_cache.scala 21:26]
  reg  valid_0_70; // @[i_cache.scala 21:26]
  reg  valid_0_71; // @[i_cache.scala 21:26]
  reg  valid_0_72; // @[i_cache.scala 21:26]
  reg  valid_0_73; // @[i_cache.scala 21:26]
  reg  valid_0_74; // @[i_cache.scala 21:26]
  reg  valid_0_75; // @[i_cache.scala 21:26]
  reg  valid_0_76; // @[i_cache.scala 21:26]
  reg  valid_0_77; // @[i_cache.scala 21:26]
  reg  valid_0_78; // @[i_cache.scala 21:26]
  reg  valid_0_79; // @[i_cache.scala 21:26]
  reg  valid_0_80; // @[i_cache.scala 21:26]
  reg  valid_0_81; // @[i_cache.scala 21:26]
  reg  valid_0_82; // @[i_cache.scala 21:26]
  reg  valid_0_83; // @[i_cache.scala 21:26]
  reg  valid_0_84; // @[i_cache.scala 21:26]
  reg  valid_0_85; // @[i_cache.scala 21:26]
  reg  valid_0_86; // @[i_cache.scala 21:26]
  reg  valid_0_87; // @[i_cache.scala 21:26]
  reg  valid_0_88; // @[i_cache.scala 21:26]
  reg  valid_0_89; // @[i_cache.scala 21:26]
  reg  valid_0_90; // @[i_cache.scala 21:26]
  reg  valid_0_91; // @[i_cache.scala 21:26]
  reg  valid_0_92; // @[i_cache.scala 21:26]
  reg  valid_0_93; // @[i_cache.scala 21:26]
  reg  valid_0_94; // @[i_cache.scala 21:26]
  reg  valid_0_95; // @[i_cache.scala 21:26]
  reg  valid_0_96; // @[i_cache.scala 21:26]
  reg  valid_0_97; // @[i_cache.scala 21:26]
  reg  valid_0_98; // @[i_cache.scala 21:26]
  reg  valid_0_99; // @[i_cache.scala 21:26]
  reg  valid_0_100; // @[i_cache.scala 21:26]
  reg  valid_0_101; // @[i_cache.scala 21:26]
  reg  valid_0_102; // @[i_cache.scala 21:26]
  reg  valid_0_103; // @[i_cache.scala 21:26]
  reg  valid_0_104; // @[i_cache.scala 21:26]
  reg  valid_0_105; // @[i_cache.scala 21:26]
  reg  valid_0_106; // @[i_cache.scala 21:26]
  reg  valid_0_107; // @[i_cache.scala 21:26]
  reg  valid_0_108; // @[i_cache.scala 21:26]
  reg  valid_0_109; // @[i_cache.scala 21:26]
  reg  valid_0_110; // @[i_cache.scala 21:26]
  reg  valid_0_111; // @[i_cache.scala 21:26]
  reg  valid_0_112; // @[i_cache.scala 21:26]
  reg  valid_0_113; // @[i_cache.scala 21:26]
  reg  valid_0_114; // @[i_cache.scala 21:26]
  reg  valid_0_115; // @[i_cache.scala 21:26]
  reg  valid_0_116; // @[i_cache.scala 21:26]
  reg  valid_0_117; // @[i_cache.scala 21:26]
  reg  valid_0_118; // @[i_cache.scala 21:26]
  reg  valid_0_119; // @[i_cache.scala 21:26]
  reg  valid_0_120; // @[i_cache.scala 21:26]
  reg  valid_0_121; // @[i_cache.scala 21:26]
  reg  valid_0_122; // @[i_cache.scala 21:26]
  reg  valid_0_123; // @[i_cache.scala 21:26]
  reg  valid_0_124; // @[i_cache.scala 21:26]
  reg  valid_0_125; // @[i_cache.scala 21:26]
  reg  valid_0_126; // @[i_cache.scala 21:26]
  reg  valid_0_127; // @[i_cache.scala 21:26]
  reg  valid_1_0; // @[i_cache.scala 22:26]
  reg  valid_1_1; // @[i_cache.scala 22:26]
  reg  valid_1_2; // @[i_cache.scala 22:26]
  reg  valid_1_3; // @[i_cache.scala 22:26]
  reg  valid_1_4; // @[i_cache.scala 22:26]
  reg  valid_1_5; // @[i_cache.scala 22:26]
  reg  valid_1_6; // @[i_cache.scala 22:26]
  reg  valid_1_7; // @[i_cache.scala 22:26]
  reg  valid_1_8; // @[i_cache.scala 22:26]
  reg  valid_1_9; // @[i_cache.scala 22:26]
  reg  valid_1_10; // @[i_cache.scala 22:26]
  reg  valid_1_11; // @[i_cache.scala 22:26]
  reg  valid_1_12; // @[i_cache.scala 22:26]
  reg  valid_1_13; // @[i_cache.scala 22:26]
  reg  valid_1_14; // @[i_cache.scala 22:26]
  reg  valid_1_15; // @[i_cache.scala 22:26]
  reg  valid_1_16; // @[i_cache.scala 22:26]
  reg  valid_1_17; // @[i_cache.scala 22:26]
  reg  valid_1_18; // @[i_cache.scala 22:26]
  reg  valid_1_19; // @[i_cache.scala 22:26]
  reg  valid_1_20; // @[i_cache.scala 22:26]
  reg  valid_1_21; // @[i_cache.scala 22:26]
  reg  valid_1_22; // @[i_cache.scala 22:26]
  reg  valid_1_23; // @[i_cache.scala 22:26]
  reg  valid_1_24; // @[i_cache.scala 22:26]
  reg  valid_1_25; // @[i_cache.scala 22:26]
  reg  valid_1_26; // @[i_cache.scala 22:26]
  reg  valid_1_27; // @[i_cache.scala 22:26]
  reg  valid_1_28; // @[i_cache.scala 22:26]
  reg  valid_1_29; // @[i_cache.scala 22:26]
  reg  valid_1_30; // @[i_cache.scala 22:26]
  reg  valid_1_31; // @[i_cache.scala 22:26]
  reg  valid_1_32; // @[i_cache.scala 22:26]
  reg  valid_1_33; // @[i_cache.scala 22:26]
  reg  valid_1_34; // @[i_cache.scala 22:26]
  reg  valid_1_35; // @[i_cache.scala 22:26]
  reg  valid_1_36; // @[i_cache.scala 22:26]
  reg  valid_1_37; // @[i_cache.scala 22:26]
  reg  valid_1_38; // @[i_cache.scala 22:26]
  reg  valid_1_39; // @[i_cache.scala 22:26]
  reg  valid_1_40; // @[i_cache.scala 22:26]
  reg  valid_1_41; // @[i_cache.scala 22:26]
  reg  valid_1_42; // @[i_cache.scala 22:26]
  reg  valid_1_43; // @[i_cache.scala 22:26]
  reg  valid_1_44; // @[i_cache.scala 22:26]
  reg  valid_1_45; // @[i_cache.scala 22:26]
  reg  valid_1_46; // @[i_cache.scala 22:26]
  reg  valid_1_47; // @[i_cache.scala 22:26]
  reg  valid_1_48; // @[i_cache.scala 22:26]
  reg  valid_1_49; // @[i_cache.scala 22:26]
  reg  valid_1_50; // @[i_cache.scala 22:26]
  reg  valid_1_51; // @[i_cache.scala 22:26]
  reg  valid_1_52; // @[i_cache.scala 22:26]
  reg  valid_1_53; // @[i_cache.scala 22:26]
  reg  valid_1_54; // @[i_cache.scala 22:26]
  reg  valid_1_55; // @[i_cache.scala 22:26]
  reg  valid_1_56; // @[i_cache.scala 22:26]
  reg  valid_1_57; // @[i_cache.scala 22:26]
  reg  valid_1_58; // @[i_cache.scala 22:26]
  reg  valid_1_59; // @[i_cache.scala 22:26]
  reg  valid_1_60; // @[i_cache.scala 22:26]
  reg  valid_1_61; // @[i_cache.scala 22:26]
  reg  valid_1_62; // @[i_cache.scala 22:26]
  reg  valid_1_63; // @[i_cache.scala 22:26]
  reg  valid_1_64; // @[i_cache.scala 22:26]
  reg  valid_1_65; // @[i_cache.scala 22:26]
  reg  valid_1_66; // @[i_cache.scala 22:26]
  reg  valid_1_67; // @[i_cache.scala 22:26]
  reg  valid_1_68; // @[i_cache.scala 22:26]
  reg  valid_1_69; // @[i_cache.scala 22:26]
  reg  valid_1_70; // @[i_cache.scala 22:26]
  reg  valid_1_71; // @[i_cache.scala 22:26]
  reg  valid_1_72; // @[i_cache.scala 22:26]
  reg  valid_1_73; // @[i_cache.scala 22:26]
  reg  valid_1_74; // @[i_cache.scala 22:26]
  reg  valid_1_75; // @[i_cache.scala 22:26]
  reg  valid_1_76; // @[i_cache.scala 22:26]
  reg  valid_1_77; // @[i_cache.scala 22:26]
  reg  valid_1_78; // @[i_cache.scala 22:26]
  reg  valid_1_79; // @[i_cache.scala 22:26]
  reg  valid_1_80; // @[i_cache.scala 22:26]
  reg  valid_1_81; // @[i_cache.scala 22:26]
  reg  valid_1_82; // @[i_cache.scala 22:26]
  reg  valid_1_83; // @[i_cache.scala 22:26]
  reg  valid_1_84; // @[i_cache.scala 22:26]
  reg  valid_1_85; // @[i_cache.scala 22:26]
  reg  valid_1_86; // @[i_cache.scala 22:26]
  reg  valid_1_87; // @[i_cache.scala 22:26]
  reg  valid_1_88; // @[i_cache.scala 22:26]
  reg  valid_1_89; // @[i_cache.scala 22:26]
  reg  valid_1_90; // @[i_cache.scala 22:26]
  reg  valid_1_91; // @[i_cache.scala 22:26]
  reg  valid_1_92; // @[i_cache.scala 22:26]
  reg  valid_1_93; // @[i_cache.scala 22:26]
  reg  valid_1_94; // @[i_cache.scala 22:26]
  reg  valid_1_95; // @[i_cache.scala 22:26]
  reg  valid_1_96; // @[i_cache.scala 22:26]
  reg  valid_1_97; // @[i_cache.scala 22:26]
  reg  valid_1_98; // @[i_cache.scala 22:26]
  reg  valid_1_99; // @[i_cache.scala 22:26]
  reg  valid_1_100; // @[i_cache.scala 22:26]
  reg  valid_1_101; // @[i_cache.scala 22:26]
  reg  valid_1_102; // @[i_cache.scala 22:26]
  reg  valid_1_103; // @[i_cache.scala 22:26]
  reg  valid_1_104; // @[i_cache.scala 22:26]
  reg  valid_1_105; // @[i_cache.scala 22:26]
  reg  valid_1_106; // @[i_cache.scala 22:26]
  reg  valid_1_107; // @[i_cache.scala 22:26]
  reg  valid_1_108; // @[i_cache.scala 22:26]
  reg  valid_1_109; // @[i_cache.scala 22:26]
  reg  valid_1_110; // @[i_cache.scala 22:26]
  reg  valid_1_111; // @[i_cache.scala 22:26]
  reg  valid_1_112; // @[i_cache.scala 22:26]
  reg  valid_1_113; // @[i_cache.scala 22:26]
  reg  valid_1_114; // @[i_cache.scala 22:26]
  reg  valid_1_115; // @[i_cache.scala 22:26]
  reg  valid_1_116; // @[i_cache.scala 22:26]
  reg  valid_1_117; // @[i_cache.scala 22:26]
  reg  valid_1_118; // @[i_cache.scala 22:26]
  reg  valid_1_119; // @[i_cache.scala 22:26]
  reg  valid_1_120; // @[i_cache.scala 22:26]
  reg  valid_1_121; // @[i_cache.scala 22:26]
  reg  valid_1_122; // @[i_cache.scala 22:26]
  reg  valid_1_123; // @[i_cache.scala 22:26]
  reg  valid_1_124; // @[i_cache.scala 22:26]
  reg  valid_1_125; // @[i_cache.scala 22:26]
  reg  valid_1_126; // @[i_cache.scala 22:26]
  reg  valid_1_127; // @[i_cache.scala 22:26]
  reg  way0_hit; // @[i_cache.scala 23:27]
  reg  way1_hit; // @[i_cache.scala 24:27]
  reg [1:0] unuse_way; // @[i_cache.scala 26:28]
  reg [63:0] receive_data; // @[i_cache.scala 27:31]
  reg  quene; // @[i_cache.scala 28:24]
  wire [6:0] index = io_from_ifu_araddr[6:0]; // @[i_cache.scala 31:35]
  wire [24:0] tag = io_from_ifu_araddr[31:7]; // @[i_cache.scala 32:33]
  wire [31:0] _GEN_1 = 7'h1 == index ? tag_0_1 : tag_0_0; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_2 = 7'h2 == index ? tag_0_2 : _GEN_1; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_3 = 7'h3 == index ? tag_0_3 : _GEN_2; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_4 = 7'h4 == index ? tag_0_4 : _GEN_3; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_5 = 7'h5 == index ? tag_0_5 : _GEN_4; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_6 = 7'h6 == index ? tag_0_6 : _GEN_5; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_7 = 7'h7 == index ? tag_0_7 : _GEN_6; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_8 = 7'h8 == index ? tag_0_8 : _GEN_7; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_9 = 7'h9 == index ? tag_0_9 : _GEN_8; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_10 = 7'ha == index ? tag_0_10 : _GEN_9; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_11 = 7'hb == index ? tag_0_11 : _GEN_10; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_12 = 7'hc == index ? tag_0_12 : _GEN_11; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_13 = 7'hd == index ? tag_0_13 : _GEN_12; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_14 = 7'he == index ? tag_0_14 : _GEN_13; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_15 = 7'hf == index ? tag_0_15 : _GEN_14; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_16 = 7'h10 == index ? tag_0_16 : _GEN_15; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_17 = 7'h11 == index ? tag_0_17 : _GEN_16; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_18 = 7'h12 == index ? tag_0_18 : _GEN_17; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_19 = 7'h13 == index ? tag_0_19 : _GEN_18; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_20 = 7'h14 == index ? tag_0_20 : _GEN_19; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_21 = 7'h15 == index ? tag_0_21 : _GEN_20; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_22 = 7'h16 == index ? tag_0_22 : _GEN_21; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_23 = 7'h17 == index ? tag_0_23 : _GEN_22; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_24 = 7'h18 == index ? tag_0_24 : _GEN_23; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_25 = 7'h19 == index ? tag_0_25 : _GEN_24; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_26 = 7'h1a == index ? tag_0_26 : _GEN_25; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_27 = 7'h1b == index ? tag_0_27 : _GEN_26; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_28 = 7'h1c == index ? tag_0_28 : _GEN_27; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_29 = 7'h1d == index ? tag_0_29 : _GEN_28; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_30 = 7'h1e == index ? tag_0_30 : _GEN_29; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_31 = 7'h1f == index ? tag_0_31 : _GEN_30; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_32 = 7'h20 == index ? tag_0_32 : _GEN_31; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_33 = 7'h21 == index ? tag_0_33 : _GEN_32; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_34 = 7'h22 == index ? tag_0_34 : _GEN_33; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_35 = 7'h23 == index ? tag_0_35 : _GEN_34; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_36 = 7'h24 == index ? tag_0_36 : _GEN_35; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_37 = 7'h25 == index ? tag_0_37 : _GEN_36; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_38 = 7'h26 == index ? tag_0_38 : _GEN_37; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_39 = 7'h27 == index ? tag_0_39 : _GEN_38; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_40 = 7'h28 == index ? tag_0_40 : _GEN_39; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_41 = 7'h29 == index ? tag_0_41 : _GEN_40; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_42 = 7'h2a == index ? tag_0_42 : _GEN_41; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_43 = 7'h2b == index ? tag_0_43 : _GEN_42; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_44 = 7'h2c == index ? tag_0_44 : _GEN_43; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_45 = 7'h2d == index ? tag_0_45 : _GEN_44; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_46 = 7'h2e == index ? tag_0_46 : _GEN_45; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_47 = 7'h2f == index ? tag_0_47 : _GEN_46; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_48 = 7'h30 == index ? tag_0_48 : _GEN_47; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_49 = 7'h31 == index ? tag_0_49 : _GEN_48; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_50 = 7'h32 == index ? tag_0_50 : _GEN_49; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_51 = 7'h33 == index ? tag_0_51 : _GEN_50; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_52 = 7'h34 == index ? tag_0_52 : _GEN_51; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_53 = 7'h35 == index ? tag_0_53 : _GEN_52; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_54 = 7'h36 == index ? tag_0_54 : _GEN_53; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_55 = 7'h37 == index ? tag_0_55 : _GEN_54; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_56 = 7'h38 == index ? tag_0_56 : _GEN_55; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_57 = 7'h39 == index ? tag_0_57 : _GEN_56; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_58 = 7'h3a == index ? tag_0_58 : _GEN_57; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_59 = 7'h3b == index ? tag_0_59 : _GEN_58; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_60 = 7'h3c == index ? tag_0_60 : _GEN_59; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_61 = 7'h3d == index ? tag_0_61 : _GEN_60; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_62 = 7'h3e == index ? tag_0_62 : _GEN_61; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_63 = 7'h3f == index ? tag_0_63 : _GEN_62; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_64 = 7'h40 == index ? tag_0_64 : _GEN_63; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_65 = 7'h41 == index ? tag_0_65 : _GEN_64; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_66 = 7'h42 == index ? tag_0_66 : _GEN_65; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_67 = 7'h43 == index ? tag_0_67 : _GEN_66; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_68 = 7'h44 == index ? tag_0_68 : _GEN_67; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_69 = 7'h45 == index ? tag_0_69 : _GEN_68; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_70 = 7'h46 == index ? tag_0_70 : _GEN_69; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_71 = 7'h47 == index ? tag_0_71 : _GEN_70; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_72 = 7'h48 == index ? tag_0_72 : _GEN_71; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_73 = 7'h49 == index ? tag_0_73 : _GEN_72; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_74 = 7'h4a == index ? tag_0_74 : _GEN_73; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_75 = 7'h4b == index ? tag_0_75 : _GEN_74; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_76 = 7'h4c == index ? tag_0_76 : _GEN_75; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_77 = 7'h4d == index ? tag_0_77 : _GEN_76; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_78 = 7'h4e == index ? tag_0_78 : _GEN_77; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_79 = 7'h4f == index ? tag_0_79 : _GEN_78; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_80 = 7'h50 == index ? tag_0_80 : _GEN_79; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_81 = 7'h51 == index ? tag_0_81 : _GEN_80; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_82 = 7'h52 == index ? tag_0_82 : _GEN_81; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_83 = 7'h53 == index ? tag_0_83 : _GEN_82; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_84 = 7'h54 == index ? tag_0_84 : _GEN_83; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_85 = 7'h55 == index ? tag_0_85 : _GEN_84; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_86 = 7'h56 == index ? tag_0_86 : _GEN_85; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_87 = 7'h57 == index ? tag_0_87 : _GEN_86; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_88 = 7'h58 == index ? tag_0_88 : _GEN_87; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_89 = 7'h59 == index ? tag_0_89 : _GEN_88; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_90 = 7'h5a == index ? tag_0_90 : _GEN_89; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_91 = 7'h5b == index ? tag_0_91 : _GEN_90; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_92 = 7'h5c == index ? tag_0_92 : _GEN_91; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_93 = 7'h5d == index ? tag_0_93 : _GEN_92; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_94 = 7'h5e == index ? tag_0_94 : _GEN_93; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_95 = 7'h5f == index ? tag_0_95 : _GEN_94; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_96 = 7'h60 == index ? tag_0_96 : _GEN_95; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_97 = 7'h61 == index ? tag_0_97 : _GEN_96; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_98 = 7'h62 == index ? tag_0_98 : _GEN_97; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_99 = 7'h63 == index ? tag_0_99 : _GEN_98; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_100 = 7'h64 == index ? tag_0_100 : _GEN_99; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_101 = 7'h65 == index ? tag_0_101 : _GEN_100; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_102 = 7'h66 == index ? tag_0_102 : _GEN_101; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_103 = 7'h67 == index ? tag_0_103 : _GEN_102; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_104 = 7'h68 == index ? tag_0_104 : _GEN_103; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_105 = 7'h69 == index ? tag_0_105 : _GEN_104; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_106 = 7'h6a == index ? tag_0_106 : _GEN_105; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_107 = 7'h6b == index ? tag_0_107 : _GEN_106; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_108 = 7'h6c == index ? tag_0_108 : _GEN_107; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_109 = 7'h6d == index ? tag_0_109 : _GEN_108; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_110 = 7'h6e == index ? tag_0_110 : _GEN_109; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_111 = 7'h6f == index ? tag_0_111 : _GEN_110; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_112 = 7'h70 == index ? tag_0_112 : _GEN_111; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_113 = 7'h71 == index ? tag_0_113 : _GEN_112; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_114 = 7'h72 == index ? tag_0_114 : _GEN_113; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_115 = 7'h73 == index ? tag_0_115 : _GEN_114; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_116 = 7'h74 == index ? tag_0_116 : _GEN_115; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_117 = 7'h75 == index ? tag_0_117 : _GEN_116; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_118 = 7'h76 == index ? tag_0_118 : _GEN_117; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_119 = 7'h77 == index ? tag_0_119 : _GEN_118; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_120 = 7'h78 == index ? tag_0_120 : _GEN_119; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_121 = 7'h79 == index ? tag_0_121 : _GEN_120; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_122 = 7'h7a == index ? tag_0_122 : _GEN_121; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_123 = 7'h7b == index ? tag_0_123 : _GEN_122; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_124 = 7'h7c == index ? tag_0_124 : _GEN_123; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_125 = 7'h7d == index ? tag_0_125 : _GEN_124; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_126 = 7'h7e == index ? tag_0_126 : _GEN_125; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_127 = 7'h7f == index ? tag_0_127 : _GEN_126; // @[i_cache.scala 34:{24,24}]
  wire [31:0] _GEN_7706 = {{7'd0}, tag}; // @[i_cache.scala 34:24]
  wire  _GEN_129 = 7'h1 == index ? valid_0_1 : valid_0_0; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_130 = 7'h2 == index ? valid_0_2 : _GEN_129; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_131 = 7'h3 == index ? valid_0_3 : _GEN_130; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_132 = 7'h4 == index ? valid_0_4 : _GEN_131; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_133 = 7'h5 == index ? valid_0_5 : _GEN_132; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_134 = 7'h6 == index ? valid_0_6 : _GEN_133; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_135 = 7'h7 == index ? valid_0_7 : _GEN_134; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_136 = 7'h8 == index ? valid_0_8 : _GEN_135; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_137 = 7'h9 == index ? valid_0_9 : _GEN_136; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_138 = 7'ha == index ? valid_0_10 : _GEN_137; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_139 = 7'hb == index ? valid_0_11 : _GEN_138; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_140 = 7'hc == index ? valid_0_12 : _GEN_139; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_141 = 7'hd == index ? valid_0_13 : _GEN_140; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_142 = 7'he == index ? valid_0_14 : _GEN_141; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_143 = 7'hf == index ? valid_0_15 : _GEN_142; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_144 = 7'h10 == index ? valid_0_16 : _GEN_143; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_145 = 7'h11 == index ? valid_0_17 : _GEN_144; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_146 = 7'h12 == index ? valid_0_18 : _GEN_145; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_147 = 7'h13 == index ? valid_0_19 : _GEN_146; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_148 = 7'h14 == index ? valid_0_20 : _GEN_147; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_149 = 7'h15 == index ? valid_0_21 : _GEN_148; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_150 = 7'h16 == index ? valid_0_22 : _GEN_149; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_151 = 7'h17 == index ? valid_0_23 : _GEN_150; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_152 = 7'h18 == index ? valid_0_24 : _GEN_151; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_153 = 7'h19 == index ? valid_0_25 : _GEN_152; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_154 = 7'h1a == index ? valid_0_26 : _GEN_153; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_155 = 7'h1b == index ? valid_0_27 : _GEN_154; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_156 = 7'h1c == index ? valid_0_28 : _GEN_155; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_157 = 7'h1d == index ? valid_0_29 : _GEN_156; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_158 = 7'h1e == index ? valid_0_30 : _GEN_157; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_159 = 7'h1f == index ? valid_0_31 : _GEN_158; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_160 = 7'h20 == index ? valid_0_32 : _GEN_159; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_161 = 7'h21 == index ? valid_0_33 : _GEN_160; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_162 = 7'h22 == index ? valid_0_34 : _GEN_161; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_163 = 7'h23 == index ? valid_0_35 : _GEN_162; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_164 = 7'h24 == index ? valid_0_36 : _GEN_163; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_165 = 7'h25 == index ? valid_0_37 : _GEN_164; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_166 = 7'h26 == index ? valid_0_38 : _GEN_165; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_167 = 7'h27 == index ? valid_0_39 : _GEN_166; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_168 = 7'h28 == index ? valid_0_40 : _GEN_167; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_169 = 7'h29 == index ? valid_0_41 : _GEN_168; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_170 = 7'h2a == index ? valid_0_42 : _GEN_169; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_171 = 7'h2b == index ? valid_0_43 : _GEN_170; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_172 = 7'h2c == index ? valid_0_44 : _GEN_171; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_173 = 7'h2d == index ? valid_0_45 : _GEN_172; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_174 = 7'h2e == index ? valid_0_46 : _GEN_173; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_175 = 7'h2f == index ? valid_0_47 : _GEN_174; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_176 = 7'h30 == index ? valid_0_48 : _GEN_175; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_177 = 7'h31 == index ? valid_0_49 : _GEN_176; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_178 = 7'h32 == index ? valid_0_50 : _GEN_177; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_179 = 7'h33 == index ? valid_0_51 : _GEN_178; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_180 = 7'h34 == index ? valid_0_52 : _GEN_179; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_181 = 7'h35 == index ? valid_0_53 : _GEN_180; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_182 = 7'h36 == index ? valid_0_54 : _GEN_181; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_183 = 7'h37 == index ? valid_0_55 : _GEN_182; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_184 = 7'h38 == index ? valid_0_56 : _GEN_183; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_185 = 7'h39 == index ? valid_0_57 : _GEN_184; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_186 = 7'h3a == index ? valid_0_58 : _GEN_185; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_187 = 7'h3b == index ? valid_0_59 : _GEN_186; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_188 = 7'h3c == index ? valid_0_60 : _GEN_187; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_189 = 7'h3d == index ? valid_0_61 : _GEN_188; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_190 = 7'h3e == index ? valid_0_62 : _GEN_189; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_191 = 7'h3f == index ? valid_0_63 : _GEN_190; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_192 = 7'h40 == index ? valid_0_64 : _GEN_191; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_193 = 7'h41 == index ? valid_0_65 : _GEN_192; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_194 = 7'h42 == index ? valid_0_66 : _GEN_193; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_195 = 7'h43 == index ? valid_0_67 : _GEN_194; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_196 = 7'h44 == index ? valid_0_68 : _GEN_195; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_197 = 7'h45 == index ? valid_0_69 : _GEN_196; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_198 = 7'h46 == index ? valid_0_70 : _GEN_197; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_199 = 7'h47 == index ? valid_0_71 : _GEN_198; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_200 = 7'h48 == index ? valid_0_72 : _GEN_199; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_201 = 7'h49 == index ? valid_0_73 : _GEN_200; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_202 = 7'h4a == index ? valid_0_74 : _GEN_201; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_203 = 7'h4b == index ? valid_0_75 : _GEN_202; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_204 = 7'h4c == index ? valid_0_76 : _GEN_203; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_205 = 7'h4d == index ? valid_0_77 : _GEN_204; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_206 = 7'h4e == index ? valid_0_78 : _GEN_205; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_207 = 7'h4f == index ? valid_0_79 : _GEN_206; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_208 = 7'h50 == index ? valid_0_80 : _GEN_207; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_209 = 7'h51 == index ? valid_0_81 : _GEN_208; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_210 = 7'h52 == index ? valid_0_82 : _GEN_209; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_211 = 7'h53 == index ? valid_0_83 : _GEN_210; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_212 = 7'h54 == index ? valid_0_84 : _GEN_211; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_213 = 7'h55 == index ? valid_0_85 : _GEN_212; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_214 = 7'h56 == index ? valid_0_86 : _GEN_213; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_215 = 7'h57 == index ? valid_0_87 : _GEN_214; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_216 = 7'h58 == index ? valid_0_88 : _GEN_215; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_217 = 7'h59 == index ? valid_0_89 : _GEN_216; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_218 = 7'h5a == index ? valid_0_90 : _GEN_217; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_219 = 7'h5b == index ? valid_0_91 : _GEN_218; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_220 = 7'h5c == index ? valid_0_92 : _GEN_219; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_221 = 7'h5d == index ? valid_0_93 : _GEN_220; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_222 = 7'h5e == index ? valid_0_94 : _GEN_221; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_223 = 7'h5f == index ? valid_0_95 : _GEN_222; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_224 = 7'h60 == index ? valid_0_96 : _GEN_223; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_225 = 7'h61 == index ? valid_0_97 : _GEN_224; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_226 = 7'h62 == index ? valid_0_98 : _GEN_225; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_227 = 7'h63 == index ? valid_0_99 : _GEN_226; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_228 = 7'h64 == index ? valid_0_100 : _GEN_227; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_229 = 7'h65 == index ? valid_0_101 : _GEN_228; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_230 = 7'h66 == index ? valid_0_102 : _GEN_229; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_231 = 7'h67 == index ? valid_0_103 : _GEN_230; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_232 = 7'h68 == index ? valid_0_104 : _GEN_231; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_233 = 7'h69 == index ? valid_0_105 : _GEN_232; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_234 = 7'h6a == index ? valid_0_106 : _GEN_233; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_235 = 7'h6b == index ? valid_0_107 : _GEN_234; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_236 = 7'h6c == index ? valid_0_108 : _GEN_235; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_237 = 7'h6d == index ? valid_0_109 : _GEN_236; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_238 = 7'h6e == index ? valid_0_110 : _GEN_237; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_239 = 7'h6f == index ? valid_0_111 : _GEN_238; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_240 = 7'h70 == index ? valid_0_112 : _GEN_239; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_241 = 7'h71 == index ? valid_0_113 : _GEN_240; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_242 = 7'h72 == index ? valid_0_114 : _GEN_241; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_243 = 7'h73 == index ? valid_0_115 : _GEN_242; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_244 = 7'h74 == index ? valid_0_116 : _GEN_243; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_245 = 7'h75 == index ? valid_0_117 : _GEN_244; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_246 = 7'h76 == index ? valid_0_118 : _GEN_245; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_247 = 7'h77 == index ? valid_0_119 : _GEN_246; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_248 = 7'h78 == index ? valid_0_120 : _GEN_247; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_249 = 7'h79 == index ? valid_0_121 : _GEN_248; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_250 = 7'h7a == index ? valid_0_122 : _GEN_249; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_251 = 7'h7b == index ? valid_0_123 : _GEN_250; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_252 = 7'h7c == index ? valid_0_124 : _GEN_251; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_253 = 7'h7d == index ? valid_0_125 : _GEN_252; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_254 = 7'h7e == index ? valid_0_126 : _GEN_253; // @[i_cache.scala 34:{50,50}]
  wire  _GEN_255 = 7'h7f == index ? valid_0_127 : _GEN_254; // @[i_cache.scala 34:{50,50}]
  wire  _T_2 = _GEN_127 == _GEN_7706 & _GEN_255; // @[i_cache.scala 34:33]
  wire [31:0] _GEN_258 = 7'h1 == index ? tag_1_1 : tag_1_0; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_259 = 7'h2 == index ? tag_1_2 : _GEN_258; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_260 = 7'h3 == index ? tag_1_3 : _GEN_259; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_261 = 7'h4 == index ? tag_1_4 : _GEN_260; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_262 = 7'h5 == index ? tag_1_5 : _GEN_261; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_263 = 7'h6 == index ? tag_1_6 : _GEN_262; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_264 = 7'h7 == index ? tag_1_7 : _GEN_263; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_265 = 7'h8 == index ? tag_1_8 : _GEN_264; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_266 = 7'h9 == index ? tag_1_9 : _GEN_265; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_267 = 7'ha == index ? tag_1_10 : _GEN_266; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_268 = 7'hb == index ? tag_1_11 : _GEN_267; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_269 = 7'hc == index ? tag_1_12 : _GEN_268; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_270 = 7'hd == index ? tag_1_13 : _GEN_269; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_271 = 7'he == index ? tag_1_14 : _GEN_270; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_272 = 7'hf == index ? tag_1_15 : _GEN_271; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_273 = 7'h10 == index ? tag_1_16 : _GEN_272; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_274 = 7'h11 == index ? tag_1_17 : _GEN_273; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_275 = 7'h12 == index ? tag_1_18 : _GEN_274; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_276 = 7'h13 == index ? tag_1_19 : _GEN_275; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_277 = 7'h14 == index ? tag_1_20 : _GEN_276; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_278 = 7'h15 == index ? tag_1_21 : _GEN_277; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_279 = 7'h16 == index ? tag_1_22 : _GEN_278; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_280 = 7'h17 == index ? tag_1_23 : _GEN_279; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_281 = 7'h18 == index ? tag_1_24 : _GEN_280; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_282 = 7'h19 == index ? tag_1_25 : _GEN_281; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_283 = 7'h1a == index ? tag_1_26 : _GEN_282; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_284 = 7'h1b == index ? tag_1_27 : _GEN_283; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_285 = 7'h1c == index ? tag_1_28 : _GEN_284; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_286 = 7'h1d == index ? tag_1_29 : _GEN_285; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_287 = 7'h1e == index ? tag_1_30 : _GEN_286; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_288 = 7'h1f == index ? tag_1_31 : _GEN_287; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_289 = 7'h20 == index ? tag_1_32 : _GEN_288; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_290 = 7'h21 == index ? tag_1_33 : _GEN_289; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_291 = 7'h22 == index ? tag_1_34 : _GEN_290; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_292 = 7'h23 == index ? tag_1_35 : _GEN_291; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_293 = 7'h24 == index ? tag_1_36 : _GEN_292; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_294 = 7'h25 == index ? tag_1_37 : _GEN_293; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_295 = 7'h26 == index ? tag_1_38 : _GEN_294; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_296 = 7'h27 == index ? tag_1_39 : _GEN_295; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_297 = 7'h28 == index ? tag_1_40 : _GEN_296; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_298 = 7'h29 == index ? tag_1_41 : _GEN_297; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_299 = 7'h2a == index ? tag_1_42 : _GEN_298; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_300 = 7'h2b == index ? tag_1_43 : _GEN_299; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_301 = 7'h2c == index ? tag_1_44 : _GEN_300; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_302 = 7'h2d == index ? tag_1_45 : _GEN_301; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_303 = 7'h2e == index ? tag_1_46 : _GEN_302; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_304 = 7'h2f == index ? tag_1_47 : _GEN_303; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_305 = 7'h30 == index ? tag_1_48 : _GEN_304; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_306 = 7'h31 == index ? tag_1_49 : _GEN_305; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_307 = 7'h32 == index ? tag_1_50 : _GEN_306; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_308 = 7'h33 == index ? tag_1_51 : _GEN_307; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_309 = 7'h34 == index ? tag_1_52 : _GEN_308; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_310 = 7'h35 == index ? tag_1_53 : _GEN_309; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_311 = 7'h36 == index ? tag_1_54 : _GEN_310; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_312 = 7'h37 == index ? tag_1_55 : _GEN_311; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_313 = 7'h38 == index ? tag_1_56 : _GEN_312; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_314 = 7'h39 == index ? tag_1_57 : _GEN_313; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_315 = 7'h3a == index ? tag_1_58 : _GEN_314; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_316 = 7'h3b == index ? tag_1_59 : _GEN_315; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_317 = 7'h3c == index ? tag_1_60 : _GEN_316; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_318 = 7'h3d == index ? tag_1_61 : _GEN_317; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_319 = 7'h3e == index ? tag_1_62 : _GEN_318; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_320 = 7'h3f == index ? tag_1_63 : _GEN_319; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_321 = 7'h40 == index ? tag_1_64 : _GEN_320; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_322 = 7'h41 == index ? tag_1_65 : _GEN_321; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_323 = 7'h42 == index ? tag_1_66 : _GEN_322; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_324 = 7'h43 == index ? tag_1_67 : _GEN_323; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_325 = 7'h44 == index ? tag_1_68 : _GEN_324; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_326 = 7'h45 == index ? tag_1_69 : _GEN_325; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_327 = 7'h46 == index ? tag_1_70 : _GEN_326; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_328 = 7'h47 == index ? tag_1_71 : _GEN_327; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_329 = 7'h48 == index ? tag_1_72 : _GEN_328; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_330 = 7'h49 == index ? tag_1_73 : _GEN_329; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_331 = 7'h4a == index ? tag_1_74 : _GEN_330; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_332 = 7'h4b == index ? tag_1_75 : _GEN_331; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_333 = 7'h4c == index ? tag_1_76 : _GEN_332; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_334 = 7'h4d == index ? tag_1_77 : _GEN_333; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_335 = 7'h4e == index ? tag_1_78 : _GEN_334; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_336 = 7'h4f == index ? tag_1_79 : _GEN_335; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_337 = 7'h50 == index ? tag_1_80 : _GEN_336; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_338 = 7'h51 == index ? tag_1_81 : _GEN_337; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_339 = 7'h52 == index ? tag_1_82 : _GEN_338; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_340 = 7'h53 == index ? tag_1_83 : _GEN_339; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_341 = 7'h54 == index ? tag_1_84 : _GEN_340; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_342 = 7'h55 == index ? tag_1_85 : _GEN_341; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_343 = 7'h56 == index ? tag_1_86 : _GEN_342; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_344 = 7'h57 == index ? tag_1_87 : _GEN_343; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_345 = 7'h58 == index ? tag_1_88 : _GEN_344; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_346 = 7'h59 == index ? tag_1_89 : _GEN_345; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_347 = 7'h5a == index ? tag_1_90 : _GEN_346; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_348 = 7'h5b == index ? tag_1_91 : _GEN_347; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_349 = 7'h5c == index ? tag_1_92 : _GEN_348; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_350 = 7'h5d == index ? tag_1_93 : _GEN_349; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_351 = 7'h5e == index ? tag_1_94 : _GEN_350; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_352 = 7'h5f == index ? tag_1_95 : _GEN_351; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_353 = 7'h60 == index ? tag_1_96 : _GEN_352; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_354 = 7'h61 == index ? tag_1_97 : _GEN_353; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_355 = 7'h62 == index ? tag_1_98 : _GEN_354; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_356 = 7'h63 == index ? tag_1_99 : _GEN_355; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_357 = 7'h64 == index ? tag_1_100 : _GEN_356; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_358 = 7'h65 == index ? tag_1_101 : _GEN_357; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_359 = 7'h66 == index ? tag_1_102 : _GEN_358; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_360 = 7'h67 == index ? tag_1_103 : _GEN_359; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_361 = 7'h68 == index ? tag_1_104 : _GEN_360; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_362 = 7'h69 == index ? tag_1_105 : _GEN_361; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_363 = 7'h6a == index ? tag_1_106 : _GEN_362; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_364 = 7'h6b == index ? tag_1_107 : _GEN_363; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_365 = 7'h6c == index ? tag_1_108 : _GEN_364; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_366 = 7'h6d == index ? tag_1_109 : _GEN_365; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_367 = 7'h6e == index ? tag_1_110 : _GEN_366; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_368 = 7'h6f == index ? tag_1_111 : _GEN_367; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_369 = 7'h70 == index ? tag_1_112 : _GEN_368; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_370 = 7'h71 == index ? tag_1_113 : _GEN_369; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_371 = 7'h72 == index ? tag_1_114 : _GEN_370; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_372 = 7'h73 == index ? tag_1_115 : _GEN_371; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_373 = 7'h74 == index ? tag_1_116 : _GEN_372; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_374 = 7'h75 == index ? tag_1_117 : _GEN_373; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_375 = 7'h76 == index ? tag_1_118 : _GEN_374; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_376 = 7'h77 == index ? tag_1_119 : _GEN_375; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_377 = 7'h78 == index ? tag_1_120 : _GEN_376; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_378 = 7'h79 == index ? tag_1_121 : _GEN_377; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_379 = 7'h7a == index ? tag_1_122 : _GEN_378; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_380 = 7'h7b == index ? tag_1_123 : _GEN_379; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_381 = 7'h7c == index ? tag_1_124 : _GEN_380; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_382 = 7'h7d == index ? tag_1_125 : _GEN_381; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_383 = 7'h7e == index ? tag_1_126 : _GEN_382; // @[i_cache.scala 39:{24,24}]
  wire [31:0] _GEN_384 = 7'h7f == index ? tag_1_127 : _GEN_383; // @[i_cache.scala 39:{24,24}]
  wire  _GEN_386 = 7'h1 == index ? valid_1_1 : valid_1_0; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_387 = 7'h2 == index ? valid_1_2 : _GEN_386; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_388 = 7'h3 == index ? valid_1_3 : _GEN_387; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_389 = 7'h4 == index ? valid_1_4 : _GEN_388; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_390 = 7'h5 == index ? valid_1_5 : _GEN_389; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_391 = 7'h6 == index ? valid_1_6 : _GEN_390; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_392 = 7'h7 == index ? valid_1_7 : _GEN_391; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_393 = 7'h8 == index ? valid_1_8 : _GEN_392; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_394 = 7'h9 == index ? valid_1_9 : _GEN_393; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_395 = 7'ha == index ? valid_1_10 : _GEN_394; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_396 = 7'hb == index ? valid_1_11 : _GEN_395; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_397 = 7'hc == index ? valid_1_12 : _GEN_396; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_398 = 7'hd == index ? valid_1_13 : _GEN_397; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_399 = 7'he == index ? valid_1_14 : _GEN_398; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_400 = 7'hf == index ? valid_1_15 : _GEN_399; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_401 = 7'h10 == index ? valid_1_16 : _GEN_400; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_402 = 7'h11 == index ? valid_1_17 : _GEN_401; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_403 = 7'h12 == index ? valid_1_18 : _GEN_402; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_404 = 7'h13 == index ? valid_1_19 : _GEN_403; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_405 = 7'h14 == index ? valid_1_20 : _GEN_404; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_406 = 7'h15 == index ? valid_1_21 : _GEN_405; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_407 = 7'h16 == index ? valid_1_22 : _GEN_406; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_408 = 7'h17 == index ? valid_1_23 : _GEN_407; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_409 = 7'h18 == index ? valid_1_24 : _GEN_408; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_410 = 7'h19 == index ? valid_1_25 : _GEN_409; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_411 = 7'h1a == index ? valid_1_26 : _GEN_410; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_412 = 7'h1b == index ? valid_1_27 : _GEN_411; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_413 = 7'h1c == index ? valid_1_28 : _GEN_412; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_414 = 7'h1d == index ? valid_1_29 : _GEN_413; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_415 = 7'h1e == index ? valid_1_30 : _GEN_414; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_416 = 7'h1f == index ? valid_1_31 : _GEN_415; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_417 = 7'h20 == index ? valid_1_32 : _GEN_416; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_418 = 7'h21 == index ? valid_1_33 : _GEN_417; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_419 = 7'h22 == index ? valid_1_34 : _GEN_418; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_420 = 7'h23 == index ? valid_1_35 : _GEN_419; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_421 = 7'h24 == index ? valid_1_36 : _GEN_420; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_422 = 7'h25 == index ? valid_1_37 : _GEN_421; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_423 = 7'h26 == index ? valid_1_38 : _GEN_422; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_424 = 7'h27 == index ? valid_1_39 : _GEN_423; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_425 = 7'h28 == index ? valid_1_40 : _GEN_424; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_426 = 7'h29 == index ? valid_1_41 : _GEN_425; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_427 = 7'h2a == index ? valid_1_42 : _GEN_426; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_428 = 7'h2b == index ? valid_1_43 : _GEN_427; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_429 = 7'h2c == index ? valid_1_44 : _GEN_428; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_430 = 7'h2d == index ? valid_1_45 : _GEN_429; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_431 = 7'h2e == index ? valid_1_46 : _GEN_430; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_432 = 7'h2f == index ? valid_1_47 : _GEN_431; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_433 = 7'h30 == index ? valid_1_48 : _GEN_432; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_434 = 7'h31 == index ? valid_1_49 : _GEN_433; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_435 = 7'h32 == index ? valid_1_50 : _GEN_434; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_436 = 7'h33 == index ? valid_1_51 : _GEN_435; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_437 = 7'h34 == index ? valid_1_52 : _GEN_436; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_438 = 7'h35 == index ? valid_1_53 : _GEN_437; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_439 = 7'h36 == index ? valid_1_54 : _GEN_438; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_440 = 7'h37 == index ? valid_1_55 : _GEN_439; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_441 = 7'h38 == index ? valid_1_56 : _GEN_440; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_442 = 7'h39 == index ? valid_1_57 : _GEN_441; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_443 = 7'h3a == index ? valid_1_58 : _GEN_442; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_444 = 7'h3b == index ? valid_1_59 : _GEN_443; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_445 = 7'h3c == index ? valid_1_60 : _GEN_444; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_446 = 7'h3d == index ? valid_1_61 : _GEN_445; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_447 = 7'h3e == index ? valid_1_62 : _GEN_446; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_448 = 7'h3f == index ? valid_1_63 : _GEN_447; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_449 = 7'h40 == index ? valid_1_64 : _GEN_448; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_450 = 7'h41 == index ? valid_1_65 : _GEN_449; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_451 = 7'h42 == index ? valid_1_66 : _GEN_450; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_452 = 7'h43 == index ? valid_1_67 : _GEN_451; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_453 = 7'h44 == index ? valid_1_68 : _GEN_452; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_454 = 7'h45 == index ? valid_1_69 : _GEN_453; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_455 = 7'h46 == index ? valid_1_70 : _GEN_454; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_456 = 7'h47 == index ? valid_1_71 : _GEN_455; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_457 = 7'h48 == index ? valid_1_72 : _GEN_456; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_458 = 7'h49 == index ? valid_1_73 : _GEN_457; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_459 = 7'h4a == index ? valid_1_74 : _GEN_458; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_460 = 7'h4b == index ? valid_1_75 : _GEN_459; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_461 = 7'h4c == index ? valid_1_76 : _GEN_460; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_462 = 7'h4d == index ? valid_1_77 : _GEN_461; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_463 = 7'h4e == index ? valid_1_78 : _GEN_462; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_464 = 7'h4f == index ? valid_1_79 : _GEN_463; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_465 = 7'h50 == index ? valid_1_80 : _GEN_464; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_466 = 7'h51 == index ? valid_1_81 : _GEN_465; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_467 = 7'h52 == index ? valid_1_82 : _GEN_466; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_468 = 7'h53 == index ? valid_1_83 : _GEN_467; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_469 = 7'h54 == index ? valid_1_84 : _GEN_468; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_470 = 7'h55 == index ? valid_1_85 : _GEN_469; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_471 = 7'h56 == index ? valid_1_86 : _GEN_470; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_472 = 7'h57 == index ? valid_1_87 : _GEN_471; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_473 = 7'h58 == index ? valid_1_88 : _GEN_472; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_474 = 7'h59 == index ? valid_1_89 : _GEN_473; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_475 = 7'h5a == index ? valid_1_90 : _GEN_474; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_476 = 7'h5b == index ? valid_1_91 : _GEN_475; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_477 = 7'h5c == index ? valid_1_92 : _GEN_476; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_478 = 7'h5d == index ? valid_1_93 : _GEN_477; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_479 = 7'h5e == index ? valid_1_94 : _GEN_478; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_480 = 7'h5f == index ? valid_1_95 : _GEN_479; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_481 = 7'h60 == index ? valid_1_96 : _GEN_480; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_482 = 7'h61 == index ? valid_1_97 : _GEN_481; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_483 = 7'h62 == index ? valid_1_98 : _GEN_482; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_484 = 7'h63 == index ? valid_1_99 : _GEN_483; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_485 = 7'h64 == index ? valid_1_100 : _GEN_484; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_486 = 7'h65 == index ? valid_1_101 : _GEN_485; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_487 = 7'h66 == index ? valid_1_102 : _GEN_486; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_488 = 7'h67 == index ? valid_1_103 : _GEN_487; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_489 = 7'h68 == index ? valid_1_104 : _GEN_488; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_490 = 7'h69 == index ? valid_1_105 : _GEN_489; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_491 = 7'h6a == index ? valid_1_106 : _GEN_490; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_492 = 7'h6b == index ? valid_1_107 : _GEN_491; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_493 = 7'h6c == index ? valid_1_108 : _GEN_492; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_494 = 7'h6d == index ? valid_1_109 : _GEN_493; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_495 = 7'h6e == index ? valid_1_110 : _GEN_494; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_496 = 7'h6f == index ? valid_1_111 : _GEN_495; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_497 = 7'h70 == index ? valid_1_112 : _GEN_496; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_498 = 7'h71 == index ? valid_1_113 : _GEN_497; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_499 = 7'h72 == index ? valid_1_114 : _GEN_498; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_500 = 7'h73 == index ? valid_1_115 : _GEN_499; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_501 = 7'h74 == index ? valid_1_116 : _GEN_500; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_502 = 7'h75 == index ? valid_1_117 : _GEN_501; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_503 = 7'h76 == index ? valid_1_118 : _GEN_502; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_504 = 7'h77 == index ? valid_1_119 : _GEN_503; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_505 = 7'h78 == index ? valid_1_120 : _GEN_504; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_506 = 7'h79 == index ? valid_1_121 : _GEN_505; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_507 = 7'h7a == index ? valid_1_122 : _GEN_506; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_508 = 7'h7b == index ? valid_1_123 : _GEN_507; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_509 = 7'h7c == index ? valid_1_124 : _GEN_508; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_510 = 7'h7d == index ? valid_1_125 : _GEN_509; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_511 = 7'h7e == index ? valid_1_126 : _GEN_510; // @[i_cache.scala 39:{50,50}]
  wire  _GEN_512 = 7'h7f == index ? valid_1_127 : _GEN_511; // @[i_cache.scala 39:{50,50}]
  wire  _T_5 = _GEN_384 == _GEN_7706 & _GEN_512; // @[i_cache.scala 39:33]
  reg [2:0] state; // @[i_cache.scala 53:24]
  wire [2:0] _GEN_517 = io_from_ifu_rready ? 3'h0 : state; // @[i_cache.scala 53:24 64:41 65:27]
  wire [2:0] _GEN_518 = way1_hit ? _GEN_517 : 3'h2; // @[i_cache.scala 68:33 73:23]
  wire [2:0] _GEN_520 = io_from_axi_rvalid ? 3'h3 : state; // @[i_cache.scala 77:37 78:23 53:24]
  wire [63:0] _GEN_521 = io_from_axi_rvalid ? io_from_axi_rdata : receive_data; // @[i_cache.scala 80:37 81:30 27:31]
  wire [63:0] _GEN_522 = 7'h0 == index ? receive_data : ram_0_0; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_523 = 7'h1 == index ? receive_data : ram_0_1; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_524 = 7'h2 == index ? receive_data : ram_0_2; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_525 = 7'h3 == index ? receive_data : ram_0_3; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_526 = 7'h4 == index ? receive_data : ram_0_4; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_527 = 7'h5 == index ? receive_data : ram_0_5; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_528 = 7'h6 == index ? receive_data : ram_0_6; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_529 = 7'h7 == index ? receive_data : ram_0_7; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_530 = 7'h8 == index ? receive_data : ram_0_8; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_531 = 7'h9 == index ? receive_data : ram_0_9; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_532 = 7'ha == index ? receive_data : ram_0_10; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_533 = 7'hb == index ? receive_data : ram_0_11; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_534 = 7'hc == index ? receive_data : ram_0_12; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_535 = 7'hd == index ? receive_data : ram_0_13; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_536 = 7'he == index ? receive_data : ram_0_14; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_537 = 7'hf == index ? receive_data : ram_0_15; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_538 = 7'h10 == index ? receive_data : ram_0_16; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_539 = 7'h11 == index ? receive_data : ram_0_17; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_540 = 7'h12 == index ? receive_data : ram_0_18; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_541 = 7'h13 == index ? receive_data : ram_0_19; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_542 = 7'h14 == index ? receive_data : ram_0_20; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_543 = 7'h15 == index ? receive_data : ram_0_21; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_544 = 7'h16 == index ? receive_data : ram_0_22; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_545 = 7'h17 == index ? receive_data : ram_0_23; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_546 = 7'h18 == index ? receive_data : ram_0_24; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_547 = 7'h19 == index ? receive_data : ram_0_25; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_548 = 7'h1a == index ? receive_data : ram_0_26; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_549 = 7'h1b == index ? receive_data : ram_0_27; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_550 = 7'h1c == index ? receive_data : ram_0_28; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_551 = 7'h1d == index ? receive_data : ram_0_29; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_552 = 7'h1e == index ? receive_data : ram_0_30; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_553 = 7'h1f == index ? receive_data : ram_0_31; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_554 = 7'h20 == index ? receive_data : ram_0_32; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_555 = 7'h21 == index ? receive_data : ram_0_33; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_556 = 7'h22 == index ? receive_data : ram_0_34; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_557 = 7'h23 == index ? receive_data : ram_0_35; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_558 = 7'h24 == index ? receive_data : ram_0_36; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_559 = 7'h25 == index ? receive_data : ram_0_37; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_560 = 7'h26 == index ? receive_data : ram_0_38; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_561 = 7'h27 == index ? receive_data : ram_0_39; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_562 = 7'h28 == index ? receive_data : ram_0_40; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_563 = 7'h29 == index ? receive_data : ram_0_41; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_564 = 7'h2a == index ? receive_data : ram_0_42; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_565 = 7'h2b == index ? receive_data : ram_0_43; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_566 = 7'h2c == index ? receive_data : ram_0_44; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_567 = 7'h2d == index ? receive_data : ram_0_45; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_568 = 7'h2e == index ? receive_data : ram_0_46; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_569 = 7'h2f == index ? receive_data : ram_0_47; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_570 = 7'h30 == index ? receive_data : ram_0_48; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_571 = 7'h31 == index ? receive_data : ram_0_49; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_572 = 7'h32 == index ? receive_data : ram_0_50; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_573 = 7'h33 == index ? receive_data : ram_0_51; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_574 = 7'h34 == index ? receive_data : ram_0_52; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_575 = 7'h35 == index ? receive_data : ram_0_53; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_576 = 7'h36 == index ? receive_data : ram_0_54; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_577 = 7'h37 == index ? receive_data : ram_0_55; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_578 = 7'h38 == index ? receive_data : ram_0_56; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_579 = 7'h39 == index ? receive_data : ram_0_57; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_580 = 7'h3a == index ? receive_data : ram_0_58; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_581 = 7'h3b == index ? receive_data : ram_0_59; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_582 = 7'h3c == index ? receive_data : ram_0_60; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_583 = 7'h3d == index ? receive_data : ram_0_61; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_584 = 7'h3e == index ? receive_data : ram_0_62; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_585 = 7'h3f == index ? receive_data : ram_0_63; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_586 = 7'h40 == index ? receive_data : ram_0_64; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_587 = 7'h41 == index ? receive_data : ram_0_65; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_588 = 7'h42 == index ? receive_data : ram_0_66; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_589 = 7'h43 == index ? receive_data : ram_0_67; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_590 = 7'h44 == index ? receive_data : ram_0_68; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_591 = 7'h45 == index ? receive_data : ram_0_69; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_592 = 7'h46 == index ? receive_data : ram_0_70; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_593 = 7'h47 == index ? receive_data : ram_0_71; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_594 = 7'h48 == index ? receive_data : ram_0_72; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_595 = 7'h49 == index ? receive_data : ram_0_73; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_596 = 7'h4a == index ? receive_data : ram_0_74; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_597 = 7'h4b == index ? receive_data : ram_0_75; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_598 = 7'h4c == index ? receive_data : ram_0_76; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_599 = 7'h4d == index ? receive_data : ram_0_77; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_600 = 7'h4e == index ? receive_data : ram_0_78; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_601 = 7'h4f == index ? receive_data : ram_0_79; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_602 = 7'h50 == index ? receive_data : ram_0_80; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_603 = 7'h51 == index ? receive_data : ram_0_81; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_604 = 7'h52 == index ? receive_data : ram_0_82; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_605 = 7'h53 == index ? receive_data : ram_0_83; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_606 = 7'h54 == index ? receive_data : ram_0_84; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_607 = 7'h55 == index ? receive_data : ram_0_85; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_608 = 7'h56 == index ? receive_data : ram_0_86; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_609 = 7'h57 == index ? receive_data : ram_0_87; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_610 = 7'h58 == index ? receive_data : ram_0_88; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_611 = 7'h59 == index ? receive_data : ram_0_89; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_612 = 7'h5a == index ? receive_data : ram_0_90; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_613 = 7'h5b == index ? receive_data : ram_0_91; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_614 = 7'h5c == index ? receive_data : ram_0_92; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_615 = 7'h5d == index ? receive_data : ram_0_93; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_616 = 7'h5e == index ? receive_data : ram_0_94; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_617 = 7'h5f == index ? receive_data : ram_0_95; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_618 = 7'h60 == index ? receive_data : ram_0_96; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_619 = 7'h61 == index ? receive_data : ram_0_97; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_620 = 7'h62 == index ? receive_data : ram_0_98; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_621 = 7'h63 == index ? receive_data : ram_0_99; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_622 = 7'h64 == index ? receive_data : ram_0_100; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_623 = 7'h65 == index ? receive_data : ram_0_101; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_624 = 7'h66 == index ? receive_data : ram_0_102; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_625 = 7'h67 == index ? receive_data : ram_0_103; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_626 = 7'h68 == index ? receive_data : ram_0_104; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_627 = 7'h69 == index ? receive_data : ram_0_105; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_628 = 7'h6a == index ? receive_data : ram_0_106; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_629 = 7'h6b == index ? receive_data : ram_0_107; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_630 = 7'h6c == index ? receive_data : ram_0_108; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_631 = 7'h6d == index ? receive_data : ram_0_109; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_632 = 7'h6e == index ? receive_data : ram_0_110; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_633 = 7'h6f == index ? receive_data : ram_0_111; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_634 = 7'h70 == index ? receive_data : ram_0_112; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_635 = 7'h71 == index ? receive_data : ram_0_113; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_636 = 7'h72 == index ? receive_data : ram_0_114; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_637 = 7'h73 == index ? receive_data : ram_0_115; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_638 = 7'h74 == index ? receive_data : ram_0_116; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_639 = 7'h75 == index ? receive_data : ram_0_117; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_640 = 7'h76 == index ? receive_data : ram_0_118; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_641 = 7'h77 == index ? receive_data : ram_0_119; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_642 = 7'h78 == index ? receive_data : ram_0_120; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_643 = 7'h79 == index ? receive_data : ram_0_121; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_644 = 7'h7a == index ? receive_data : ram_0_122; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_645 = 7'h7b == index ? receive_data : ram_0_123; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_646 = 7'h7c == index ? receive_data : ram_0_124; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_647 = 7'h7d == index ? receive_data : ram_0_125; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_648 = 7'h7e == index ? receive_data : ram_0_126; // @[i_cache.scala 17:24 87:{30,30}]
  wire [63:0] _GEN_649 = 7'h7f == index ? receive_data : ram_0_127; // @[i_cache.scala 17:24 87:{30,30}]
  wire [31:0] _GEN_650 = 7'h0 == index ? _GEN_7706 : tag_0_0; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_651 = 7'h1 == index ? _GEN_7706 : tag_0_1; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_652 = 7'h2 == index ? _GEN_7706 : tag_0_2; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_653 = 7'h3 == index ? _GEN_7706 : tag_0_3; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_654 = 7'h4 == index ? _GEN_7706 : tag_0_4; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_655 = 7'h5 == index ? _GEN_7706 : tag_0_5; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_656 = 7'h6 == index ? _GEN_7706 : tag_0_6; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_657 = 7'h7 == index ? _GEN_7706 : tag_0_7; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_658 = 7'h8 == index ? _GEN_7706 : tag_0_8; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_659 = 7'h9 == index ? _GEN_7706 : tag_0_9; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_660 = 7'ha == index ? _GEN_7706 : tag_0_10; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_661 = 7'hb == index ? _GEN_7706 : tag_0_11; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_662 = 7'hc == index ? _GEN_7706 : tag_0_12; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_663 = 7'hd == index ? _GEN_7706 : tag_0_13; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_664 = 7'he == index ? _GEN_7706 : tag_0_14; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_665 = 7'hf == index ? _GEN_7706 : tag_0_15; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_666 = 7'h10 == index ? _GEN_7706 : tag_0_16; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_667 = 7'h11 == index ? _GEN_7706 : tag_0_17; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_668 = 7'h12 == index ? _GEN_7706 : tag_0_18; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_669 = 7'h13 == index ? _GEN_7706 : tag_0_19; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_670 = 7'h14 == index ? _GEN_7706 : tag_0_20; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_671 = 7'h15 == index ? _GEN_7706 : tag_0_21; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_672 = 7'h16 == index ? _GEN_7706 : tag_0_22; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_673 = 7'h17 == index ? _GEN_7706 : tag_0_23; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_674 = 7'h18 == index ? _GEN_7706 : tag_0_24; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_675 = 7'h19 == index ? _GEN_7706 : tag_0_25; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_676 = 7'h1a == index ? _GEN_7706 : tag_0_26; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_677 = 7'h1b == index ? _GEN_7706 : tag_0_27; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_678 = 7'h1c == index ? _GEN_7706 : tag_0_28; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_679 = 7'h1d == index ? _GEN_7706 : tag_0_29; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_680 = 7'h1e == index ? _GEN_7706 : tag_0_30; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_681 = 7'h1f == index ? _GEN_7706 : tag_0_31; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_682 = 7'h20 == index ? _GEN_7706 : tag_0_32; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_683 = 7'h21 == index ? _GEN_7706 : tag_0_33; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_684 = 7'h22 == index ? _GEN_7706 : tag_0_34; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_685 = 7'h23 == index ? _GEN_7706 : tag_0_35; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_686 = 7'h24 == index ? _GEN_7706 : tag_0_36; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_687 = 7'h25 == index ? _GEN_7706 : tag_0_37; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_688 = 7'h26 == index ? _GEN_7706 : tag_0_38; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_689 = 7'h27 == index ? _GEN_7706 : tag_0_39; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_690 = 7'h28 == index ? _GEN_7706 : tag_0_40; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_691 = 7'h29 == index ? _GEN_7706 : tag_0_41; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_692 = 7'h2a == index ? _GEN_7706 : tag_0_42; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_693 = 7'h2b == index ? _GEN_7706 : tag_0_43; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_694 = 7'h2c == index ? _GEN_7706 : tag_0_44; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_695 = 7'h2d == index ? _GEN_7706 : tag_0_45; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_696 = 7'h2e == index ? _GEN_7706 : tag_0_46; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_697 = 7'h2f == index ? _GEN_7706 : tag_0_47; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_698 = 7'h30 == index ? _GEN_7706 : tag_0_48; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_699 = 7'h31 == index ? _GEN_7706 : tag_0_49; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_700 = 7'h32 == index ? _GEN_7706 : tag_0_50; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_701 = 7'h33 == index ? _GEN_7706 : tag_0_51; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_702 = 7'h34 == index ? _GEN_7706 : tag_0_52; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_703 = 7'h35 == index ? _GEN_7706 : tag_0_53; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_704 = 7'h36 == index ? _GEN_7706 : tag_0_54; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_705 = 7'h37 == index ? _GEN_7706 : tag_0_55; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_706 = 7'h38 == index ? _GEN_7706 : tag_0_56; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_707 = 7'h39 == index ? _GEN_7706 : tag_0_57; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_708 = 7'h3a == index ? _GEN_7706 : tag_0_58; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_709 = 7'h3b == index ? _GEN_7706 : tag_0_59; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_710 = 7'h3c == index ? _GEN_7706 : tag_0_60; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_711 = 7'h3d == index ? _GEN_7706 : tag_0_61; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_712 = 7'h3e == index ? _GEN_7706 : tag_0_62; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_713 = 7'h3f == index ? _GEN_7706 : tag_0_63; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_714 = 7'h40 == index ? _GEN_7706 : tag_0_64; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_715 = 7'h41 == index ? _GEN_7706 : tag_0_65; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_716 = 7'h42 == index ? _GEN_7706 : tag_0_66; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_717 = 7'h43 == index ? _GEN_7706 : tag_0_67; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_718 = 7'h44 == index ? _GEN_7706 : tag_0_68; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_719 = 7'h45 == index ? _GEN_7706 : tag_0_69; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_720 = 7'h46 == index ? _GEN_7706 : tag_0_70; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_721 = 7'h47 == index ? _GEN_7706 : tag_0_71; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_722 = 7'h48 == index ? _GEN_7706 : tag_0_72; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_723 = 7'h49 == index ? _GEN_7706 : tag_0_73; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_724 = 7'h4a == index ? _GEN_7706 : tag_0_74; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_725 = 7'h4b == index ? _GEN_7706 : tag_0_75; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_726 = 7'h4c == index ? _GEN_7706 : tag_0_76; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_727 = 7'h4d == index ? _GEN_7706 : tag_0_77; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_728 = 7'h4e == index ? _GEN_7706 : tag_0_78; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_729 = 7'h4f == index ? _GEN_7706 : tag_0_79; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_730 = 7'h50 == index ? _GEN_7706 : tag_0_80; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_731 = 7'h51 == index ? _GEN_7706 : tag_0_81; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_732 = 7'h52 == index ? _GEN_7706 : tag_0_82; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_733 = 7'h53 == index ? _GEN_7706 : tag_0_83; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_734 = 7'h54 == index ? _GEN_7706 : tag_0_84; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_735 = 7'h55 == index ? _GEN_7706 : tag_0_85; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_736 = 7'h56 == index ? _GEN_7706 : tag_0_86; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_737 = 7'h57 == index ? _GEN_7706 : tag_0_87; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_738 = 7'h58 == index ? _GEN_7706 : tag_0_88; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_739 = 7'h59 == index ? _GEN_7706 : tag_0_89; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_740 = 7'h5a == index ? _GEN_7706 : tag_0_90; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_741 = 7'h5b == index ? _GEN_7706 : tag_0_91; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_742 = 7'h5c == index ? _GEN_7706 : tag_0_92; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_743 = 7'h5d == index ? _GEN_7706 : tag_0_93; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_744 = 7'h5e == index ? _GEN_7706 : tag_0_94; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_745 = 7'h5f == index ? _GEN_7706 : tag_0_95; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_746 = 7'h60 == index ? _GEN_7706 : tag_0_96; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_747 = 7'h61 == index ? _GEN_7706 : tag_0_97; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_748 = 7'h62 == index ? _GEN_7706 : tag_0_98; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_749 = 7'h63 == index ? _GEN_7706 : tag_0_99; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_750 = 7'h64 == index ? _GEN_7706 : tag_0_100; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_751 = 7'h65 == index ? _GEN_7706 : tag_0_101; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_752 = 7'h66 == index ? _GEN_7706 : tag_0_102; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_753 = 7'h67 == index ? _GEN_7706 : tag_0_103; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_754 = 7'h68 == index ? _GEN_7706 : tag_0_104; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_755 = 7'h69 == index ? _GEN_7706 : tag_0_105; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_756 = 7'h6a == index ? _GEN_7706 : tag_0_106; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_757 = 7'h6b == index ? _GEN_7706 : tag_0_107; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_758 = 7'h6c == index ? _GEN_7706 : tag_0_108; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_759 = 7'h6d == index ? _GEN_7706 : tag_0_109; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_760 = 7'h6e == index ? _GEN_7706 : tag_0_110; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_761 = 7'h6f == index ? _GEN_7706 : tag_0_111; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_762 = 7'h70 == index ? _GEN_7706 : tag_0_112; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_763 = 7'h71 == index ? _GEN_7706 : tag_0_113; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_764 = 7'h72 == index ? _GEN_7706 : tag_0_114; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_765 = 7'h73 == index ? _GEN_7706 : tag_0_115; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_766 = 7'h74 == index ? _GEN_7706 : tag_0_116; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_767 = 7'h75 == index ? _GEN_7706 : tag_0_117; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_768 = 7'h76 == index ? _GEN_7706 : tag_0_118; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_769 = 7'h77 == index ? _GEN_7706 : tag_0_119; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_770 = 7'h78 == index ? _GEN_7706 : tag_0_120; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_771 = 7'h79 == index ? _GEN_7706 : tag_0_121; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_772 = 7'h7a == index ? _GEN_7706 : tag_0_122; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_773 = 7'h7b == index ? _GEN_7706 : tag_0_123; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_774 = 7'h7c == index ? _GEN_7706 : tag_0_124; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_775 = 7'h7d == index ? _GEN_7706 : tag_0_125; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_776 = 7'h7e == index ? _GEN_7706 : tag_0_126; // @[i_cache.scala 19:24 88:{30,30}]
  wire [31:0] _GEN_777 = 7'h7f == index ? _GEN_7706 : tag_0_127; // @[i_cache.scala 19:24 88:{30,30}]
  wire  _GEN_7710 = 7'h0 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_778 = 7'h0 == index | valid_0_0; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7712 = 7'h1 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_779 = 7'h1 == index | valid_0_1; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7714 = 7'h2 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_780 = 7'h2 == index | valid_0_2; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7718 = 7'h3 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_781 = 7'h3 == index | valid_0_3; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7727 = 7'h4 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_782 = 7'h4 == index | valid_0_4; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7729 = 7'h5 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_783 = 7'h5 == index | valid_0_5; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7731 = 7'h6 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_784 = 7'h6 == index | valid_0_6; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7733 = 7'h7 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_785 = 7'h7 == index | valid_0_7; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7738 = 7'h8 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_786 = 7'h8 == index | valid_0_8; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7739 = 7'h9 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_787 = 7'h9 == index | valid_0_9; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7740 = 7'ha == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_788 = 7'ha == index | valid_0_10; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7741 = 7'hb == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_789 = 7'hb == index | valid_0_11; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7742 = 7'hc == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_790 = 7'hc == index | valid_0_12; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7743 = 7'hd == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_791 = 7'hd == index | valid_0_13; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7744 = 7'he == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_792 = 7'he == index | valid_0_14; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7745 = 7'hf == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_793 = 7'hf == index | valid_0_15; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7746 = 7'h10 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_794 = 7'h10 == index | valid_0_16; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7747 = 7'h11 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_795 = 7'h11 == index | valid_0_17; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7748 = 7'h12 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_796 = 7'h12 == index | valid_0_18; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7749 = 7'h13 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_797 = 7'h13 == index | valid_0_19; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7750 = 7'h14 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_798 = 7'h14 == index | valid_0_20; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7751 = 7'h15 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_799 = 7'h15 == index | valid_0_21; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7752 = 7'h16 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_800 = 7'h16 == index | valid_0_22; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7753 = 7'h17 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_801 = 7'h17 == index | valid_0_23; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7754 = 7'h18 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_802 = 7'h18 == index | valid_0_24; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7755 = 7'h19 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_803 = 7'h19 == index | valid_0_25; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7756 = 7'h1a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_804 = 7'h1a == index | valid_0_26; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7757 = 7'h1b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_805 = 7'h1b == index | valid_0_27; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7758 = 7'h1c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_806 = 7'h1c == index | valid_0_28; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7759 = 7'h1d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_807 = 7'h1d == index | valid_0_29; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7760 = 7'h1e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_808 = 7'h1e == index | valid_0_30; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7761 = 7'h1f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_809 = 7'h1f == index | valid_0_31; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7762 = 7'h20 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_810 = 7'h20 == index | valid_0_32; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7763 = 7'h21 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_811 = 7'h21 == index | valid_0_33; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7764 = 7'h22 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_812 = 7'h22 == index | valid_0_34; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7765 = 7'h23 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_813 = 7'h23 == index | valid_0_35; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7766 = 7'h24 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_814 = 7'h24 == index | valid_0_36; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7767 = 7'h25 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_815 = 7'h25 == index | valid_0_37; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7768 = 7'h26 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_816 = 7'h26 == index | valid_0_38; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7769 = 7'h27 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_817 = 7'h27 == index | valid_0_39; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7770 = 7'h28 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_818 = 7'h28 == index | valid_0_40; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7771 = 7'h29 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_819 = 7'h29 == index | valid_0_41; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7772 = 7'h2a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_820 = 7'h2a == index | valid_0_42; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7773 = 7'h2b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_821 = 7'h2b == index | valid_0_43; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7774 = 7'h2c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_822 = 7'h2c == index | valid_0_44; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7775 = 7'h2d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_823 = 7'h2d == index | valid_0_45; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7776 = 7'h2e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_824 = 7'h2e == index | valid_0_46; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7777 = 7'h2f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_825 = 7'h2f == index | valid_0_47; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7778 = 7'h30 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_826 = 7'h30 == index | valid_0_48; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7779 = 7'h31 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_827 = 7'h31 == index | valid_0_49; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7780 = 7'h32 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_828 = 7'h32 == index | valid_0_50; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7781 = 7'h33 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_829 = 7'h33 == index | valid_0_51; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7782 = 7'h34 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_830 = 7'h34 == index | valid_0_52; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7783 = 7'h35 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_831 = 7'h35 == index | valid_0_53; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7784 = 7'h36 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_832 = 7'h36 == index | valid_0_54; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7785 = 7'h37 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_833 = 7'h37 == index | valid_0_55; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7786 = 7'h38 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_834 = 7'h38 == index | valid_0_56; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7787 = 7'h39 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_835 = 7'h39 == index | valid_0_57; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7788 = 7'h3a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_836 = 7'h3a == index | valid_0_58; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7789 = 7'h3b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_837 = 7'h3b == index | valid_0_59; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7790 = 7'h3c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_838 = 7'h3c == index | valid_0_60; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7791 = 7'h3d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_839 = 7'h3d == index | valid_0_61; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7792 = 7'h3e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_840 = 7'h3e == index | valid_0_62; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7793 = 7'h3f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_841 = 7'h3f == index | valid_0_63; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7794 = 7'h40 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_842 = 7'h40 == index | valid_0_64; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7795 = 7'h41 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_843 = 7'h41 == index | valid_0_65; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7796 = 7'h42 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_844 = 7'h42 == index | valid_0_66; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7797 = 7'h43 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_845 = 7'h43 == index | valid_0_67; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7798 = 7'h44 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_846 = 7'h44 == index | valid_0_68; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7799 = 7'h45 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_847 = 7'h45 == index | valid_0_69; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7800 = 7'h46 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_848 = 7'h46 == index | valid_0_70; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7801 = 7'h47 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_849 = 7'h47 == index | valid_0_71; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7802 = 7'h48 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_850 = 7'h48 == index | valid_0_72; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7803 = 7'h49 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_851 = 7'h49 == index | valid_0_73; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7804 = 7'h4a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_852 = 7'h4a == index | valid_0_74; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7805 = 7'h4b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_853 = 7'h4b == index | valid_0_75; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7806 = 7'h4c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_854 = 7'h4c == index | valid_0_76; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7807 = 7'h4d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_855 = 7'h4d == index | valid_0_77; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7808 = 7'h4e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_856 = 7'h4e == index | valid_0_78; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7809 = 7'h4f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_857 = 7'h4f == index | valid_0_79; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7810 = 7'h50 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_858 = 7'h50 == index | valid_0_80; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7811 = 7'h51 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_859 = 7'h51 == index | valid_0_81; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7812 = 7'h52 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_860 = 7'h52 == index | valid_0_82; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7813 = 7'h53 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_861 = 7'h53 == index | valid_0_83; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7814 = 7'h54 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_862 = 7'h54 == index | valid_0_84; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7815 = 7'h55 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_863 = 7'h55 == index | valid_0_85; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7816 = 7'h56 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_864 = 7'h56 == index | valid_0_86; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7817 = 7'h57 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_865 = 7'h57 == index | valid_0_87; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7818 = 7'h58 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_866 = 7'h58 == index | valid_0_88; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7819 = 7'h59 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_867 = 7'h59 == index | valid_0_89; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7820 = 7'h5a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_868 = 7'h5a == index | valid_0_90; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7821 = 7'h5b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_869 = 7'h5b == index | valid_0_91; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7822 = 7'h5c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_870 = 7'h5c == index | valid_0_92; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7823 = 7'h5d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_871 = 7'h5d == index | valid_0_93; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7824 = 7'h5e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_872 = 7'h5e == index | valid_0_94; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7825 = 7'h5f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_873 = 7'h5f == index | valid_0_95; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7826 = 7'h60 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_874 = 7'h60 == index | valid_0_96; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7827 = 7'h61 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_875 = 7'h61 == index | valid_0_97; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7828 = 7'h62 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_876 = 7'h62 == index | valid_0_98; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7829 = 7'h63 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_877 = 7'h63 == index | valid_0_99; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7830 = 7'h64 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_878 = 7'h64 == index | valid_0_100; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7831 = 7'h65 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_879 = 7'h65 == index | valid_0_101; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7832 = 7'h66 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_880 = 7'h66 == index | valid_0_102; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7833 = 7'h67 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_881 = 7'h67 == index | valid_0_103; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7834 = 7'h68 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_882 = 7'h68 == index | valid_0_104; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7835 = 7'h69 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_883 = 7'h69 == index | valid_0_105; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7836 = 7'h6a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_884 = 7'h6a == index | valid_0_106; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7837 = 7'h6b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_885 = 7'h6b == index | valid_0_107; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7838 = 7'h6c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_886 = 7'h6c == index | valid_0_108; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7839 = 7'h6d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_887 = 7'h6d == index | valid_0_109; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7840 = 7'h6e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_888 = 7'h6e == index | valid_0_110; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7841 = 7'h6f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_889 = 7'h6f == index | valid_0_111; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7842 = 7'h70 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_890 = 7'h70 == index | valid_0_112; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7843 = 7'h71 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_891 = 7'h71 == index | valid_0_113; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7844 = 7'h72 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_892 = 7'h72 == index | valid_0_114; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7845 = 7'h73 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_893 = 7'h73 == index | valid_0_115; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7846 = 7'h74 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_894 = 7'h74 == index | valid_0_116; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7847 = 7'h75 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_895 = 7'h75 == index | valid_0_117; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7848 = 7'h76 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_896 = 7'h76 == index | valid_0_118; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7849 = 7'h77 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_897 = 7'h77 == index | valid_0_119; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7850 = 7'h78 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_898 = 7'h78 == index | valid_0_120; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7851 = 7'h79 == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_899 = 7'h79 == index | valid_0_121; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7852 = 7'h7a == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_900 = 7'h7a == index | valid_0_122; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7853 = 7'h7b == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_901 = 7'h7b == index | valid_0_123; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7854 = 7'h7c == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_902 = 7'h7c == index | valid_0_124; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7855 = 7'h7d == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_903 = 7'h7d == index | valid_0_125; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7856 = 7'h7e == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_904 = 7'h7e == index | valid_0_126; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_7857 = 7'h7f == index; // @[i_cache.scala 21:26 89:{32,32}]
  wire  _GEN_905 = 7'h7f == index | valid_0_127; // @[i_cache.scala 21:26 89:{32,32}]
  wire [63:0] _GEN_906 = 7'h0 == index ? receive_data : ram_1_0; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_907 = 7'h1 == index ? receive_data : ram_1_1; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_908 = 7'h2 == index ? receive_data : ram_1_2; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_909 = 7'h3 == index ? receive_data : ram_1_3; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_910 = 7'h4 == index ? receive_data : ram_1_4; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_911 = 7'h5 == index ? receive_data : ram_1_5; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_912 = 7'h6 == index ? receive_data : ram_1_6; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_913 = 7'h7 == index ? receive_data : ram_1_7; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_914 = 7'h8 == index ? receive_data : ram_1_8; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_915 = 7'h9 == index ? receive_data : ram_1_9; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_916 = 7'ha == index ? receive_data : ram_1_10; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_917 = 7'hb == index ? receive_data : ram_1_11; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_918 = 7'hc == index ? receive_data : ram_1_12; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_919 = 7'hd == index ? receive_data : ram_1_13; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_920 = 7'he == index ? receive_data : ram_1_14; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_921 = 7'hf == index ? receive_data : ram_1_15; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_922 = 7'h10 == index ? receive_data : ram_1_16; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_923 = 7'h11 == index ? receive_data : ram_1_17; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_924 = 7'h12 == index ? receive_data : ram_1_18; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_925 = 7'h13 == index ? receive_data : ram_1_19; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_926 = 7'h14 == index ? receive_data : ram_1_20; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_927 = 7'h15 == index ? receive_data : ram_1_21; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_928 = 7'h16 == index ? receive_data : ram_1_22; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_929 = 7'h17 == index ? receive_data : ram_1_23; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_930 = 7'h18 == index ? receive_data : ram_1_24; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_931 = 7'h19 == index ? receive_data : ram_1_25; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_932 = 7'h1a == index ? receive_data : ram_1_26; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_933 = 7'h1b == index ? receive_data : ram_1_27; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_934 = 7'h1c == index ? receive_data : ram_1_28; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_935 = 7'h1d == index ? receive_data : ram_1_29; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_936 = 7'h1e == index ? receive_data : ram_1_30; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_937 = 7'h1f == index ? receive_data : ram_1_31; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_938 = 7'h20 == index ? receive_data : ram_1_32; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_939 = 7'h21 == index ? receive_data : ram_1_33; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_940 = 7'h22 == index ? receive_data : ram_1_34; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_941 = 7'h23 == index ? receive_data : ram_1_35; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_942 = 7'h24 == index ? receive_data : ram_1_36; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_943 = 7'h25 == index ? receive_data : ram_1_37; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_944 = 7'h26 == index ? receive_data : ram_1_38; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_945 = 7'h27 == index ? receive_data : ram_1_39; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_946 = 7'h28 == index ? receive_data : ram_1_40; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_947 = 7'h29 == index ? receive_data : ram_1_41; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_948 = 7'h2a == index ? receive_data : ram_1_42; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_949 = 7'h2b == index ? receive_data : ram_1_43; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_950 = 7'h2c == index ? receive_data : ram_1_44; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_951 = 7'h2d == index ? receive_data : ram_1_45; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_952 = 7'h2e == index ? receive_data : ram_1_46; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_953 = 7'h2f == index ? receive_data : ram_1_47; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_954 = 7'h30 == index ? receive_data : ram_1_48; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_955 = 7'h31 == index ? receive_data : ram_1_49; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_956 = 7'h32 == index ? receive_data : ram_1_50; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_957 = 7'h33 == index ? receive_data : ram_1_51; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_958 = 7'h34 == index ? receive_data : ram_1_52; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_959 = 7'h35 == index ? receive_data : ram_1_53; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_960 = 7'h36 == index ? receive_data : ram_1_54; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_961 = 7'h37 == index ? receive_data : ram_1_55; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_962 = 7'h38 == index ? receive_data : ram_1_56; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_963 = 7'h39 == index ? receive_data : ram_1_57; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_964 = 7'h3a == index ? receive_data : ram_1_58; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_965 = 7'h3b == index ? receive_data : ram_1_59; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_966 = 7'h3c == index ? receive_data : ram_1_60; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_967 = 7'h3d == index ? receive_data : ram_1_61; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_968 = 7'h3e == index ? receive_data : ram_1_62; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_969 = 7'h3f == index ? receive_data : ram_1_63; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_970 = 7'h40 == index ? receive_data : ram_1_64; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_971 = 7'h41 == index ? receive_data : ram_1_65; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_972 = 7'h42 == index ? receive_data : ram_1_66; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_973 = 7'h43 == index ? receive_data : ram_1_67; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_974 = 7'h44 == index ? receive_data : ram_1_68; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_975 = 7'h45 == index ? receive_data : ram_1_69; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_976 = 7'h46 == index ? receive_data : ram_1_70; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_977 = 7'h47 == index ? receive_data : ram_1_71; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_978 = 7'h48 == index ? receive_data : ram_1_72; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_979 = 7'h49 == index ? receive_data : ram_1_73; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_980 = 7'h4a == index ? receive_data : ram_1_74; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_981 = 7'h4b == index ? receive_data : ram_1_75; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_982 = 7'h4c == index ? receive_data : ram_1_76; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_983 = 7'h4d == index ? receive_data : ram_1_77; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_984 = 7'h4e == index ? receive_data : ram_1_78; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_985 = 7'h4f == index ? receive_data : ram_1_79; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_986 = 7'h50 == index ? receive_data : ram_1_80; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_987 = 7'h51 == index ? receive_data : ram_1_81; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_988 = 7'h52 == index ? receive_data : ram_1_82; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_989 = 7'h53 == index ? receive_data : ram_1_83; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_990 = 7'h54 == index ? receive_data : ram_1_84; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_991 = 7'h55 == index ? receive_data : ram_1_85; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_992 = 7'h56 == index ? receive_data : ram_1_86; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_993 = 7'h57 == index ? receive_data : ram_1_87; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_994 = 7'h58 == index ? receive_data : ram_1_88; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_995 = 7'h59 == index ? receive_data : ram_1_89; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_996 = 7'h5a == index ? receive_data : ram_1_90; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_997 = 7'h5b == index ? receive_data : ram_1_91; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_998 = 7'h5c == index ? receive_data : ram_1_92; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_999 = 7'h5d == index ? receive_data : ram_1_93; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1000 = 7'h5e == index ? receive_data : ram_1_94; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1001 = 7'h5f == index ? receive_data : ram_1_95; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1002 = 7'h60 == index ? receive_data : ram_1_96; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1003 = 7'h61 == index ? receive_data : ram_1_97; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1004 = 7'h62 == index ? receive_data : ram_1_98; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1005 = 7'h63 == index ? receive_data : ram_1_99; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1006 = 7'h64 == index ? receive_data : ram_1_100; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1007 = 7'h65 == index ? receive_data : ram_1_101; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1008 = 7'h66 == index ? receive_data : ram_1_102; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1009 = 7'h67 == index ? receive_data : ram_1_103; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1010 = 7'h68 == index ? receive_data : ram_1_104; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1011 = 7'h69 == index ? receive_data : ram_1_105; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1012 = 7'h6a == index ? receive_data : ram_1_106; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1013 = 7'h6b == index ? receive_data : ram_1_107; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1014 = 7'h6c == index ? receive_data : ram_1_108; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1015 = 7'h6d == index ? receive_data : ram_1_109; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1016 = 7'h6e == index ? receive_data : ram_1_110; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1017 = 7'h6f == index ? receive_data : ram_1_111; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1018 = 7'h70 == index ? receive_data : ram_1_112; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1019 = 7'h71 == index ? receive_data : ram_1_113; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1020 = 7'h72 == index ? receive_data : ram_1_114; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1021 = 7'h73 == index ? receive_data : ram_1_115; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1022 = 7'h74 == index ? receive_data : ram_1_116; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1023 = 7'h75 == index ? receive_data : ram_1_117; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1024 = 7'h76 == index ? receive_data : ram_1_118; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1025 = 7'h77 == index ? receive_data : ram_1_119; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1026 = 7'h78 == index ? receive_data : ram_1_120; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1027 = 7'h79 == index ? receive_data : ram_1_121; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1028 = 7'h7a == index ? receive_data : ram_1_122; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1029 = 7'h7b == index ? receive_data : ram_1_123; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1030 = 7'h7c == index ? receive_data : ram_1_124; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1031 = 7'h7d == index ? receive_data : ram_1_125; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1032 = 7'h7e == index ? receive_data : ram_1_126; // @[i_cache.scala 18:24 92:{30,30}]
  wire [63:0] _GEN_1033 = 7'h7f == index ? receive_data : ram_1_127; // @[i_cache.scala 18:24 92:{30,30}]
  wire [31:0] _GEN_1034 = 7'h0 == index ? _GEN_7706 : tag_1_0; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1035 = 7'h1 == index ? _GEN_7706 : tag_1_1; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1036 = 7'h2 == index ? _GEN_7706 : tag_1_2; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1037 = 7'h3 == index ? _GEN_7706 : tag_1_3; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1038 = 7'h4 == index ? _GEN_7706 : tag_1_4; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1039 = 7'h5 == index ? _GEN_7706 : tag_1_5; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1040 = 7'h6 == index ? _GEN_7706 : tag_1_6; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1041 = 7'h7 == index ? _GEN_7706 : tag_1_7; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1042 = 7'h8 == index ? _GEN_7706 : tag_1_8; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1043 = 7'h9 == index ? _GEN_7706 : tag_1_9; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1044 = 7'ha == index ? _GEN_7706 : tag_1_10; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1045 = 7'hb == index ? _GEN_7706 : tag_1_11; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1046 = 7'hc == index ? _GEN_7706 : tag_1_12; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1047 = 7'hd == index ? _GEN_7706 : tag_1_13; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1048 = 7'he == index ? _GEN_7706 : tag_1_14; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1049 = 7'hf == index ? _GEN_7706 : tag_1_15; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1050 = 7'h10 == index ? _GEN_7706 : tag_1_16; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1051 = 7'h11 == index ? _GEN_7706 : tag_1_17; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1052 = 7'h12 == index ? _GEN_7706 : tag_1_18; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1053 = 7'h13 == index ? _GEN_7706 : tag_1_19; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1054 = 7'h14 == index ? _GEN_7706 : tag_1_20; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1055 = 7'h15 == index ? _GEN_7706 : tag_1_21; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1056 = 7'h16 == index ? _GEN_7706 : tag_1_22; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1057 = 7'h17 == index ? _GEN_7706 : tag_1_23; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1058 = 7'h18 == index ? _GEN_7706 : tag_1_24; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1059 = 7'h19 == index ? _GEN_7706 : tag_1_25; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1060 = 7'h1a == index ? _GEN_7706 : tag_1_26; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1061 = 7'h1b == index ? _GEN_7706 : tag_1_27; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1062 = 7'h1c == index ? _GEN_7706 : tag_1_28; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1063 = 7'h1d == index ? _GEN_7706 : tag_1_29; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1064 = 7'h1e == index ? _GEN_7706 : tag_1_30; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1065 = 7'h1f == index ? _GEN_7706 : tag_1_31; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1066 = 7'h20 == index ? _GEN_7706 : tag_1_32; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1067 = 7'h21 == index ? _GEN_7706 : tag_1_33; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1068 = 7'h22 == index ? _GEN_7706 : tag_1_34; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1069 = 7'h23 == index ? _GEN_7706 : tag_1_35; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1070 = 7'h24 == index ? _GEN_7706 : tag_1_36; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1071 = 7'h25 == index ? _GEN_7706 : tag_1_37; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1072 = 7'h26 == index ? _GEN_7706 : tag_1_38; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1073 = 7'h27 == index ? _GEN_7706 : tag_1_39; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1074 = 7'h28 == index ? _GEN_7706 : tag_1_40; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1075 = 7'h29 == index ? _GEN_7706 : tag_1_41; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1076 = 7'h2a == index ? _GEN_7706 : tag_1_42; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1077 = 7'h2b == index ? _GEN_7706 : tag_1_43; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1078 = 7'h2c == index ? _GEN_7706 : tag_1_44; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1079 = 7'h2d == index ? _GEN_7706 : tag_1_45; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1080 = 7'h2e == index ? _GEN_7706 : tag_1_46; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1081 = 7'h2f == index ? _GEN_7706 : tag_1_47; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1082 = 7'h30 == index ? _GEN_7706 : tag_1_48; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1083 = 7'h31 == index ? _GEN_7706 : tag_1_49; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1084 = 7'h32 == index ? _GEN_7706 : tag_1_50; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1085 = 7'h33 == index ? _GEN_7706 : tag_1_51; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1086 = 7'h34 == index ? _GEN_7706 : tag_1_52; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1087 = 7'h35 == index ? _GEN_7706 : tag_1_53; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1088 = 7'h36 == index ? _GEN_7706 : tag_1_54; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1089 = 7'h37 == index ? _GEN_7706 : tag_1_55; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1090 = 7'h38 == index ? _GEN_7706 : tag_1_56; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1091 = 7'h39 == index ? _GEN_7706 : tag_1_57; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1092 = 7'h3a == index ? _GEN_7706 : tag_1_58; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1093 = 7'h3b == index ? _GEN_7706 : tag_1_59; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1094 = 7'h3c == index ? _GEN_7706 : tag_1_60; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1095 = 7'h3d == index ? _GEN_7706 : tag_1_61; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1096 = 7'h3e == index ? _GEN_7706 : tag_1_62; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1097 = 7'h3f == index ? _GEN_7706 : tag_1_63; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1098 = 7'h40 == index ? _GEN_7706 : tag_1_64; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1099 = 7'h41 == index ? _GEN_7706 : tag_1_65; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1100 = 7'h42 == index ? _GEN_7706 : tag_1_66; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1101 = 7'h43 == index ? _GEN_7706 : tag_1_67; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1102 = 7'h44 == index ? _GEN_7706 : tag_1_68; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1103 = 7'h45 == index ? _GEN_7706 : tag_1_69; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1104 = 7'h46 == index ? _GEN_7706 : tag_1_70; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1105 = 7'h47 == index ? _GEN_7706 : tag_1_71; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1106 = 7'h48 == index ? _GEN_7706 : tag_1_72; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1107 = 7'h49 == index ? _GEN_7706 : tag_1_73; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1108 = 7'h4a == index ? _GEN_7706 : tag_1_74; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1109 = 7'h4b == index ? _GEN_7706 : tag_1_75; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1110 = 7'h4c == index ? _GEN_7706 : tag_1_76; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1111 = 7'h4d == index ? _GEN_7706 : tag_1_77; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1112 = 7'h4e == index ? _GEN_7706 : tag_1_78; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1113 = 7'h4f == index ? _GEN_7706 : tag_1_79; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1114 = 7'h50 == index ? _GEN_7706 : tag_1_80; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1115 = 7'h51 == index ? _GEN_7706 : tag_1_81; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1116 = 7'h52 == index ? _GEN_7706 : tag_1_82; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1117 = 7'h53 == index ? _GEN_7706 : tag_1_83; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1118 = 7'h54 == index ? _GEN_7706 : tag_1_84; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1119 = 7'h55 == index ? _GEN_7706 : tag_1_85; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1120 = 7'h56 == index ? _GEN_7706 : tag_1_86; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1121 = 7'h57 == index ? _GEN_7706 : tag_1_87; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1122 = 7'h58 == index ? _GEN_7706 : tag_1_88; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1123 = 7'h59 == index ? _GEN_7706 : tag_1_89; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1124 = 7'h5a == index ? _GEN_7706 : tag_1_90; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1125 = 7'h5b == index ? _GEN_7706 : tag_1_91; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1126 = 7'h5c == index ? _GEN_7706 : tag_1_92; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1127 = 7'h5d == index ? _GEN_7706 : tag_1_93; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1128 = 7'h5e == index ? _GEN_7706 : tag_1_94; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1129 = 7'h5f == index ? _GEN_7706 : tag_1_95; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1130 = 7'h60 == index ? _GEN_7706 : tag_1_96; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1131 = 7'h61 == index ? _GEN_7706 : tag_1_97; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1132 = 7'h62 == index ? _GEN_7706 : tag_1_98; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1133 = 7'h63 == index ? _GEN_7706 : tag_1_99; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1134 = 7'h64 == index ? _GEN_7706 : tag_1_100; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1135 = 7'h65 == index ? _GEN_7706 : tag_1_101; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1136 = 7'h66 == index ? _GEN_7706 : tag_1_102; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1137 = 7'h67 == index ? _GEN_7706 : tag_1_103; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1138 = 7'h68 == index ? _GEN_7706 : tag_1_104; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1139 = 7'h69 == index ? _GEN_7706 : tag_1_105; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1140 = 7'h6a == index ? _GEN_7706 : tag_1_106; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1141 = 7'h6b == index ? _GEN_7706 : tag_1_107; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1142 = 7'h6c == index ? _GEN_7706 : tag_1_108; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1143 = 7'h6d == index ? _GEN_7706 : tag_1_109; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1144 = 7'h6e == index ? _GEN_7706 : tag_1_110; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1145 = 7'h6f == index ? _GEN_7706 : tag_1_111; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1146 = 7'h70 == index ? _GEN_7706 : tag_1_112; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1147 = 7'h71 == index ? _GEN_7706 : tag_1_113; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1148 = 7'h72 == index ? _GEN_7706 : tag_1_114; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1149 = 7'h73 == index ? _GEN_7706 : tag_1_115; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1150 = 7'h74 == index ? _GEN_7706 : tag_1_116; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1151 = 7'h75 == index ? _GEN_7706 : tag_1_117; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1152 = 7'h76 == index ? _GEN_7706 : tag_1_118; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1153 = 7'h77 == index ? _GEN_7706 : tag_1_119; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1154 = 7'h78 == index ? _GEN_7706 : tag_1_120; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1155 = 7'h79 == index ? _GEN_7706 : tag_1_121; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1156 = 7'h7a == index ? _GEN_7706 : tag_1_122; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1157 = 7'h7b == index ? _GEN_7706 : tag_1_123; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1158 = 7'h7c == index ? _GEN_7706 : tag_1_124; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1159 = 7'h7d == index ? _GEN_7706 : tag_1_125; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1160 = 7'h7e == index ? _GEN_7706 : tag_1_126; // @[i_cache.scala 20:24 93:{30,30}]
  wire [31:0] _GEN_1161 = 7'h7f == index ? _GEN_7706 : tag_1_127; // @[i_cache.scala 20:24 93:{30,30}]
  wire  _GEN_1162 = _GEN_7710 | valid_1_0; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1163 = _GEN_7712 | valid_1_1; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1164 = _GEN_7714 | valid_1_2; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1165 = _GEN_7718 | valid_1_3; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1166 = _GEN_7727 | valid_1_4; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1167 = _GEN_7729 | valid_1_5; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1168 = _GEN_7731 | valid_1_6; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1169 = _GEN_7733 | valid_1_7; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1170 = _GEN_7738 | valid_1_8; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1171 = _GEN_7739 | valid_1_9; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1172 = _GEN_7740 | valid_1_10; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1173 = _GEN_7741 | valid_1_11; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1174 = _GEN_7742 | valid_1_12; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1175 = _GEN_7743 | valid_1_13; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1176 = _GEN_7744 | valid_1_14; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1177 = _GEN_7745 | valid_1_15; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1178 = _GEN_7746 | valid_1_16; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1179 = _GEN_7747 | valid_1_17; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1180 = _GEN_7748 | valid_1_18; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1181 = _GEN_7749 | valid_1_19; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1182 = _GEN_7750 | valid_1_20; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1183 = _GEN_7751 | valid_1_21; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1184 = _GEN_7752 | valid_1_22; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1185 = _GEN_7753 | valid_1_23; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1186 = _GEN_7754 | valid_1_24; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1187 = _GEN_7755 | valid_1_25; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1188 = _GEN_7756 | valid_1_26; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1189 = _GEN_7757 | valid_1_27; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1190 = _GEN_7758 | valid_1_28; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1191 = _GEN_7759 | valid_1_29; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1192 = _GEN_7760 | valid_1_30; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1193 = _GEN_7761 | valid_1_31; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1194 = _GEN_7762 | valid_1_32; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1195 = _GEN_7763 | valid_1_33; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1196 = _GEN_7764 | valid_1_34; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1197 = _GEN_7765 | valid_1_35; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1198 = _GEN_7766 | valid_1_36; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1199 = _GEN_7767 | valid_1_37; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1200 = _GEN_7768 | valid_1_38; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1201 = _GEN_7769 | valid_1_39; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1202 = _GEN_7770 | valid_1_40; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1203 = _GEN_7771 | valid_1_41; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1204 = _GEN_7772 | valid_1_42; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1205 = _GEN_7773 | valid_1_43; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1206 = _GEN_7774 | valid_1_44; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1207 = _GEN_7775 | valid_1_45; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1208 = _GEN_7776 | valid_1_46; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1209 = _GEN_7777 | valid_1_47; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1210 = _GEN_7778 | valid_1_48; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1211 = _GEN_7779 | valid_1_49; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1212 = _GEN_7780 | valid_1_50; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1213 = _GEN_7781 | valid_1_51; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1214 = _GEN_7782 | valid_1_52; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1215 = _GEN_7783 | valid_1_53; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1216 = _GEN_7784 | valid_1_54; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1217 = _GEN_7785 | valid_1_55; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1218 = _GEN_7786 | valid_1_56; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1219 = _GEN_7787 | valid_1_57; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1220 = _GEN_7788 | valid_1_58; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1221 = _GEN_7789 | valid_1_59; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1222 = _GEN_7790 | valid_1_60; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1223 = _GEN_7791 | valid_1_61; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1224 = _GEN_7792 | valid_1_62; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1225 = _GEN_7793 | valid_1_63; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1226 = _GEN_7794 | valid_1_64; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1227 = _GEN_7795 | valid_1_65; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1228 = _GEN_7796 | valid_1_66; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1229 = _GEN_7797 | valid_1_67; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1230 = _GEN_7798 | valid_1_68; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1231 = _GEN_7799 | valid_1_69; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1232 = _GEN_7800 | valid_1_70; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1233 = _GEN_7801 | valid_1_71; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1234 = _GEN_7802 | valid_1_72; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1235 = _GEN_7803 | valid_1_73; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1236 = _GEN_7804 | valid_1_74; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1237 = _GEN_7805 | valid_1_75; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1238 = _GEN_7806 | valid_1_76; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1239 = _GEN_7807 | valid_1_77; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1240 = _GEN_7808 | valid_1_78; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1241 = _GEN_7809 | valid_1_79; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1242 = _GEN_7810 | valid_1_80; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1243 = _GEN_7811 | valid_1_81; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1244 = _GEN_7812 | valid_1_82; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1245 = _GEN_7813 | valid_1_83; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1246 = _GEN_7814 | valid_1_84; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1247 = _GEN_7815 | valid_1_85; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1248 = _GEN_7816 | valid_1_86; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1249 = _GEN_7817 | valid_1_87; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1250 = _GEN_7818 | valid_1_88; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1251 = _GEN_7819 | valid_1_89; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1252 = _GEN_7820 | valid_1_90; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1253 = _GEN_7821 | valid_1_91; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1254 = _GEN_7822 | valid_1_92; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1255 = _GEN_7823 | valid_1_93; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1256 = _GEN_7824 | valid_1_94; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1257 = _GEN_7825 | valid_1_95; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1258 = _GEN_7826 | valid_1_96; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1259 = _GEN_7827 | valid_1_97; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1260 = _GEN_7828 | valid_1_98; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1261 = _GEN_7829 | valid_1_99; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1262 = _GEN_7830 | valid_1_100; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1263 = _GEN_7831 | valid_1_101; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1264 = _GEN_7832 | valid_1_102; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1265 = _GEN_7833 | valid_1_103; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1266 = _GEN_7834 | valid_1_104; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1267 = _GEN_7835 | valid_1_105; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1268 = _GEN_7836 | valid_1_106; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1269 = _GEN_7837 | valid_1_107; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1270 = _GEN_7838 | valid_1_108; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1271 = _GEN_7839 | valid_1_109; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1272 = _GEN_7840 | valid_1_110; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1273 = _GEN_7841 | valid_1_111; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1274 = _GEN_7842 | valid_1_112; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1275 = _GEN_7843 | valid_1_113; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1276 = _GEN_7844 | valid_1_114; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1277 = _GEN_7845 | valid_1_115; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1278 = _GEN_7846 | valid_1_116; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1279 = _GEN_7847 | valid_1_117; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1280 = _GEN_7848 | valid_1_118; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1281 = _GEN_7849 | valid_1_119; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1282 = _GEN_7850 | valid_1_120; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1283 = _GEN_7851 | valid_1_121; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1284 = _GEN_7852 | valid_1_122; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1285 = _GEN_7853 | valid_1_123; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1286 = _GEN_7854 | valid_1_124; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1287 = _GEN_7855 | valid_1_125; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1288 = _GEN_7856 | valid_1_126; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _GEN_1289 = _GEN_7857 | valid_1_127; // @[i_cache.scala 22:26 94:{32,32}]
  wire  _T_14 = ~quene; // @[i_cache.scala 97:27]
  wire [63:0] _GEN_2058 = ~quene ? _GEN_522 : ram_0_0; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2059 = ~quene ? _GEN_523 : ram_0_1; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2060 = ~quene ? _GEN_524 : ram_0_2; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2061 = ~quene ? _GEN_525 : ram_0_3; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2062 = ~quene ? _GEN_526 : ram_0_4; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2063 = ~quene ? _GEN_527 : ram_0_5; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2064 = ~quene ? _GEN_528 : ram_0_6; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2065 = ~quene ? _GEN_529 : ram_0_7; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2066 = ~quene ? _GEN_530 : ram_0_8; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2067 = ~quene ? _GEN_531 : ram_0_9; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2068 = ~quene ? _GEN_532 : ram_0_10; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2069 = ~quene ? _GEN_533 : ram_0_11; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2070 = ~quene ? _GEN_534 : ram_0_12; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2071 = ~quene ? _GEN_535 : ram_0_13; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2072 = ~quene ? _GEN_536 : ram_0_14; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2073 = ~quene ? _GEN_537 : ram_0_15; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2074 = ~quene ? _GEN_538 : ram_0_16; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2075 = ~quene ? _GEN_539 : ram_0_17; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2076 = ~quene ? _GEN_540 : ram_0_18; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2077 = ~quene ? _GEN_541 : ram_0_19; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2078 = ~quene ? _GEN_542 : ram_0_20; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2079 = ~quene ? _GEN_543 : ram_0_21; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2080 = ~quene ? _GEN_544 : ram_0_22; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2081 = ~quene ? _GEN_545 : ram_0_23; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2082 = ~quene ? _GEN_546 : ram_0_24; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2083 = ~quene ? _GEN_547 : ram_0_25; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2084 = ~quene ? _GEN_548 : ram_0_26; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2085 = ~quene ? _GEN_549 : ram_0_27; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2086 = ~quene ? _GEN_550 : ram_0_28; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2087 = ~quene ? _GEN_551 : ram_0_29; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2088 = ~quene ? _GEN_552 : ram_0_30; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2089 = ~quene ? _GEN_553 : ram_0_31; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2090 = ~quene ? _GEN_554 : ram_0_32; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2091 = ~quene ? _GEN_555 : ram_0_33; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2092 = ~quene ? _GEN_556 : ram_0_34; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2093 = ~quene ? _GEN_557 : ram_0_35; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2094 = ~quene ? _GEN_558 : ram_0_36; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2095 = ~quene ? _GEN_559 : ram_0_37; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2096 = ~quene ? _GEN_560 : ram_0_38; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2097 = ~quene ? _GEN_561 : ram_0_39; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2098 = ~quene ? _GEN_562 : ram_0_40; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2099 = ~quene ? _GEN_563 : ram_0_41; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2100 = ~quene ? _GEN_564 : ram_0_42; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2101 = ~quene ? _GEN_565 : ram_0_43; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2102 = ~quene ? _GEN_566 : ram_0_44; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2103 = ~quene ? _GEN_567 : ram_0_45; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2104 = ~quene ? _GEN_568 : ram_0_46; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2105 = ~quene ? _GEN_569 : ram_0_47; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2106 = ~quene ? _GEN_570 : ram_0_48; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2107 = ~quene ? _GEN_571 : ram_0_49; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2108 = ~quene ? _GEN_572 : ram_0_50; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2109 = ~quene ? _GEN_573 : ram_0_51; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2110 = ~quene ? _GEN_574 : ram_0_52; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2111 = ~quene ? _GEN_575 : ram_0_53; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2112 = ~quene ? _GEN_576 : ram_0_54; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2113 = ~quene ? _GEN_577 : ram_0_55; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2114 = ~quene ? _GEN_578 : ram_0_56; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2115 = ~quene ? _GEN_579 : ram_0_57; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2116 = ~quene ? _GEN_580 : ram_0_58; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2117 = ~quene ? _GEN_581 : ram_0_59; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2118 = ~quene ? _GEN_582 : ram_0_60; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2119 = ~quene ? _GEN_583 : ram_0_61; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2120 = ~quene ? _GEN_584 : ram_0_62; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2121 = ~quene ? _GEN_585 : ram_0_63; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2122 = ~quene ? _GEN_586 : ram_0_64; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2123 = ~quene ? _GEN_587 : ram_0_65; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2124 = ~quene ? _GEN_588 : ram_0_66; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2125 = ~quene ? _GEN_589 : ram_0_67; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2126 = ~quene ? _GEN_590 : ram_0_68; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2127 = ~quene ? _GEN_591 : ram_0_69; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2128 = ~quene ? _GEN_592 : ram_0_70; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2129 = ~quene ? _GEN_593 : ram_0_71; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2130 = ~quene ? _GEN_594 : ram_0_72; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2131 = ~quene ? _GEN_595 : ram_0_73; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2132 = ~quene ? _GEN_596 : ram_0_74; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2133 = ~quene ? _GEN_597 : ram_0_75; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2134 = ~quene ? _GEN_598 : ram_0_76; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2135 = ~quene ? _GEN_599 : ram_0_77; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2136 = ~quene ? _GEN_600 : ram_0_78; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2137 = ~quene ? _GEN_601 : ram_0_79; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2138 = ~quene ? _GEN_602 : ram_0_80; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2139 = ~quene ? _GEN_603 : ram_0_81; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2140 = ~quene ? _GEN_604 : ram_0_82; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2141 = ~quene ? _GEN_605 : ram_0_83; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2142 = ~quene ? _GEN_606 : ram_0_84; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2143 = ~quene ? _GEN_607 : ram_0_85; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2144 = ~quene ? _GEN_608 : ram_0_86; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2145 = ~quene ? _GEN_609 : ram_0_87; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2146 = ~quene ? _GEN_610 : ram_0_88; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2147 = ~quene ? _GEN_611 : ram_0_89; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2148 = ~quene ? _GEN_612 : ram_0_90; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2149 = ~quene ? _GEN_613 : ram_0_91; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2150 = ~quene ? _GEN_614 : ram_0_92; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2151 = ~quene ? _GEN_615 : ram_0_93; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2152 = ~quene ? _GEN_616 : ram_0_94; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2153 = ~quene ? _GEN_617 : ram_0_95; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2154 = ~quene ? _GEN_618 : ram_0_96; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2155 = ~quene ? _GEN_619 : ram_0_97; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2156 = ~quene ? _GEN_620 : ram_0_98; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2157 = ~quene ? _GEN_621 : ram_0_99; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2158 = ~quene ? _GEN_622 : ram_0_100; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2159 = ~quene ? _GEN_623 : ram_0_101; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2160 = ~quene ? _GEN_624 : ram_0_102; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2161 = ~quene ? _GEN_625 : ram_0_103; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2162 = ~quene ? _GEN_626 : ram_0_104; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2163 = ~quene ? _GEN_627 : ram_0_105; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2164 = ~quene ? _GEN_628 : ram_0_106; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2165 = ~quene ? _GEN_629 : ram_0_107; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2166 = ~quene ? _GEN_630 : ram_0_108; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2167 = ~quene ? _GEN_631 : ram_0_109; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2168 = ~quene ? _GEN_632 : ram_0_110; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2169 = ~quene ? _GEN_633 : ram_0_111; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2170 = ~quene ? _GEN_634 : ram_0_112; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2171 = ~quene ? _GEN_635 : ram_0_113; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2172 = ~quene ? _GEN_636 : ram_0_114; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2173 = ~quene ? _GEN_637 : ram_0_115; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2174 = ~quene ? _GEN_638 : ram_0_116; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2175 = ~quene ? _GEN_639 : ram_0_117; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2176 = ~quene ? _GEN_640 : ram_0_118; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2177 = ~quene ? _GEN_641 : ram_0_119; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2178 = ~quene ? _GEN_642 : ram_0_120; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2179 = ~quene ? _GEN_643 : ram_0_121; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2180 = ~quene ? _GEN_644 : ram_0_122; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2181 = ~quene ? _GEN_645 : ram_0_123; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2182 = ~quene ? _GEN_646 : ram_0_124; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2183 = ~quene ? _GEN_647 : ram_0_125; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2184 = ~quene ? _GEN_648 : ram_0_126; // @[i_cache.scala 17:24 97:34]
  wire [63:0] _GEN_2185 = ~quene ? _GEN_649 : ram_0_127; // @[i_cache.scala 17:24 97:34]
  wire [31:0] _GEN_2186 = ~quene ? _GEN_650 : tag_0_0; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2187 = ~quene ? _GEN_651 : tag_0_1; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2188 = ~quene ? _GEN_652 : tag_0_2; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2189 = ~quene ? _GEN_653 : tag_0_3; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2190 = ~quene ? _GEN_654 : tag_0_4; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2191 = ~quene ? _GEN_655 : tag_0_5; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2192 = ~quene ? _GEN_656 : tag_0_6; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2193 = ~quene ? _GEN_657 : tag_0_7; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2194 = ~quene ? _GEN_658 : tag_0_8; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2195 = ~quene ? _GEN_659 : tag_0_9; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2196 = ~quene ? _GEN_660 : tag_0_10; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2197 = ~quene ? _GEN_661 : tag_0_11; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2198 = ~quene ? _GEN_662 : tag_0_12; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2199 = ~quene ? _GEN_663 : tag_0_13; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2200 = ~quene ? _GEN_664 : tag_0_14; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2201 = ~quene ? _GEN_665 : tag_0_15; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2202 = ~quene ? _GEN_666 : tag_0_16; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2203 = ~quene ? _GEN_667 : tag_0_17; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2204 = ~quene ? _GEN_668 : tag_0_18; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2205 = ~quene ? _GEN_669 : tag_0_19; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2206 = ~quene ? _GEN_670 : tag_0_20; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2207 = ~quene ? _GEN_671 : tag_0_21; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2208 = ~quene ? _GEN_672 : tag_0_22; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2209 = ~quene ? _GEN_673 : tag_0_23; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2210 = ~quene ? _GEN_674 : tag_0_24; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2211 = ~quene ? _GEN_675 : tag_0_25; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2212 = ~quene ? _GEN_676 : tag_0_26; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2213 = ~quene ? _GEN_677 : tag_0_27; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2214 = ~quene ? _GEN_678 : tag_0_28; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2215 = ~quene ? _GEN_679 : tag_0_29; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2216 = ~quene ? _GEN_680 : tag_0_30; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2217 = ~quene ? _GEN_681 : tag_0_31; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2218 = ~quene ? _GEN_682 : tag_0_32; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2219 = ~quene ? _GEN_683 : tag_0_33; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2220 = ~quene ? _GEN_684 : tag_0_34; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2221 = ~quene ? _GEN_685 : tag_0_35; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2222 = ~quene ? _GEN_686 : tag_0_36; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2223 = ~quene ? _GEN_687 : tag_0_37; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2224 = ~quene ? _GEN_688 : tag_0_38; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2225 = ~quene ? _GEN_689 : tag_0_39; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2226 = ~quene ? _GEN_690 : tag_0_40; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2227 = ~quene ? _GEN_691 : tag_0_41; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2228 = ~quene ? _GEN_692 : tag_0_42; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2229 = ~quene ? _GEN_693 : tag_0_43; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2230 = ~quene ? _GEN_694 : tag_0_44; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2231 = ~quene ? _GEN_695 : tag_0_45; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2232 = ~quene ? _GEN_696 : tag_0_46; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2233 = ~quene ? _GEN_697 : tag_0_47; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2234 = ~quene ? _GEN_698 : tag_0_48; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2235 = ~quene ? _GEN_699 : tag_0_49; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2236 = ~quene ? _GEN_700 : tag_0_50; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2237 = ~quene ? _GEN_701 : tag_0_51; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2238 = ~quene ? _GEN_702 : tag_0_52; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2239 = ~quene ? _GEN_703 : tag_0_53; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2240 = ~quene ? _GEN_704 : tag_0_54; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2241 = ~quene ? _GEN_705 : tag_0_55; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2242 = ~quene ? _GEN_706 : tag_0_56; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2243 = ~quene ? _GEN_707 : tag_0_57; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2244 = ~quene ? _GEN_708 : tag_0_58; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2245 = ~quene ? _GEN_709 : tag_0_59; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2246 = ~quene ? _GEN_710 : tag_0_60; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2247 = ~quene ? _GEN_711 : tag_0_61; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2248 = ~quene ? _GEN_712 : tag_0_62; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2249 = ~quene ? _GEN_713 : tag_0_63; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2250 = ~quene ? _GEN_714 : tag_0_64; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2251 = ~quene ? _GEN_715 : tag_0_65; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2252 = ~quene ? _GEN_716 : tag_0_66; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2253 = ~quene ? _GEN_717 : tag_0_67; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2254 = ~quene ? _GEN_718 : tag_0_68; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2255 = ~quene ? _GEN_719 : tag_0_69; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2256 = ~quene ? _GEN_720 : tag_0_70; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2257 = ~quene ? _GEN_721 : tag_0_71; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2258 = ~quene ? _GEN_722 : tag_0_72; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2259 = ~quene ? _GEN_723 : tag_0_73; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2260 = ~quene ? _GEN_724 : tag_0_74; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2261 = ~quene ? _GEN_725 : tag_0_75; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2262 = ~quene ? _GEN_726 : tag_0_76; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2263 = ~quene ? _GEN_727 : tag_0_77; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2264 = ~quene ? _GEN_728 : tag_0_78; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2265 = ~quene ? _GEN_729 : tag_0_79; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2266 = ~quene ? _GEN_730 : tag_0_80; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2267 = ~quene ? _GEN_731 : tag_0_81; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2268 = ~quene ? _GEN_732 : tag_0_82; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2269 = ~quene ? _GEN_733 : tag_0_83; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2270 = ~quene ? _GEN_734 : tag_0_84; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2271 = ~quene ? _GEN_735 : tag_0_85; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2272 = ~quene ? _GEN_736 : tag_0_86; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2273 = ~quene ? _GEN_737 : tag_0_87; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2274 = ~quene ? _GEN_738 : tag_0_88; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2275 = ~quene ? _GEN_739 : tag_0_89; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2276 = ~quene ? _GEN_740 : tag_0_90; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2277 = ~quene ? _GEN_741 : tag_0_91; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2278 = ~quene ? _GEN_742 : tag_0_92; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2279 = ~quene ? _GEN_743 : tag_0_93; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2280 = ~quene ? _GEN_744 : tag_0_94; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2281 = ~quene ? _GEN_745 : tag_0_95; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2282 = ~quene ? _GEN_746 : tag_0_96; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2283 = ~quene ? _GEN_747 : tag_0_97; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2284 = ~quene ? _GEN_748 : tag_0_98; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2285 = ~quene ? _GEN_749 : tag_0_99; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2286 = ~quene ? _GEN_750 : tag_0_100; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2287 = ~quene ? _GEN_751 : tag_0_101; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2288 = ~quene ? _GEN_752 : tag_0_102; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2289 = ~quene ? _GEN_753 : tag_0_103; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2290 = ~quene ? _GEN_754 : tag_0_104; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2291 = ~quene ? _GEN_755 : tag_0_105; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2292 = ~quene ? _GEN_756 : tag_0_106; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2293 = ~quene ? _GEN_757 : tag_0_107; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2294 = ~quene ? _GEN_758 : tag_0_108; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2295 = ~quene ? _GEN_759 : tag_0_109; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2296 = ~quene ? _GEN_760 : tag_0_110; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2297 = ~quene ? _GEN_761 : tag_0_111; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2298 = ~quene ? _GEN_762 : tag_0_112; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2299 = ~quene ? _GEN_763 : tag_0_113; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2300 = ~quene ? _GEN_764 : tag_0_114; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2301 = ~quene ? _GEN_765 : tag_0_115; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2302 = ~quene ? _GEN_766 : tag_0_116; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2303 = ~quene ? _GEN_767 : tag_0_117; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2304 = ~quene ? _GEN_768 : tag_0_118; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2305 = ~quene ? _GEN_769 : tag_0_119; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2306 = ~quene ? _GEN_770 : tag_0_120; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2307 = ~quene ? _GEN_771 : tag_0_121; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2308 = ~quene ? _GEN_772 : tag_0_122; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2309 = ~quene ? _GEN_773 : tag_0_123; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2310 = ~quene ? _GEN_774 : tag_0_124; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2311 = ~quene ? _GEN_775 : tag_0_125; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2312 = ~quene ? _GEN_776 : tag_0_126; // @[i_cache.scala 19:24 97:34]
  wire [31:0] _GEN_2313 = ~quene ? _GEN_777 : tag_0_127; // @[i_cache.scala 19:24 97:34]
  wire  _GEN_2314 = ~quene ? _GEN_778 : valid_0_0; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2315 = ~quene ? _GEN_779 : valid_0_1; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2316 = ~quene ? _GEN_780 : valid_0_2; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2317 = ~quene ? _GEN_781 : valid_0_3; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2318 = ~quene ? _GEN_782 : valid_0_4; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2319 = ~quene ? _GEN_783 : valid_0_5; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2320 = ~quene ? _GEN_784 : valid_0_6; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2321 = ~quene ? _GEN_785 : valid_0_7; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2322 = ~quene ? _GEN_786 : valid_0_8; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2323 = ~quene ? _GEN_787 : valid_0_9; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2324 = ~quene ? _GEN_788 : valid_0_10; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2325 = ~quene ? _GEN_789 : valid_0_11; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2326 = ~quene ? _GEN_790 : valid_0_12; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2327 = ~quene ? _GEN_791 : valid_0_13; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2328 = ~quene ? _GEN_792 : valid_0_14; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2329 = ~quene ? _GEN_793 : valid_0_15; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2330 = ~quene ? _GEN_794 : valid_0_16; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2331 = ~quene ? _GEN_795 : valid_0_17; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2332 = ~quene ? _GEN_796 : valid_0_18; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2333 = ~quene ? _GEN_797 : valid_0_19; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2334 = ~quene ? _GEN_798 : valid_0_20; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2335 = ~quene ? _GEN_799 : valid_0_21; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2336 = ~quene ? _GEN_800 : valid_0_22; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2337 = ~quene ? _GEN_801 : valid_0_23; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2338 = ~quene ? _GEN_802 : valid_0_24; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2339 = ~quene ? _GEN_803 : valid_0_25; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2340 = ~quene ? _GEN_804 : valid_0_26; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2341 = ~quene ? _GEN_805 : valid_0_27; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2342 = ~quene ? _GEN_806 : valid_0_28; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2343 = ~quene ? _GEN_807 : valid_0_29; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2344 = ~quene ? _GEN_808 : valid_0_30; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2345 = ~quene ? _GEN_809 : valid_0_31; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2346 = ~quene ? _GEN_810 : valid_0_32; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2347 = ~quene ? _GEN_811 : valid_0_33; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2348 = ~quene ? _GEN_812 : valid_0_34; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2349 = ~quene ? _GEN_813 : valid_0_35; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2350 = ~quene ? _GEN_814 : valid_0_36; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2351 = ~quene ? _GEN_815 : valid_0_37; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2352 = ~quene ? _GEN_816 : valid_0_38; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2353 = ~quene ? _GEN_817 : valid_0_39; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2354 = ~quene ? _GEN_818 : valid_0_40; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2355 = ~quene ? _GEN_819 : valid_0_41; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2356 = ~quene ? _GEN_820 : valid_0_42; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2357 = ~quene ? _GEN_821 : valid_0_43; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2358 = ~quene ? _GEN_822 : valid_0_44; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2359 = ~quene ? _GEN_823 : valid_0_45; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2360 = ~quene ? _GEN_824 : valid_0_46; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2361 = ~quene ? _GEN_825 : valid_0_47; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2362 = ~quene ? _GEN_826 : valid_0_48; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2363 = ~quene ? _GEN_827 : valid_0_49; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2364 = ~quene ? _GEN_828 : valid_0_50; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2365 = ~quene ? _GEN_829 : valid_0_51; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2366 = ~quene ? _GEN_830 : valid_0_52; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2367 = ~quene ? _GEN_831 : valid_0_53; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2368 = ~quene ? _GEN_832 : valid_0_54; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2369 = ~quene ? _GEN_833 : valid_0_55; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2370 = ~quene ? _GEN_834 : valid_0_56; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2371 = ~quene ? _GEN_835 : valid_0_57; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2372 = ~quene ? _GEN_836 : valid_0_58; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2373 = ~quene ? _GEN_837 : valid_0_59; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2374 = ~quene ? _GEN_838 : valid_0_60; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2375 = ~quene ? _GEN_839 : valid_0_61; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2376 = ~quene ? _GEN_840 : valid_0_62; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2377 = ~quene ? _GEN_841 : valid_0_63; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2378 = ~quene ? _GEN_842 : valid_0_64; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2379 = ~quene ? _GEN_843 : valid_0_65; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2380 = ~quene ? _GEN_844 : valid_0_66; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2381 = ~quene ? _GEN_845 : valid_0_67; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2382 = ~quene ? _GEN_846 : valid_0_68; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2383 = ~quene ? _GEN_847 : valid_0_69; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2384 = ~quene ? _GEN_848 : valid_0_70; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2385 = ~quene ? _GEN_849 : valid_0_71; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2386 = ~quene ? _GEN_850 : valid_0_72; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2387 = ~quene ? _GEN_851 : valid_0_73; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2388 = ~quene ? _GEN_852 : valid_0_74; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2389 = ~quene ? _GEN_853 : valid_0_75; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2390 = ~quene ? _GEN_854 : valid_0_76; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2391 = ~quene ? _GEN_855 : valid_0_77; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2392 = ~quene ? _GEN_856 : valid_0_78; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2393 = ~quene ? _GEN_857 : valid_0_79; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2394 = ~quene ? _GEN_858 : valid_0_80; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2395 = ~quene ? _GEN_859 : valid_0_81; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2396 = ~quene ? _GEN_860 : valid_0_82; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2397 = ~quene ? _GEN_861 : valid_0_83; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2398 = ~quene ? _GEN_862 : valid_0_84; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2399 = ~quene ? _GEN_863 : valid_0_85; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2400 = ~quene ? _GEN_864 : valid_0_86; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2401 = ~quene ? _GEN_865 : valid_0_87; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2402 = ~quene ? _GEN_866 : valid_0_88; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2403 = ~quene ? _GEN_867 : valid_0_89; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2404 = ~quene ? _GEN_868 : valid_0_90; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2405 = ~quene ? _GEN_869 : valid_0_91; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2406 = ~quene ? _GEN_870 : valid_0_92; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2407 = ~quene ? _GEN_871 : valid_0_93; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2408 = ~quene ? _GEN_872 : valid_0_94; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2409 = ~quene ? _GEN_873 : valid_0_95; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2410 = ~quene ? _GEN_874 : valid_0_96; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2411 = ~quene ? _GEN_875 : valid_0_97; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2412 = ~quene ? _GEN_876 : valid_0_98; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2413 = ~quene ? _GEN_877 : valid_0_99; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2414 = ~quene ? _GEN_878 : valid_0_100; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2415 = ~quene ? _GEN_879 : valid_0_101; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2416 = ~quene ? _GEN_880 : valid_0_102; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2417 = ~quene ? _GEN_881 : valid_0_103; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2418 = ~quene ? _GEN_882 : valid_0_104; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2419 = ~quene ? _GEN_883 : valid_0_105; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2420 = ~quene ? _GEN_884 : valid_0_106; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2421 = ~quene ? _GEN_885 : valid_0_107; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2422 = ~quene ? _GEN_886 : valid_0_108; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2423 = ~quene ? _GEN_887 : valid_0_109; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2424 = ~quene ? _GEN_888 : valid_0_110; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2425 = ~quene ? _GEN_889 : valid_0_111; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2426 = ~quene ? _GEN_890 : valid_0_112; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2427 = ~quene ? _GEN_891 : valid_0_113; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2428 = ~quene ? _GEN_892 : valid_0_114; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2429 = ~quene ? _GEN_893 : valid_0_115; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2430 = ~quene ? _GEN_894 : valid_0_116; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2431 = ~quene ? _GEN_895 : valid_0_117; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2432 = ~quene ? _GEN_896 : valid_0_118; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2433 = ~quene ? _GEN_897 : valid_0_119; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2434 = ~quene ? _GEN_898 : valid_0_120; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2435 = ~quene ? _GEN_899 : valid_0_121; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2436 = ~quene ? _GEN_900 : valid_0_122; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2437 = ~quene ? _GEN_901 : valid_0_123; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2438 = ~quene ? _GEN_902 : valid_0_124; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2439 = ~quene ? _GEN_903 : valid_0_125; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2440 = ~quene ? _GEN_904 : valid_0_126; // @[i_cache.scala 21:26 97:34]
  wire  _GEN_2441 = ~quene ? _GEN_905 : valid_0_127; // @[i_cache.scala 21:26 97:34]
  wire [63:0] _GEN_2443 = ~quene ? ram_1_0 : _GEN_906; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2444 = ~quene ? ram_1_1 : _GEN_907; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2445 = ~quene ? ram_1_2 : _GEN_908; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2446 = ~quene ? ram_1_3 : _GEN_909; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2447 = ~quene ? ram_1_4 : _GEN_910; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2448 = ~quene ? ram_1_5 : _GEN_911; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2449 = ~quene ? ram_1_6 : _GEN_912; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2450 = ~quene ? ram_1_7 : _GEN_913; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2451 = ~quene ? ram_1_8 : _GEN_914; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2452 = ~quene ? ram_1_9 : _GEN_915; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2453 = ~quene ? ram_1_10 : _GEN_916; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2454 = ~quene ? ram_1_11 : _GEN_917; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2455 = ~quene ? ram_1_12 : _GEN_918; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2456 = ~quene ? ram_1_13 : _GEN_919; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2457 = ~quene ? ram_1_14 : _GEN_920; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2458 = ~quene ? ram_1_15 : _GEN_921; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2459 = ~quene ? ram_1_16 : _GEN_922; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2460 = ~quene ? ram_1_17 : _GEN_923; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2461 = ~quene ? ram_1_18 : _GEN_924; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2462 = ~quene ? ram_1_19 : _GEN_925; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2463 = ~quene ? ram_1_20 : _GEN_926; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2464 = ~quene ? ram_1_21 : _GEN_927; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2465 = ~quene ? ram_1_22 : _GEN_928; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2466 = ~quene ? ram_1_23 : _GEN_929; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2467 = ~quene ? ram_1_24 : _GEN_930; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2468 = ~quene ? ram_1_25 : _GEN_931; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2469 = ~quene ? ram_1_26 : _GEN_932; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2470 = ~quene ? ram_1_27 : _GEN_933; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2471 = ~quene ? ram_1_28 : _GEN_934; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2472 = ~quene ? ram_1_29 : _GEN_935; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2473 = ~quene ? ram_1_30 : _GEN_936; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2474 = ~quene ? ram_1_31 : _GEN_937; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2475 = ~quene ? ram_1_32 : _GEN_938; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2476 = ~quene ? ram_1_33 : _GEN_939; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2477 = ~quene ? ram_1_34 : _GEN_940; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2478 = ~quene ? ram_1_35 : _GEN_941; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2479 = ~quene ? ram_1_36 : _GEN_942; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2480 = ~quene ? ram_1_37 : _GEN_943; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2481 = ~quene ? ram_1_38 : _GEN_944; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2482 = ~quene ? ram_1_39 : _GEN_945; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2483 = ~quene ? ram_1_40 : _GEN_946; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2484 = ~quene ? ram_1_41 : _GEN_947; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2485 = ~quene ? ram_1_42 : _GEN_948; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2486 = ~quene ? ram_1_43 : _GEN_949; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2487 = ~quene ? ram_1_44 : _GEN_950; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2488 = ~quene ? ram_1_45 : _GEN_951; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2489 = ~quene ? ram_1_46 : _GEN_952; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2490 = ~quene ? ram_1_47 : _GEN_953; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2491 = ~quene ? ram_1_48 : _GEN_954; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2492 = ~quene ? ram_1_49 : _GEN_955; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2493 = ~quene ? ram_1_50 : _GEN_956; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2494 = ~quene ? ram_1_51 : _GEN_957; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2495 = ~quene ? ram_1_52 : _GEN_958; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2496 = ~quene ? ram_1_53 : _GEN_959; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2497 = ~quene ? ram_1_54 : _GEN_960; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2498 = ~quene ? ram_1_55 : _GEN_961; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2499 = ~quene ? ram_1_56 : _GEN_962; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2500 = ~quene ? ram_1_57 : _GEN_963; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2501 = ~quene ? ram_1_58 : _GEN_964; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2502 = ~quene ? ram_1_59 : _GEN_965; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2503 = ~quene ? ram_1_60 : _GEN_966; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2504 = ~quene ? ram_1_61 : _GEN_967; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2505 = ~quene ? ram_1_62 : _GEN_968; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2506 = ~quene ? ram_1_63 : _GEN_969; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2507 = ~quene ? ram_1_64 : _GEN_970; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2508 = ~quene ? ram_1_65 : _GEN_971; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2509 = ~quene ? ram_1_66 : _GEN_972; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2510 = ~quene ? ram_1_67 : _GEN_973; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2511 = ~quene ? ram_1_68 : _GEN_974; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2512 = ~quene ? ram_1_69 : _GEN_975; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2513 = ~quene ? ram_1_70 : _GEN_976; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2514 = ~quene ? ram_1_71 : _GEN_977; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2515 = ~quene ? ram_1_72 : _GEN_978; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2516 = ~quene ? ram_1_73 : _GEN_979; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2517 = ~quene ? ram_1_74 : _GEN_980; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2518 = ~quene ? ram_1_75 : _GEN_981; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2519 = ~quene ? ram_1_76 : _GEN_982; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2520 = ~quene ? ram_1_77 : _GEN_983; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2521 = ~quene ? ram_1_78 : _GEN_984; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2522 = ~quene ? ram_1_79 : _GEN_985; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2523 = ~quene ? ram_1_80 : _GEN_986; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2524 = ~quene ? ram_1_81 : _GEN_987; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2525 = ~quene ? ram_1_82 : _GEN_988; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2526 = ~quene ? ram_1_83 : _GEN_989; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2527 = ~quene ? ram_1_84 : _GEN_990; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2528 = ~quene ? ram_1_85 : _GEN_991; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2529 = ~quene ? ram_1_86 : _GEN_992; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2530 = ~quene ? ram_1_87 : _GEN_993; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2531 = ~quene ? ram_1_88 : _GEN_994; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2532 = ~quene ? ram_1_89 : _GEN_995; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2533 = ~quene ? ram_1_90 : _GEN_996; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2534 = ~quene ? ram_1_91 : _GEN_997; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2535 = ~quene ? ram_1_92 : _GEN_998; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2536 = ~quene ? ram_1_93 : _GEN_999; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2537 = ~quene ? ram_1_94 : _GEN_1000; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2538 = ~quene ? ram_1_95 : _GEN_1001; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2539 = ~quene ? ram_1_96 : _GEN_1002; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2540 = ~quene ? ram_1_97 : _GEN_1003; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2541 = ~quene ? ram_1_98 : _GEN_1004; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2542 = ~quene ? ram_1_99 : _GEN_1005; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2543 = ~quene ? ram_1_100 : _GEN_1006; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2544 = ~quene ? ram_1_101 : _GEN_1007; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2545 = ~quene ? ram_1_102 : _GEN_1008; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2546 = ~quene ? ram_1_103 : _GEN_1009; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2547 = ~quene ? ram_1_104 : _GEN_1010; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2548 = ~quene ? ram_1_105 : _GEN_1011; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2549 = ~quene ? ram_1_106 : _GEN_1012; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2550 = ~quene ? ram_1_107 : _GEN_1013; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2551 = ~quene ? ram_1_108 : _GEN_1014; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2552 = ~quene ? ram_1_109 : _GEN_1015; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2553 = ~quene ? ram_1_110 : _GEN_1016; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2554 = ~quene ? ram_1_111 : _GEN_1017; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2555 = ~quene ? ram_1_112 : _GEN_1018; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2556 = ~quene ? ram_1_113 : _GEN_1019; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2557 = ~quene ? ram_1_114 : _GEN_1020; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2558 = ~quene ? ram_1_115 : _GEN_1021; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2559 = ~quene ? ram_1_116 : _GEN_1022; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2560 = ~quene ? ram_1_117 : _GEN_1023; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2561 = ~quene ? ram_1_118 : _GEN_1024; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2562 = ~quene ? ram_1_119 : _GEN_1025; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2563 = ~quene ? ram_1_120 : _GEN_1026; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2564 = ~quene ? ram_1_121 : _GEN_1027; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2565 = ~quene ? ram_1_122 : _GEN_1028; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2566 = ~quene ? ram_1_123 : _GEN_1029; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2567 = ~quene ? ram_1_124 : _GEN_1030; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2568 = ~quene ? ram_1_125 : _GEN_1031; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2569 = ~quene ? ram_1_126 : _GEN_1032; // @[i_cache.scala 18:24 97:34]
  wire [63:0] _GEN_2570 = ~quene ? ram_1_127 : _GEN_1033; // @[i_cache.scala 18:24 97:34]
  wire [31:0] _GEN_2571 = ~quene ? tag_1_0 : _GEN_1034; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2572 = ~quene ? tag_1_1 : _GEN_1035; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2573 = ~quene ? tag_1_2 : _GEN_1036; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2574 = ~quene ? tag_1_3 : _GEN_1037; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2575 = ~quene ? tag_1_4 : _GEN_1038; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2576 = ~quene ? tag_1_5 : _GEN_1039; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2577 = ~quene ? tag_1_6 : _GEN_1040; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2578 = ~quene ? tag_1_7 : _GEN_1041; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2579 = ~quene ? tag_1_8 : _GEN_1042; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2580 = ~quene ? tag_1_9 : _GEN_1043; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2581 = ~quene ? tag_1_10 : _GEN_1044; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2582 = ~quene ? tag_1_11 : _GEN_1045; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2583 = ~quene ? tag_1_12 : _GEN_1046; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2584 = ~quene ? tag_1_13 : _GEN_1047; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2585 = ~quene ? tag_1_14 : _GEN_1048; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2586 = ~quene ? tag_1_15 : _GEN_1049; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2587 = ~quene ? tag_1_16 : _GEN_1050; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2588 = ~quene ? tag_1_17 : _GEN_1051; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2589 = ~quene ? tag_1_18 : _GEN_1052; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2590 = ~quene ? tag_1_19 : _GEN_1053; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2591 = ~quene ? tag_1_20 : _GEN_1054; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2592 = ~quene ? tag_1_21 : _GEN_1055; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2593 = ~quene ? tag_1_22 : _GEN_1056; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2594 = ~quene ? tag_1_23 : _GEN_1057; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2595 = ~quene ? tag_1_24 : _GEN_1058; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2596 = ~quene ? tag_1_25 : _GEN_1059; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2597 = ~quene ? tag_1_26 : _GEN_1060; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2598 = ~quene ? tag_1_27 : _GEN_1061; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2599 = ~quene ? tag_1_28 : _GEN_1062; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2600 = ~quene ? tag_1_29 : _GEN_1063; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2601 = ~quene ? tag_1_30 : _GEN_1064; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2602 = ~quene ? tag_1_31 : _GEN_1065; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2603 = ~quene ? tag_1_32 : _GEN_1066; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2604 = ~quene ? tag_1_33 : _GEN_1067; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2605 = ~quene ? tag_1_34 : _GEN_1068; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2606 = ~quene ? tag_1_35 : _GEN_1069; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2607 = ~quene ? tag_1_36 : _GEN_1070; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2608 = ~quene ? tag_1_37 : _GEN_1071; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2609 = ~quene ? tag_1_38 : _GEN_1072; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2610 = ~quene ? tag_1_39 : _GEN_1073; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2611 = ~quene ? tag_1_40 : _GEN_1074; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2612 = ~quene ? tag_1_41 : _GEN_1075; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2613 = ~quene ? tag_1_42 : _GEN_1076; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2614 = ~quene ? tag_1_43 : _GEN_1077; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2615 = ~quene ? tag_1_44 : _GEN_1078; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2616 = ~quene ? tag_1_45 : _GEN_1079; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2617 = ~quene ? tag_1_46 : _GEN_1080; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2618 = ~quene ? tag_1_47 : _GEN_1081; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2619 = ~quene ? tag_1_48 : _GEN_1082; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2620 = ~quene ? tag_1_49 : _GEN_1083; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2621 = ~quene ? tag_1_50 : _GEN_1084; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2622 = ~quene ? tag_1_51 : _GEN_1085; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2623 = ~quene ? tag_1_52 : _GEN_1086; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2624 = ~quene ? tag_1_53 : _GEN_1087; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2625 = ~quene ? tag_1_54 : _GEN_1088; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2626 = ~quene ? tag_1_55 : _GEN_1089; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2627 = ~quene ? tag_1_56 : _GEN_1090; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2628 = ~quene ? tag_1_57 : _GEN_1091; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2629 = ~quene ? tag_1_58 : _GEN_1092; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2630 = ~quene ? tag_1_59 : _GEN_1093; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2631 = ~quene ? tag_1_60 : _GEN_1094; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2632 = ~quene ? tag_1_61 : _GEN_1095; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2633 = ~quene ? tag_1_62 : _GEN_1096; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2634 = ~quene ? tag_1_63 : _GEN_1097; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2635 = ~quene ? tag_1_64 : _GEN_1098; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2636 = ~quene ? tag_1_65 : _GEN_1099; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2637 = ~quene ? tag_1_66 : _GEN_1100; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2638 = ~quene ? tag_1_67 : _GEN_1101; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2639 = ~quene ? tag_1_68 : _GEN_1102; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2640 = ~quene ? tag_1_69 : _GEN_1103; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2641 = ~quene ? tag_1_70 : _GEN_1104; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2642 = ~quene ? tag_1_71 : _GEN_1105; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2643 = ~quene ? tag_1_72 : _GEN_1106; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2644 = ~quene ? tag_1_73 : _GEN_1107; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2645 = ~quene ? tag_1_74 : _GEN_1108; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2646 = ~quene ? tag_1_75 : _GEN_1109; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2647 = ~quene ? tag_1_76 : _GEN_1110; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2648 = ~quene ? tag_1_77 : _GEN_1111; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2649 = ~quene ? tag_1_78 : _GEN_1112; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2650 = ~quene ? tag_1_79 : _GEN_1113; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2651 = ~quene ? tag_1_80 : _GEN_1114; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2652 = ~quene ? tag_1_81 : _GEN_1115; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2653 = ~quene ? tag_1_82 : _GEN_1116; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2654 = ~quene ? tag_1_83 : _GEN_1117; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2655 = ~quene ? tag_1_84 : _GEN_1118; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2656 = ~quene ? tag_1_85 : _GEN_1119; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2657 = ~quene ? tag_1_86 : _GEN_1120; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2658 = ~quene ? tag_1_87 : _GEN_1121; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2659 = ~quene ? tag_1_88 : _GEN_1122; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2660 = ~quene ? tag_1_89 : _GEN_1123; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2661 = ~quene ? tag_1_90 : _GEN_1124; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2662 = ~quene ? tag_1_91 : _GEN_1125; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2663 = ~quene ? tag_1_92 : _GEN_1126; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2664 = ~quene ? tag_1_93 : _GEN_1127; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2665 = ~quene ? tag_1_94 : _GEN_1128; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2666 = ~quene ? tag_1_95 : _GEN_1129; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2667 = ~quene ? tag_1_96 : _GEN_1130; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2668 = ~quene ? tag_1_97 : _GEN_1131; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2669 = ~quene ? tag_1_98 : _GEN_1132; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2670 = ~quene ? tag_1_99 : _GEN_1133; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2671 = ~quene ? tag_1_100 : _GEN_1134; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2672 = ~quene ? tag_1_101 : _GEN_1135; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2673 = ~quene ? tag_1_102 : _GEN_1136; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2674 = ~quene ? tag_1_103 : _GEN_1137; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2675 = ~quene ? tag_1_104 : _GEN_1138; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2676 = ~quene ? tag_1_105 : _GEN_1139; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2677 = ~quene ? tag_1_106 : _GEN_1140; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2678 = ~quene ? tag_1_107 : _GEN_1141; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2679 = ~quene ? tag_1_108 : _GEN_1142; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2680 = ~quene ? tag_1_109 : _GEN_1143; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2681 = ~quene ? tag_1_110 : _GEN_1144; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2682 = ~quene ? tag_1_111 : _GEN_1145; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2683 = ~quene ? tag_1_112 : _GEN_1146; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2684 = ~quene ? tag_1_113 : _GEN_1147; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2685 = ~quene ? tag_1_114 : _GEN_1148; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2686 = ~quene ? tag_1_115 : _GEN_1149; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2687 = ~quene ? tag_1_116 : _GEN_1150; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2688 = ~quene ? tag_1_117 : _GEN_1151; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2689 = ~quene ? tag_1_118 : _GEN_1152; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2690 = ~quene ? tag_1_119 : _GEN_1153; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2691 = ~quene ? tag_1_120 : _GEN_1154; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2692 = ~quene ? tag_1_121 : _GEN_1155; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2693 = ~quene ? tag_1_122 : _GEN_1156; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2694 = ~quene ? tag_1_123 : _GEN_1157; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2695 = ~quene ? tag_1_124 : _GEN_1158; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2696 = ~quene ? tag_1_125 : _GEN_1159; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2697 = ~quene ? tag_1_126 : _GEN_1160; // @[i_cache.scala 20:24 97:34]
  wire [31:0] _GEN_2698 = ~quene ? tag_1_127 : _GEN_1161; // @[i_cache.scala 20:24 97:34]
  wire  _GEN_2699 = ~quene ? valid_1_0 : _GEN_1162; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2700 = ~quene ? valid_1_1 : _GEN_1163; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2701 = ~quene ? valid_1_2 : _GEN_1164; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2702 = ~quene ? valid_1_3 : _GEN_1165; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2703 = ~quene ? valid_1_4 : _GEN_1166; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2704 = ~quene ? valid_1_5 : _GEN_1167; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2705 = ~quene ? valid_1_6 : _GEN_1168; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2706 = ~quene ? valid_1_7 : _GEN_1169; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2707 = ~quene ? valid_1_8 : _GEN_1170; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2708 = ~quene ? valid_1_9 : _GEN_1171; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2709 = ~quene ? valid_1_10 : _GEN_1172; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2710 = ~quene ? valid_1_11 : _GEN_1173; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2711 = ~quene ? valid_1_12 : _GEN_1174; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2712 = ~quene ? valid_1_13 : _GEN_1175; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2713 = ~quene ? valid_1_14 : _GEN_1176; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2714 = ~quene ? valid_1_15 : _GEN_1177; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2715 = ~quene ? valid_1_16 : _GEN_1178; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2716 = ~quene ? valid_1_17 : _GEN_1179; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2717 = ~quene ? valid_1_18 : _GEN_1180; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2718 = ~quene ? valid_1_19 : _GEN_1181; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2719 = ~quene ? valid_1_20 : _GEN_1182; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2720 = ~quene ? valid_1_21 : _GEN_1183; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2721 = ~quene ? valid_1_22 : _GEN_1184; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2722 = ~quene ? valid_1_23 : _GEN_1185; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2723 = ~quene ? valid_1_24 : _GEN_1186; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2724 = ~quene ? valid_1_25 : _GEN_1187; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2725 = ~quene ? valid_1_26 : _GEN_1188; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2726 = ~quene ? valid_1_27 : _GEN_1189; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2727 = ~quene ? valid_1_28 : _GEN_1190; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2728 = ~quene ? valid_1_29 : _GEN_1191; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2729 = ~quene ? valid_1_30 : _GEN_1192; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2730 = ~quene ? valid_1_31 : _GEN_1193; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2731 = ~quene ? valid_1_32 : _GEN_1194; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2732 = ~quene ? valid_1_33 : _GEN_1195; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2733 = ~quene ? valid_1_34 : _GEN_1196; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2734 = ~quene ? valid_1_35 : _GEN_1197; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2735 = ~quene ? valid_1_36 : _GEN_1198; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2736 = ~quene ? valid_1_37 : _GEN_1199; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2737 = ~quene ? valid_1_38 : _GEN_1200; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2738 = ~quene ? valid_1_39 : _GEN_1201; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2739 = ~quene ? valid_1_40 : _GEN_1202; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2740 = ~quene ? valid_1_41 : _GEN_1203; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2741 = ~quene ? valid_1_42 : _GEN_1204; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2742 = ~quene ? valid_1_43 : _GEN_1205; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2743 = ~quene ? valid_1_44 : _GEN_1206; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2744 = ~quene ? valid_1_45 : _GEN_1207; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2745 = ~quene ? valid_1_46 : _GEN_1208; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2746 = ~quene ? valid_1_47 : _GEN_1209; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2747 = ~quene ? valid_1_48 : _GEN_1210; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2748 = ~quene ? valid_1_49 : _GEN_1211; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2749 = ~quene ? valid_1_50 : _GEN_1212; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2750 = ~quene ? valid_1_51 : _GEN_1213; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2751 = ~quene ? valid_1_52 : _GEN_1214; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2752 = ~quene ? valid_1_53 : _GEN_1215; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2753 = ~quene ? valid_1_54 : _GEN_1216; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2754 = ~quene ? valid_1_55 : _GEN_1217; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2755 = ~quene ? valid_1_56 : _GEN_1218; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2756 = ~quene ? valid_1_57 : _GEN_1219; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2757 = ~quene ? valid_1_58 : _GEN_1220; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2758 = ~quene ? valid_1_59 : _GEN_1221; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2759 = ~quene ? valid_1_60 : _GEN_1222; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2760 = ~quene ? valid_1_61 : _GEN_1223; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2761 = ~quene ? valid_1_62 : _GEN_1224; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2762 = ~quene ? valid_1_63 : _GEN_1225; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2763 = ~quene ? valid_1_64 : _GEN_1226; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2764 = ~quene ? valid_1_65 : _GEN_1227; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2765 = ~quene ? valid_1_66 : _GEN_1228; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2766 = ~quene ? valid_1_67 : _GEN_1229; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2767 = ~quene ? valid_1_68 : _GEN_1230; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2768 = ~quene ? valid_1_69 : _GEN_1231; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2769 = ~quene ? valid_1_70 : _GEN_1232; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2770 = ~quene ? valid_1_71 : _GEN_1233; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2771 = ~quene ? valid_1_72 : _GEN_1234; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2772 = ~quene ? valid_1_73 : _GEN_1235; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2773 = ~quene ? valid_1_74 : _GEN_1236; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2774 = ~quene ? valid_1_75 : _GEN_1237; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2775 = ~quene ? valid_1_76 : _GEN_1238; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2776 = ~quene ? valid_1_77 : _GEN_1239; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2777 = ~quene ? valid_1_78 : _GEN_1240; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2778 = ~quene ? valid_1_79 : _GEN_1241; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2779 = ~quene ? valid_1_80 : _GEN_1242; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2780 = ~quene ? valid_1_81 : _GEN_1243; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2781 = ~quene ? valid_1_82 : _GEN_1244; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2782 = ~quene ? valid_1_83 : _GEN_1245; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2783 = ~quene ? valid_1_84 : _GEN_1246; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2784 = ~quene ? valid_1_85 : _GEN_1247; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2785 = ~quene ? valid_1_86 : _GEN_1248; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2786 = ~quene ? valid_1_87 : _GEN_1249; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2787 = ~quene ? valid_1_88 : _GEN_1250; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2788 = ~quene ? valid_1_89 : _GEN_1251; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2789 = ~quene ? valid_1_90 : _GEN_1252; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2790 = ~quene ? valid_1_91 : _GEN_1253; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2791 = ~quene ? valid_1_92 : _GEN_1254; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2792 = ~quene ? valid_1_93 : _GEN_1255; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2793 = ~quene ? valid_1_94 : _GEN_1256; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2794 = ~quene ? valid_1_95 : _GEN_1257; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2795 = ~quene ? valid_1_96 : _GEN_1258; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2796 = ~quene ? valid_1_97 : _GEN_1259; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2797 = ~quene ? valid_1_98 : _GEN_1260; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2798 = ~quene ? valid_1_99 : _GEN_1261; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2799 = ~quene ? valid_1_100 : _GEN_1262; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2800 = ~quene ? valid_1_101 : _GEN_1263; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2801 = ~quene ? valid_1_102 : _GEN_1264; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2802 = ~quene ? valid_1_103 : _GEN_1265; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2803 = ~quene ? valid_1_104 : _GEN_1266; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2804 = ~quene ? valid_1_105 : _GEN_1267; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2805 = ~quene ? valid_1_106 : _GEN_1268; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2806 = ~quene ? valid_1_107 : _GEN_1269; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2807 = ~quene ? valid_1_108 : _GEN_1270; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2808 = ~quene ? valid_1_109 : _GEN_1271; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2809 = ~quene ? valid_1_110 : _GEN_1272; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2810 = ~quene ? valid_1_111 : _GEN_1273; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2811 = ~quene ? valid_1_112 : _GEN_1274; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2812 = ~quene ? valid_1_113 : _GEN_1275; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2813 = ~quene ? valid_1_114 : _GEN_1276; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2814 = ~quene ? valid_1_115 : _GEN_1277; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2815 = ~quene ? valid_1_116 : _GEN_1278; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2816 = ~quene ? valid_1_117 : _GEN_1279; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2817 = ~quene ? valid_1_118 : _GEN_1280; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2818 = ~quene ? valid_1_119 : _GEN_1281; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2819 = ~quene ? valid_1_120 : _GEN_1282; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2820 = ~quene ? valid_1_121 : _GEN_1283; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2821 = ~quene ? valid_1_122 : _GEN_1284; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2822 = ~quene ? valid_1_123 : _GEN_1285; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2823 = ~quene ? valid_1_124 : _GEN_1286; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2824 = ~quene ? valid_1_125 : _GEN_1287; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2825 = ~quene ? valid_1_126 : _GEN_1288; // @[i_cache.scala 22:26 97:34]
  wire  _GEN_2826 = ~quene ? valid_1_127 : _GEN_1289; // @[i_cache.scala 22:26 97:34]
  wire [63:0] _GEN_2827 = unuse_way == 2'h2 ? _GEN_906 : _GEN_2443; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2828 = unuse_way == 2'h2 ? _GEN_907 : _GEN_2444; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2829 = unuse_way == 2'h2 ? _GEN_908 : _GEN_2445; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2830 = unuse_way == 2'h2 ? _GEN_909 : _GEN_2446; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2831 = unuse_way == 2'h2 ? _GEN_910 : _GEN_2447; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2832 = unuse_way == 2'h2 ? _GEN_911 : _GEN_2448; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2833 = unuse_way == 2'h2 ? _GEN_912 : _GEN_2449; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2834 = unuse_way == 2'h2 ? _GEN_913 : _GEN_2450; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2835 = unuse_way == 2'h2 ? _GEN_914 : _GEN_2451; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2836 = unuse_way == 2'h2 ? _GEN_915 : _GEN_2452; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2837 = unuse_way == 2'h2 ? _GEN_916 : _GEN_2453; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2838 = unuse_way == 2'h2 ? _GEN_917 : _GEN_2454; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2839 = unuse_way == 2'h2 ? _GEN_918 : _GEN_2455; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2840 = unuse_way == 2'h2 ? _GEN_919 : _GEN_2456; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2841 = unuse_way == 2'h2 ? _GEN_920 : _GEN_2457; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2842 = unuse_way == 2'h2 ? _GEN_921 : _GEN_2458; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2843 = unuse_way == 2'h2 ? _GEN_922 : _GEN_2459; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2844 = unuse_way == 2'h2 ? _GEN_923 : _GEN_2460; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2845 = unuse_way == 2'h2 ? _GEN_924 : _GEN_2461; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2846 = unuse_way == 2'h2 ? _GEN_925 : _GEN_2462; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2847 = unuse_way == 2'h2 ? _GEN_926 : _GEN_2463; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2848 = unuse_way == 2'h2 ? _GEN_927 : _GEN_2464; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2849 = unuse_way == 2'h2 ? _GEN_928 : _GEN_2465; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2850 = unuse_way == 2'h2 ? _GEN_929 : _GEN_2466; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2851 = unuse_way == 2'h2 ? _GEN_930 : _GEN_2467; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2852 = unuse_way == 2'h2 ? _GEN_931 : _GEN_2468; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2853 = unuse_way == 2'h2 ? _GEN_932 : _GEN_2469; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2854 = unuse_way == 2'h2 ? _GEN_933 : _GEN_2470; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2855 = unuse_way == 2'h2 ? _GEN_934 : _GEN_2471; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2856 = unuse_way == 2'h2 ? _GEN_935 : _GEN_2472; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2857 = unuse_way == 2'h2 ? _GEN_936 : _GEN_2473; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2858 = unuse_way == 2'h2 ? _GEN_937 : _GEN_2474; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2859 = unuse_way == 2'h2 ? _GEN_938 : _GEN_2475; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2860 = unuse_way == 2'h2 ? _GEN_939 : _GEN_2476; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2861 = unuse_way == 2'h2 ? _GEN_940 : _GEN_2477; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2862 = unuse_way == 2'h2 ? _GEN_941 : _GEN_2478; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2863 = unuse_way == 2'h2 ? _GEN_942 : _GEN_2479; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2864 = unuse_way == 2'h2 ? _GEN_943 : _GEN_2480; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2865 = unuse_way == 2'h2 ? _GEN_944 : _GEN_2481; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2866 = unuse_way == 2'h2 ? _GEN_945 : _GEN_2482; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2867 = unuse_way == 2'h2 ? _GEN_946 : _GEN_2483; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2868 = unuse_way == 2'h2 ? _GEN_947 : _GEN_2484; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2869 = unuse_way == 2'h2 ? _GEN_948 : _GEN_2485; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2870 = unuse_way == 2'h2 ? _GEN_949 : _GEN_2486; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2871 = unuse_way == 2'h2 ? _GEN_950 : _GEN_2487; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2872 = unuse_way == 2'h2 ? _GEN_951 : _GEN_2488; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2873 = unuse_way == 2'h2 ? _GEN_952 : _GEN_2489; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2874 = unuse_way == 2'h2 ? _GEN_953 : _GEN_2490; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2875 = unuse_way == 2'h2 ? _GEN_954 : _GEN_2491; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2876 = unuse_way == 2'h2 ? _GEN_955 : _GEN_2492; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2877 = unuse_way == 2'h2 ? _GEN_956 : _GEN_2493; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2878 = unuse_way == 2'h2 ? _GEN_957 : _GEN_2494; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2879 = unuse_way == 2'h2 ? _GEN_958 : _GEN_2495; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2880 = unuse_way == 2'h2 ? _GEN_959 : _GEN_2496; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2881 = unuse_way == 2'h2 ? _GEN_960 : _GEN_2497; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2882 = unuse_way == 2'h2 ? _GEN_961 : _GEN_2498; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2883 = unuse_way == 2'h2 ? _GEN_962 : _GEN_2499; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2884 = unuse_way == 2'h2 ? _GEN_963 : _GEN_2500; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2885 = unuse_way == 2'h2 ? _GEN_964 : _GEN_2501; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2886 = unuse_way == 2'h2 ? _GEN_965 : _GEN_2502; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2887 = unuse_way == 2'h2 ? _GEN_966 : _GEN_2503; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2888 = unuse_way == 2'h2 ? _GEN_967 : _GEN_2504; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2889 = unuse_way == 2'h2 ? _GEN_968 : _GEN_2505; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2890 = unuse_way == 2'h2 ? _GEN_969 : _GEN_2506; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2891 = unuse_way == 2'h2 ? _GEN_970 : _GEN_2507; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2892 = unuse_way == 2'h2 ? _GEN_971 : _GEN_2508; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2893 = unuse_way == 2'h2 ? _GEN_972 : _GEN_2509; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2894 = unuse_way == 2'h2 ? _GEN_973 : _GEN_2510; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2895 = unuse_way == 2'h2 ? _GEN_974 : _GEN_2511; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2896 = unuse_way == 2'h2 ? _GEN_975 : _GEN_2512; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2897 = unuse_way == 2'h2 ? _GEN_976 : _GEN_2513; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2898 = unuse_way == 2'h2 ? _GEN_977 : _GEN_2514; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2899 = unuse_way == 2'h2 ? _GEN_978 : _GEN_2515; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2900 = unuse_way == 2'h2 ? _GEN_979 : _GEN_2516; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2901 = unuse_way == 2'h2 ? _GEN_980 : _GEN_2517; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2902 = unuse_way == 2'h2 ? _GEN_981 : _GEN_2518; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2903 = unuse_way == 2'h2 ? _GEN_982 : _GEN_2519; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2904 = unuse_way == 2'h2 ? _GEN_983 : _GEN_2520; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2905 = unuse_way == 2'h2 ? _GEN_984 : _GEN_2521; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2906 = unuse_way == 2'h2 ? _GEN_985 : _GEN_2522; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2907 = unuse_way == 2'h2 ? _GEN_986 : _GEN_2523; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2908 = unuse_way == 2'h2 ? _GEN_987 : _GEN_2524; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2909 = unuse_way == 2'h2 ? _GEN_988 : _GEN_2525; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2910 = unuse_way == 2'h2 ? _GEN_989 : _GEN_2526; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2911 = unuse_way == 2'h2 ? _GEN_990 : _GEN_2527; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2912 = unuse_way == 2'h2 ? _GEN_991 : _GEN_2528; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2913 = unuse_way == 2'h2 ? _GEN_992 : _GEN_2529; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2914 = unuse_way == 2'h2 ? _GEN_993 : _GEN_2530; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2915 = unuse_way == 2'h2 ? _GEN_994 : _GEN_2531; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2916 = unuse_way == 2'h2 ? _GEN_995 : _GEN_2532; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2917 = unuse_way == 2'h2 ? _GEN_996 : _GEN_2533; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2918 = unuse_way == 2'h2 ? _GEN_997 : _GEN_2534; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2919 = unuse_way == 2'h2 ? _GEN_998 : _GEN_2535; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2920 = unuse_way == 2'h2 ? _GEN_999 : _GEN_2536; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2921 = unuse_way == 2'h2 ? _GEN_1000 : _GEN_2537; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2922 = unuse_way == 2'h2 ? _GEN_1001 : _GEN_2538; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2923 = unuse_way == 2'h2 ? _GEN_1002 : _GEN_2539; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2924 = unuse_way == 2'h2 ? _GEN_1003 : _GEN_2540; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2925 = unuse_way == 2'h2 ? _GEN_1004 : _GEN_2541; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2926 = unuse_way == 2'h2 ? _GEN_1005 : _GEN_2542; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2927 = unuse_way == 2'h2 ? _GEN_1006 : _GEN_2543; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2928 = unuse_way == 2'h2 ? _GEN_1007 : _GEN_2544; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2929 = unuse_way == 2'h2 ? _GEN_1008 : _GEN_2545; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2930 = unuse_way == 2'h2 ? _GEN_1009 : _GEN_2546; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2931 = unuse_way == 2'h2 ? _GEN_1010 : _GEN_2547; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2932 = unuse_way == 2'h2 ? _GEN_1011 : _GEN_2548; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2933 = unuse_way == 2'h2 ? _GEN_1012 : _GEN_2549; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2934 = unuse_way == 2'h2 ? _GEN_1013 : _GEN_2550; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2935 = unuse_way == 2'h2 ? _GEN_1014 : _GEN_2551; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2936 = unuse_way == 2'h2 ? _GEN_1015 : _GEN_2552; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2937 = unuse_way == 2'h2 ? _GEN_1016 : _GEN_2553; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2938 = unuse_way == 2'h2 ? _GEN_1017 : _GEN_2554; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2939 = unuse_way == 2'h2 ? _GEN_1018 : _GEN_2555; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2940 = unuse_way == 2'h2 ? _GEN_1019 : _GEN_2556; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2941 = unuse_way == 2'h2 ? _GEN_1020 : _GEN_2557; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2942 = unuse_way == 2'h2 ? _GEN_1021 : _GEN_2558; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2943 = unuse_way == 2'h2 ? _GEN_1022 : _GEN_2559; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2944 = unuse_way == 2'h2 ? _GEN_1023 : _GEN_2560; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2945 = unuse_way == 2'h2 ? _GEN_1024 : _GEN_2561; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2946 = unuse_way == 2'h2 ? _GEN_1025 : _GEN_2562; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2947 = unuse_way == 2'h2 ? _GEN_1026 : _GEN_2563; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2948 = unuse_way == 2'h2 ? _GEN_1027 : _GEN_2564; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2949 = unuse_way == 2'h2 ? _GEN_1028 : _GEN_2565; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2950 = unuse_way == 2'h2 ? _GEN_1029 : _GEN_2566; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2951 = unuse_way == 2'h2 ? _GEN_1030 : _GEN_2567; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2952 = unuse_way == 2'h2 ? _GEN_1031 : _GEN_2568; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2953 = unuse_way == 2'h2 ? _GEN_1032 : _GEN_2569; // @[i_cache.scala 91:40]
  wire [63:0] _GEN_2954 = unuse_way == 2'h2 ? _GEN_1033 : _GEN_2570; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2955 = unuse_way == 2'h2 ? _GEN_1034 : _GEN_2571; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2956 = unuse_way == 2'h2 ? _GEN_1035 : _GEN_2572; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2957 = unuse_way == 2'h2 ? _GEN_1036 : _GEN_2573; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2958 = unuse_way == 2'h2 ? _GEN_1037 : _GEN_2574; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2959 = unuse_way == 2'h2 ? _GEN_1038 : _GEN_2575; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2960 = unuse_way == 2'h2 ? _GEN_1039 : _GEN_2576; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2961 = unuse_way == 2'h2 ? _GEN_1040 : _GEN_2577; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2962 = unuse_way == 2'h2 ? _GEN_1041 : _GEN_2578; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2963 = unuse_way == 2'h2 ? _GEN_1042 : _GEN_2579; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2964 = unuse_way == 2'h2 ? _GEN_1043 : _GEN_2580; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2965 = unuse_way == 2'h2 ? _GEN_1044 : _GEN_2581; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2966 = unuse_way == 2'h2 ? _GEN_1045 : _GEN_2582; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2967 = unuse_way == 2'h2 ? _GEN_1046 : _GEN_2583; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2968 = unuse_way == 2'h2 ? _GEN_1047 : _GEN_2584; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2969 = unuse_way == 2'h2 ? _GEN_1048 : _GEN_2585; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2970 = unuse_way == 2'h2 ? _GEN_1049 : _GEN_2586; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2971 = unuse_way == 2'h2 ? _GEN_1050 : _GEN_2587; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2972 = unuse_way == 2'h2 ? _GEN_1051 : _GEN_2588; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2973 = unuse_way == 2'h2 ? _GEN_1052 : _GEN_2589; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2974 = unuse_way == 2'h2 ? _GEN_1053 : _GEN_2590; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2975 = unuse_way == 2'h2 ? _GEN_1054 : _GEN_2591; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2976 = unuse_way == 2'h2 ? _GEN_1055 : _GEN_2592; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2977 = unuse_way == 2'h2 ? _GEN_1056 : _GEN_2593; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2978 = unuse_way == 2'h2 ? _GEN_1057 : _GEN_2594; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2979 = unuse_way == 2'h2 ? _GEN_1058 : _GEN_2595; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2980 = unuse_way == 2'h2 ? _GEN_1059 : _GEN_2596; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2981 = unuse_way == 2'h2 ? _GEN_1060 : _GEN_2597; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2982 = unuse_way == 2'h2 ? _GEN_1061 : _GEN_2598; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2983 = unuse_way == 2'h2 ? _GEN_1062 : _GEN_2599; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2984 = unuse_way == 2'h2 ? _GEN_1063 : _GEN_2600; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2985 = unuse_way == 2'h2 ? _GEN_1064 : _GEN_2601; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2986 = unuse_way == 2'h2 ? _GEN_1065 : _GEN_2602; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2987 = unuse_way == 2'h2 ? _GEN_1066 : _GEN_2603; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2988 = unuse_way == 2'h2 ? _GEN_1067 : _GEN_2604; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2989 = unuse_way == 2'h2 ? _GEN_1068 : _GEN_2605; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2990 = unuse_way == 2'h2 ? _GEN_1069 : _GEN_2606; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2991 = unuse_way == 2'h2 ? _GEN_1070 : _GEN_2607; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2992 = unuse_way == 2'h2 ? _GEN_1071 : _GEN_2608; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2993 = unuse_way == 2'h2 ? _GEN_1072 : _GEN_2609; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2994 = unuse_way == 2'h2 ? _GEN_1073 : _GEN_2610; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2995 = unuse_way == 2'h2 ? _GEN_1074 : _GEN_2611; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2996 = unuse_way == 2'h2 ? _GEN_1075 : _GEN_2612; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2997 = unuse_way == 2'h2 ? _GEN_1076 : _GEN_2613; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2998 = unuse_way == 2'h2 ? _GEN_1077 : _GEN_2614; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_2999 = unuse_way == 2'h2 ? _GEN_1078 : _GEN_2615; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3000 = unuse_way == 2'h2 ? _GEN_1079 : _GEN_2616; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3001 = unuse_way == 2'h2 ? _GEN_1080 : _GEN_2617; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3002 = unuse_way == 2'h2 ? _GEN_1081 : _GEN_2618; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3003 = unuse_way == 2'h2 ? _GEN_1082 : _GEN_2619; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3004 = unuse_way == 2'h2 ? _GEN_1083 : _GEN_2620; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3005 = unuse_way == 2'h2 ? _GEN_1084 : _GEN_2621; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3006 = unuse_way == 2'h2 ? _GEN_1085 : _GEN_2622; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3007 = unuse_way == 2'h2 ? _GEN_1086 : _GEN_2623; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3008 = unuse_way == 2'h2 ? _GEN_1087 : _GEN_2624; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3009 = unuse_way == 2'h2 ? _GEN_1088 : _GEN_2625; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3010 = unuse_way == 2'h2 ? _GEN_1089 : _GEN_2626; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3011 = unuse_way == 2'h2 ? _GEN_1090 : _GEN_2627; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3012 = unuse_way == 2'h2 ? _GEN_1091 : _GEN_2628; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3013 = unuse_way == 2'h2 ? _GEN_1092 : _GEN_2629; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3014 = unuse_way == 2'h2 ? _GEN_1093 : _GEN_2630; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3015 = unuse_way == 2'h2 ? _GEN_1094 : _GEN_2631; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3016 = unuse_way == 2'h2 ? _GEN_1095 : _GEN_2632; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3017 = unuse_way == 2'h2 ? _GEN_1096 : _GEN_2633; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3018 = unuse_way == 2'h2 ? _GEN_1097 : _GEN_2634; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3019 = unuse_way == 2'h2 ? _GEN_1098 : _GEN_2635; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3020 = unuse_way == 2'h2 ? _GEN_1099 : _GEN_2636; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3021 = unuse_way == 2'h2 ? _GEN_1100 : _GEN_2637; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3022 = unuse_way == 2'h2 ? _GEN_1101 : _GEN_2638; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3023 = unuse_way == 2'h2 ? _GEN_1102 : _GEN_2639; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3024 = unuse_way == 2'h2 ? _GEN_1103 : _GEN_2640; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3025 = unuse_way == 2'h2 ? _GEN_1104 : _GEN_2641; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3026 = unuse_way == 2'h2 ? _GEN_1105 : _GEN_2642; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3027 = unuse_way == 2'h2 ? _GEN_1106 : _GEN_2643; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3028 = unuse_way == 2'h2 ? _GEN_1107 : _GEN_2644; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3029 = unuse_way == 2'h2 ? _GEN_1108 : _GEN_2645; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3030 = unuse_way == 2'h2 ? _GEN_1109 : _GEN_2646; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3031 = unuse_way == 2'h2 ? _GEN_1110 : _GEN_2647; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3032 = unuse_way == 2'h2 ? _GEN_1111 : _GEN_2648; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3033 = unuse_way == 2'h2 ? _GEN_1112 : _GEN_2649; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3034 = unuse_way == 2'h2 ? _GEN_1113 : _GEN_2650; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3035 = unuse_way == 2'h2 ? _GEN_1114 : _GEN_2651; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3036 = unuse_way == 2'h2 ? _GEN_1115 : _GEN_2652; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3037 = unuse_way == 2'h2 ? _GEN_1116 : _GEN_2653; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3038 = unuse_way == 2'h2 ? _GEN_1117 : _GEN_2654; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3039 = unuse_way == 2'h2 ? _GEN_1118 : _GEN_2655; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3040 = unuse_way == 2'h2 ? _GEN_1119 : _GEN_2656; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3041 = unuse_way == 2'h2 ? _GEN_1120 : _GEN_2657; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3042 = unuse_way == 2'h2 ? _GEN_1121 : _GEN_2658; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3043 = unuse_way == 2'h2 ? _GEN_1122 : _GEN_2659; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3044 = unuse_way == 2'h2 ? _GEN_1123 : _GEN_2660; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3045 = unuse_way == 2'h2 ? _GEN_1124 : _GEN_2661; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3046 = unuse_way == 2'h2 ? _GEN_1125 : _GEN_2662; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3047 = unuse_way == 2'h2 ? _GEN_1126 : _GEN_2663; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3048 = unuse_way == 2'h2 ? _GEN_1127 : _GEN_2664; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3049 = unuse_way == 2'h2 ? _GEN_1128 : _GEN_2665; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3050 = unuse_way == 2'h2 ? _GEN_1129 : _GEN_2666; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3051 = unuse_way == 2'h2 ? _GEN_1130 : _GEN_2667; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3052 = unuse_way == 2'h2 ? _GEN_1131 : _GEN_2668; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3053 = unuse_way == 2'h2 ? _GEN_1132 : _GEN_2669; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3054 = unuse_way == 2'h2 ? _GEN_1133 : _GEN_2670; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3055 = unuse_way == 2'h2 ? _GEN_1134 : _GEN_2671; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3056 = unuse_way == 2'h2 ? _GEN_1135 : _GEN_2672; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3057 = unuse_way == 2'h2 ? _GEN_1136 : _GEN_2673; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3058 = unuse_way == 2'h2 ? _GEN_1137 : _GEN_2674; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3059 = unuse_way == 2'h2 ? _GEN_1138 : _GEN_2675; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3060 = unuse_way == 2'h2 ? _GEN_1139 : _GEN_2676; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3061 = unuse_way == 2'h2 ? _GEN_1140 : _GEN_2677; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3062 = unuse_way == 2'h2 ? _GEN_1141 : _GEN_2678; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3063 = unuse_way == 2'h2 ? _GEN_1142 : _GEN_2679; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3064 = unuse_way == 2'h2 ? _GEN_1143 : _GEN_2680; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3065 = unuse_way == 2'h2 ? _GEN_1144 : _GEN_2681; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3066 = unuse_way == 2'h2 ? _GEN_1145 : _GEN_2682; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3067 = unuse_way == 2'h2 ? _GEN_1146 : _GEN_2683; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3068 = unuse_way == 2'h2 ? _GEN_1147 : _GEN_2684; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3069 = unuse_way == 2'h2 ? _GEN_1148 : _GEN_2685; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3070 = unuse_way == 2'h2 ? _GEN_1149 : _GEN_2686; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3071 = unuse_way == 2'h2 ? _GEN_1150 : _GEN_2687; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3072 = unuse_way == 2'h2 ? _GEN_1151 : _GEN_2688; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3073 = unuse_way == 2'h2 ? _GEN_1152 : _GEN_2689; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3074 = unuse_way == 2'h2 ? _GEN_1153 : _GEN_2690; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3075 = unuse_way == 2'h2 ? _GEN_1154 : _GEN_2691; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3076 = unuse_way == 2'h2 ? _GEN_1155 : _GEN_2692; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3077 = unuse_way == 2'h2 ? _GEN_1156 : _GEN_2693; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3078 = unuse_way == 2'h2 ? _GEN_1157 : _GEN_2694; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3079 = unuse_way == 2'h2 ? _GEN_1158 : _GEN_2695; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3080 = unuse_way == 2'h2 ? _GEN_1159 : _GEN_2696; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3081 = unuse_way == 2'h2 ? _GEN_1160 : _GEN_2697; // @[i_cache.scala 91:40]
  wire [31:0] _GEN_3082 = unuse_way == 2'h2 ? _GEN_1161 : _GEN_2698; // @[i_cache.scala 91:40]
  wire  _GEN_3083 = unuse_way == 2'h2 ? _GEN_1162 : _GEN_2699; // @[i_cache.scala 91:40]
  wire  _GEN_3084 = unuse_way == 2'h2 ? _GEN_1163 : _GEN_2700; // @[i_cache.scala 91:40]
  wire  _GEN_3085 = unuse_way == 2'h2 ? _GEN_1164 : _GEN_2701; // @[i_cache.scala 91:40]
  wire  _GEN_3086 = unuse_way == 2'h2 ? _GEN_1165 : _GEN_2702; // @[i_cache.scala 91:40]
  wire  _GEN_3087 = unuse_way == 2'h2 ? _GEN_1166 : _GEN_2703; // @[i_cache.scala 91:40]
  wire  _GEN_3088 = unuse_way == 2'h2 ? _GEN_1167 : _GEN_2704; // @[i_cache.scala 91:40]
  wire  _GEN_3089 = unuse_way == 2'h2 ? _GEN_1168 : _GEN_2705; // @[i_cache.scala 91:40]
  wire  _GEN_3090 = unuse_way == 2'h2 ? _GEN_1169 : _GEN_2706; // @[i_cache.scala 91:40]
  wire  _GEN_3091 = unuse_way == 2'h2 ? _GEN_1170 : _GEN_2707; // @[i_cache.scala 91:40]
  wire  _GEN_3092 = unuse_way == 2'h2 ? _GEN_1171 : _GEN_2708; // @[i_cache.scala 91:40]
  wire  _GEN_3093 = unuse_way == 2'h2 ? _GEN_1172 : _GEN_2709; // @[i_cache.scala 91:40]
  wire  _GEN_3094 = unuse_way == 2'h2 ? _GEN_1173 : _GEN_2710; // @[i_cache.scala 91:40]
  wire  _GEN_3095 = unuse_way == 2'h2 ? _GEN_1174 : _GEN_2711; // @[i_cache.scala 91:40]
  wire  _GEN_3096 = unuse_way == 2'h2 ? _GEN_1175 : _GEN_2712; // @[i_cache.scala 91:40]
  wire  _GEN_3097 = unuse_way == 2'h2 ? _GEN_1176 : _GEN_2713; // @[i_cache.scala 91:40]
  wire  _GEN_3098 = unuse_way == 2'h2 ? _GEN_1177 : _GEN_2714; // @[i_cache.scala 91:40]
  wire  _GEN_3099 = unuse_way == 2'h2 ? _GEN_1178 : _GEN_2715; // @[i_cache.scala 91:40]
  wire  _GEN_3100 = unuse_way == 2'h2 ? _GEN_1179 : _GEN_2716; // @[i_cache.scala 91:40]
  wire  _GEN_3101 = unuse_way == 2'h2 ? _GEN_1180 : _GEN_2717; // @[i_cache.scala 91:40]
  wire  _GEN_3102 = unuse_way == 2'h2 ? _GEN_1181 : _GEN_2718; // @[i_cache.scala 91:40]
  wire  _GEN_3103 = unuse_way == 2'h2 ? _GEN_1182 : _GEN_2719; // @[i_cache.scala 91:40]
  wire  _GEN_3104 = unuse_way == 2'h2 ? _GEN_1183 : _GEN_2720; // @[i_cache.scala 91:40]
  wire  _GEN_3105 = unuse_way == 2'h2 ? _GEN_1184 : _GEN_2721; // @[i_cache.scala 91:40]
  wire  _GEN_3106 = unuse_way == 2'h2 ? _GEN_1185 : _GEN_2722; // @[i_cache.scala 91:40]
  wire  _GEN_3107 = unuse_way == 2'h2 ? _GEN_1186 : _GEN_2723; // @[i_cache.scala 91:40]
  wire  _GEN_3108 = unuse_way == 2'h2 ? _GEN_1187 : _GEN_2724; // @[i_cache.scala 91:40]
  wire  _GEN_3109 = unuse_way == 2'h2 ? _GEN_1188 : _GEN_2725; // @[i_cache.scala 91:40]
  wire  _GEN_3110 = unuse_way == 2'h2 ? _GEN_1189 : _GEN_2726; // @[i_cache.scala 91:40]
  wire  _GEN_3111 = unuse_way == 2'h2 ? _GEN_1190 : _GEN_2727; // @[i_cache.scala 91:40]
  wire  _GEN_3112 = unuse_way == 2'h2 ? _GEN_1191 : _GEN_2728; // @[i_cache.scala 91:40]
  wire  _GEN_3113 = unuse_way == 2'h2 ? _GEN_1192 : _GEN_2729; // @[i_cache.scala 91:40]
  wire  _GEN_3114 = unuse_way == 2'h2 ? _GEN_1193 : _GEN_2730; // @[i_cache.scala 91:40]
  wire  _GEN_3115 = unuse_way == 2'h2 ? _GEN_1194 : _GEN_2731; // @[i_cache.scala 91:40]
  wire  _GEN_3116 = unuse_way == 2'h2 ? _GEN_1195 : _GEN_2732; // @[i_cache.scala 91:40]
  wire  _GEN_3117 = unuse_way == 2'h2 ? _GEN_1196 : _GEN_2733; // @[i_cache.scala 91:40]
  wire  _GEN_3118 = unuse_way == 2'h2 ? _GEN_1197 : _GEN_2734; // @[i_cache.scala 91:40]
  wire  _GEN_3119 = unuse_way == 2'h2 ? _GEN_1198 : _GEN_2735; // @[i_cache.scala 91:40]
  wire  _GEN_3120 = unuse_way == 2'h2 ? _GEN_1199 : _GEN_2736; // @[i_cache.scala 91:40]
  wire  _GEN_3121 = unuse_way == 2'h2 ? _GEN_1200 : _GEN_2737; // @[i_cache.scala 91:40]
  wire  _GEN_3122 = unuse_way == 2'h2 ? _GEN_1201 : _GEN_2738; // @[i_cache.scala 91:40]
  wire  _GEN_3123 = unuse_way == 2'h2 ? _GEN_1202 : _GEN_2739; // @[i_cache.scala 91:40]
  wire  _GEN_3124 = unuse_way == 2'h2 ? _GEN_1203 : _GEN_2740; // @[i_cache.scala 91:40]
  wire  _GEN_3125 = unuse_way == 2'h2 ? _GEN_1204 : _GEN_2741; // @[i_cache.scala 91:40]
  wire  _GEN_3126 = unuse_way == 2'h2 ? _GEN_1205 : _GEN_2742; // @[i_cache.scala 91:40]
  wire  _GEN_3127 = unuse_way == 2'h2 ? _GEN_1206 : _GEN_2743; // @[i_cache.scala 91:40]
  wire  _GEN_3128 = unuse_way == 2'h2 ? _GEN_1207 : _GEN_2744; // @[i_cache.scala 91:40]
  wire  _GEN_3129 = unuse_way == 2'h2 ? _GEN_1208 : _GEN_2745; // @[i_cache.scala 91:40]
  wire  _GEN_3130 = unuse_way == 2'h2 ? _GEN_1209 : _GEN_2746; // @[i_cache.scala 91:40]
  wire  _GEN_3131 = unuse_way == 2'h2 ? _GEN_1210 : _GEN_2747; // @[i_cache.scala 91:40]
  wire  _GEN_3132 = unuse_way == 2'h2 ? _GEN_1211 : _GEN_2748; // @[i_cache.scala 91:40]
  wire  _GEN_3133 = unuse_way == 2'h2 ? _GEN_1212 : _GEN_2749; // @[i_cache.scala 91:40]
  wire  _GEN_3134 = unuse_way == 2'h2 ? _GEN_1213 : _GEN_2750; // @[i_cache.scala 91:40]
  wire  _GEN_3135 = unuse_way == 2'h2 ? _GEN_1214 : _GEN_2751; // @[i_cache.scala 91:40]
  wire  _GEN_3136 = unuse_way == 2'h2 ? _GEN_1215 : _GEN_2752; // @[i_cache.scala 91:40]
  wire  _GEN_3137 = unuse_way == 2'h2 ? _GEN_1216 : _GEN_2753; // @[i_cache.scala 91:40]
  wire  _GEN_3138 = unuse_way == 2'h2 ? _GEN_1217 : _GEN_2754; // @[i_cache.scala 91:40]
  wire  _GEN_3139 = unuse_way == 2'h2 ? _GEN_1218 : _GEN_2755; // @[i_cache.scala 91:40]
  wire  _GEN_3140 = unuse_way == 2'h2 ? _GEN_1219 : _GEN_2756; // @[i_cache.scala 91:40]
  wire  _GEN_3141 = unuse_way == 2'h2 ? _GEN_1220 : _GEN_2757; // @[i_cache.scala 91:40]
  wire  _GEN_3142 = unuse_way == 2'h2 ? _GEN_1221 : _GEN_2758; // @[i_cache.scala 91:40]
  wire  _GEN_3143 = unuse_way == 2'h2 ? _GEN_1222 : _GEN_2759; // @[i_cache.scala 91:40]
  wire  _GEN_3144 = unuse_way == 2'h2 ? _GEN_1223 : _GEN_2760; // @[i_cache.scala 91:40]
  wire  _GEN_3145 = unuse_way == 2'h2 ? _GEN_1224 : _GEN_2761; // @[i_cache.scala 91:40]
  wire  _GEN_3146 = unuse_way == 2'h2 ? _GEN_1225 : _GEN_2762; // @[i_cache.scala 91:40]
  wire  _GEN_3147 = unuse_way == 2'h2 ? _GEN_1226 : _GEN_2763; // @[i_cache.scala 91:40]
  wire  _GEN_3148 = unuse_way == 2'h2 ? _GEN_1227 : _GEN_2764; // @[i_cache.scala 91:40]
  wire  _GEN_3149 = unuse_way == 2'h2 ? _GEN_1228 : _GEN_2765; // @[i_cache.scala 91:40]
  wire  _GEN_3150 = unuse_way == 2'h2 ? _GEN_1229 : _GEN_2766; // @[i_cache.scala 91:40]
  wire  _GEN_3151 = unuse_way == 2'h2 ? _GEN_1230 : _GEN_2767; // @[i_cache.scala 91:40]
  wire  _GEN_3152 = unuse_way == 2'h2 ? _GEN_1231 : _GEN_2768; // @[i_cache.scala 91:40]
  wire  _GEN_3153 = unuse_way == 2'h2 ? _GEN_1232 : _GEN_2769; // @[i_cache.scala 91:40]
  wire  _GEN_3154 = unuse_way == 2'h2 ? _GEN_1233 : _GEN_2770; // @[i_cache.scala 91:40]
  wire  _GEN_3155 = unuse_way == 2'h2 ? _GEN_1234 : _GEN_2771; // @[i_cache.scala 91:40]
  wire  _GEN_3156 = unuse_way == 2'h2 ? _GEN_1235 : _GEN_2772; // @[i_cache.scala 91:40]
  wire  _GEN_3157 = unuse_way == 2'h2 ? _GEN_1236 : _GEN_2773; // @[i_cache.scala 91:40]
  wire  _GEN_3158 = unuse_way == 2'h2 ? _GEN_1237 : _GEN_2774; // @[i_cache.scala 91:40]
  wire  _GEN_3159 = unuse_way == 2'h2 ? _GEN_1238 : _GEN_2775; // @[i_cache.scala 91:40]
  wire  _GEN_3160 = unuse_way == 2'h2 ? _GEN_1239 : _GEN_2776; // @[i_cache.scala 91:40]
  wire  _GEN_3161 = unuse_way == 2'h2 ? _GEN_1240 : _GEN_2777; // @[i_cache.scala 91:40]
  wire  _GEN_3162 = unuse_way == 2'h2 ? _GEN_1241 : _GEN_2778; // @[i_cache.scala 91:40]
  wire  _GEN_3163 = unuse_way == 2'h2 ? _GEN_1242 : _GEN_2779; // @[i_cache.scala 91:40]
  wire  _GEN_3164 = unuse_way == 2'h2 ? _GEN_1243 : _GEN_2780; // @[i_cache.scala 91:40]
  wire  _GEN_3165 = unuse_way == 2'h2 ? _GEN_1244 : _GEN_2781; // @[i_cache.scala 91:40]
  wire  _GEN_3166 = unuse_way == 2'h2 ? _GEN_1245 : _GEN_2782; // @[i_cache.scala 91:40]
  wire  _GEN_3167 = unuse_way == 2'h2 ? _GEN_1246 : _GEN_2783; // @[i_cache.scala 91:40]
  wire  _GEN_3168 = unuse_way == 2'h2 ? _GEN_1247 : _GEN_2784; // @[i_cache.scala 91:40]
  wire  _GEN_3169 = unuse_way == 2'h2 ? _GEN_1248 : _GEN_2785; // @[i_cache.scala 91:40]
  wire  _GEN_3170 = unuse_way == 2'h2 ? _GEN_1249 : _GEN_2786; // @[i_cache.scala 91:40]
  wire  _GEN_3171 = unuse_way == 2'h2 ? _GEN_1250 : _GEN_2787; // @[i_cache.scala 91:40]
  wire  _GEN_3172 = unuse_way == 2'h2 ? _GEN_1251 : _GEN_2788; // @[i_cache.scala 91:40]
  wire  _GEN_3173 = unuse_way == 2'h2 ? _GEN_1252 : _GEN_2789; // @[i_cache.scala 91:40]
  wire  _GEN_3174 = unuse_way == 2'h2 ? _GEN_1253 : _GEN_2790; // @[i_cache.scala 91:40]
  wire  _GEN_3175 = unuse_way == 2'h2 ? _GEN_1254 : _GEN_2791; // @[i_cache.scala 91:40]
  wire  _GEN_3176 = unuse_way == 2'h2 ? _GEN_1255 : _GEN_2792; // @[i_cache.scala 91:40]
  wire  _GEN_3177 = unuse_way == 2'h2 ? _GEN_1256 : _GEN_2793; // @[i_cache.scala 91:40]
  wire  _GEN_3178 = unuse_way == 2'h2 ? _GEN_1257 : _GEN_2794; // @[i_cache.scala 91:40]
  wire  _GEN_3179 = unuse_way == 2'h2 ? _GEN_1258 : _GEN_2795; // @[i_cache.scala 91:40]
  wire  _GEN_3180 = unuse_way == 2'h2 ? _GEN_1259 : _GEN_2796; // @[i_cache.scala 91:40]
  wire  _GEN_3181 = unuse_way == 2'h2 ? _GEN_1260 : _GEN_2797; // @[i_cache.scala 91:40]
  wire  _GEN_3182 = unuse_way == 2'h2 ? _GEN_1261 : _GEN_2798; // @[i_cache.scala 91:40]
  wire  _GEN_3183 = unuse_way == 2'h2 ? _GEN_1262 : _GEN_2799; // @[i_cache.scala 91:40]
  wire  _GEN_3184 = unuse_way == 2'h2 ? _GEN_1263 : _GEN_2800; // @[i_cache.scala 91:40]
  wire  _GEN_3185 = unuse_way == 2'h2 ? _GEN_1264 : _GEN_2801; // @[i_cache.scala 91:40]
  wire  _GEN_3186 = unuse_way == 2'h2 ? _GEN_1265 : _GEN_2802; // @[i_cache.scala 91:40]
  wire  _GEN_3187 = unuse_way == 2'h2 ? _GEN_1266 : _GEN_2803; // @[i_cache.scala 91:40]
  wire  _GEN_3188 = unuse_way == 2'h2 ? _GEN_1267 : _GEN_2804; // @[i_cache.scala 91:40]
  wire  _GEN_3189 = unuse_way == 2'h2 ? _GEN_1268 : _GEN_2805; // @[i_cache.scala 91:40]
  wire  _GEN_3190 = unuse_way == 2'h2 ? _GEN_1269 : _GEN_2806; // @[i_cache.scala 91:40]
  wire  _GEN_3191 = unuse_way == 2'h2 ? _GEN_1270 : _GEN_2807; // @[i_cache.scala 91:40]
  wire  _GEN_3192 = unuse_way == 2'h2 ? _GEN_1271 : _GEN_2808; // @[i_cache.scala 91:40]
  wire  _GEN_3193 = unuse_way == 2'h2 ? _GEN_1272 : _GEN_2809; // @[i_cache.scala 91:40]
  wire  _GEN_3194 = unuse_way == 2'h2 ? _GEN_1273 : _GEN_2810; // @[i_cache.scala 91:40]
  wire  _GEN_3195 = unuse_way == 2'h2 ? _GEN_1274 : _GEN_2811; // @[i_cache.scala 91:40]
  wire  _GEN_3196 = unuse_way == 2'h2 ? _GEN_1275 : _GEN_2812; // @[i_cache.scala 91:40]
  wire  _GEN_3197 = unuse_way == 2'h2 ? _GEN_1276 : _GEN_2813; // @[i_cache.scala 91:40]
  wire  _GEN_3198 = unuse_way == 2'h2 ? _GEN_1277 : _GEN_2814; // @[i_cache.scala 91:40]
  wire  _GEN_3199 = unuse_way == 2'h2 ? _GEN_1278 : _GEN_2815; // @[i_cache.scala 91:40]
  wire  _GEN_3200 = unuse_way == 2'h2 ? _GEN_1279 : _GEN_2816; // @[i_cache.scala 91:40]
  wire  _GEN_3201 = unuse_way == 2'h2 ? _GEN_1280 : _GEN_2817; // @[i_cache.scala 91:40]
  wire  _GEN_3202 = unuse_way == 2'h2 ? _GEN_1281 : _GEN_2818; // @[i_cache.scala 91:40]
  wire  _GEN_3203 = unuse_way == 2'h2 ? _GEN_1282 : _GEN_2819; // @[i_cache.scala 91:40]
  wire  _GEN_3204 = unuse_way == 2'h2 ? _GEN_1283 : _GEN_2820; // @[i_cache.scala 91:40]
  wire  _GEN_3205 = unuse_way == 2'h2 ? _GEN_1284 : _GEN_2821; // @[i_cache.scala 91:40]
  wire  _GEN_3206 = unuse_way == 2'h2 ? _GEN_1285 : _GEN_2822; // @[i_cache.scala 91:40]
  wire  _GEN_3207 = unuse_way == 2'h2 ? _GEN_1286 : _GEN_2823; // @[i_cache.scala 91:40]
  wire  _GEN_3208 = unuse_way == 2'h2 ? _GEN_1287 : _GEN_2824; // @[i_cache.scala 91:40]
  wire  _GEN_3209 = unuse_way == 2'h2 ? _GEN_1288 : _GEN_2825; // @[i_cache.scala 91:40]
  wire  _GEN_3210 = unuse_way == 2'h2 ? _GEN_1289 : _GEN_2826; // @[i_cache.scala 91:40]
  wire  _GEN_3211 = unuse_way == 2'h2 ? 1'h0 : _T_14; // @[i_cache.scala 91:40 95:23]
  wire [63:0] _GEN_3212 = unuse_way == 2'h2 ? ram_0_0 : _GEN_2058; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3213 = unuse_way == 2'h2 ? ram_0_1 : _GEN_2059; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3214 = unuse_way == 2'h2 ? ram_0_2 : _GEN_2060; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3215 = unuse_way == 2'h2 ? ram_0_3 : _GEN_2061; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3216 = unuse_way == 2'h2 ? ram_0_4 : _GEN_2062; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3217 = unuse_way == 2'h2 ? ram_0_5 : _GEN_2063; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3218 = unuse_way == 2'h2 ? ram_0_6 : _GEN_2064; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3219 = unuse_way == 2'h2 ? ram_0_7 : _GEN_2065; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3220 = unuse_way == 2'h2 ? ram_0_8 : _GEN_2066; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3221 = unuse_way == 2'h2 ? ram_0_9 : _GEN_2067; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3222 = unuse_way == 2'h2 ? ram_0_10 : _GEN_2068; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3223 = unuse_way == 2'h2 ? ram_0_11 : _GEN_2069; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3224 = unuse_way == 2'h2 ? ram_0_12 : _GEN_2070; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3225 = unuse_way == 2'h2 ? ram_0_13 : _GEN_2071; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3226 = unuse_way == 2'h2 ? ram_0_14 : _GEN_2072; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3227 = unuse_way == 2'h2 ? ram_0_15 : _GEN_2073; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3228 = unuse_way == 2'h2 ? ram_0_16 : _GEN_2074; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3229 = unuse_way == 2'h2 ? ram_0_17 : _GEN_2075; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3230 = unuse_way == 2'h2 ? ram_0_18 : _GEN_2076; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3231 = unuse_way == 2'h2 ? ram_0_19 : _GEN_2077; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3232 = unuse_way == 2'h2 ? ram_0_20 : _GEN_2078; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3233 = unuse_way == 2'h2 ? ram_0_21 : _GEN_2079; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3234 = unuse_way == 2'h2 ? ram_0_22 : _GEN_2080; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3235 = unuse_way == 2'h2 ? ram_0_23 : _GEN_2081; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3236 = unuse_way == 2'h2 ? ram_0_24 : _GEN_2082; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3237 = unuse_way == 2'h2 ? ram_0_25 : _GEN_2083; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3238 = unuse_way == 2'h2 ? ram_0_26 : _GEN_2084; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3239 = unuse_way == 2'h2 ? ram_0_27 : _GEN_2085; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3240 = unuse_way == 2'h2 ? ram_0_28 : _GEN_2086; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3241 = unuse_way == 2'h2 ? ram_0_29 : _GEN_2087; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3242 = unuse_way == 2'h2 ? ram_0_30 : _GEN_2088; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3243 = unuse_way == 2'h2 ? ram_0_31 : _GEN_2089; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3244 = unuse_way == 2'h2 ? ram_0_32 : _GEN_2090; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3245 = unuse_way == 2'h2 ? ram_0_33 : _GEN_2091; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3246 = unuse_way == 2'h2 ? ram_0_34 : _GEN_2092; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3247 = unuse_way == 2'h2 ? ram_0_35 : _GEN_2093; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3248 = unuse_way == 2'h2 ? ram_0_36 : _GEN_2094; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3249 = unuse_way == 2'h2 ? ram_0_37 : _GEN_2095; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3250 = unuse_way == 2'h2 ? ram_0_38 : _GEN_2096; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3251 = unuse_way == 2'h2 ? ram_0_39 : _GEN_2097; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3252 = unuse_way == 2'h2 ? ram_0_40 : _GEN_2098; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3253 = unuse_way == 2'h2 ? ram_0_41 : _GEN_2099; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3254 = unuse_way == 2'h2 ? ram_0_42 : _GEN_2100; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3255 = unuse_way == 2'h2 ? ram_0_43 : _GEN_2101; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3256 = unuse_way == 2'h2 ? ram_0_44 : _GEN_2102; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3257 = unuse_way == 2'h2 ? ram_0_45 : _GEN_2103; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3258 = unuse_way == 2'h2 ? ram_0_46 : _GEN_2104; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3259 = unuse_way == 2'h2 ? ram_0_47 : _GEN_2105; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3260 = unuse_way == 2'h2 ? ram_0_48 : _GEN_2106; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3261 = unuse_way == 2'h2 ? ram_0_49 : _GEN_2107; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3262 = unuse_way == 2'h2 ? ram_0_50 : _GEN_2108; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3263 = unuse_way == 2'h2 ? ram_0_51 : _GEN_2109; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3264 = unuse_way == 2'h2 ? ram_0_52 : _GEN_2110; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3265 = unuse_way == 2'h2 ? ram_0_53 : _GEN_2111; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3266 = unuse_way == 2'h2 ? ram_0_54 : _GEN_2112; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3267 = unuse_way == 2'h2 ? ram_0_55 : _GEN_2113; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3268 = unuse_way == 2'h2 ? ram_0_56 : _GEN_2114; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3269 = unuse_way == 2'h2 ? ram_0_57 : _GEN_2115; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3270 = unuse_way == 2'h2 ? ram_0_58 : _GEN_2116; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3271 = unuse_way == 2'h2 ? ram_0_59 : _GEN_2117; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3272 = unuse_way == 2'h2 ? ram_0_60 : _GEN_2118; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3273 = unuse_way == 2'h2 ? ram_0_61 : _GEN_2119; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3274 = unuse_way == 2'h2 ? ram_0_62 : _GEN_2120; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3275 = unuse_way == 2'h2 ? ram_0_63 : _GEN_2121; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3276 = unuse_way == 2'h2 ? ram_0_64 : _GEN_2122; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3277 = unuse_way == 2'h2 ? ram_0_65 : _GEN_2123; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3278 = unuse_way == 2'h2 ? ram_0_66 : _GEN_2124; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3279 = unuse_way == 2'h2 ? ram_0_67 : _GEN_2125; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3280 = unuse_way == 2'h2 ? ram_0_68 : _GEN_2126; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3281 = unuse_way == 2'h2 ? ram_0_69 : _GEN_2127; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3282 = unuse_way == 2'h2 ? ram_0_70 : _GEN_2128; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3283 = unuse_way == 2'h2 ? ram_0_71 : _GEN_2129; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3284 = unuse_way == 2'h2 ? ram_0_72 : _GEN_2130; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3285 = unuse_way == 2'h2 ? ram_0_73 : _GEN_2131; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3286 = unuse_way == 2'h2 ? ram_0_74 : _GEN_2132; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3287 = unuse_way == 2'h2 ? ram_0_75 : _GEN_2133; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3288 = unuse_way == 2'h2 ? ram_0_76 : _GEN_2134; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3289 = unuse_way == 2'h2 ? ram_0_77 : _GEN_2135; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3290 = unuse_way == 2'h2 ? ram_0_78 : _GEN_2136; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3291 = unuse_way == 2'h2 ? ram_0_79 : _GEN_2137; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3292 = unuse_way == 2'h2 ? ram_0_80 : _GEN_2138; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3293 = unuse_way == 2'h2 ? ram_0_81 : _GEN_2139; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3294 = unuse_way == 2'h2 ? ram_0_82 : _GEN_2140; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3295 = unuse_way == 2'h2 ? ram_0_83 : _GEN_2141; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3296 = unuse_way == 2'h2 ? ram_0_84 : _GEN_2142; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3297 = unuse_way == 2'h2 ? ram_0_85 : _GEN_2143; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3298 = unuse_way == 2'h2 ? ram_0_86 : _GEN_2144; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3299 = unuse_way == 2'h2 ? ram_0_87 : _GEN_2145; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3300 = unuse_way == 2'h2 ? ram_0_88 : _GEN_2146; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3301 = unuse_way == 2'h2 ? ram_0_89 : _GEN_2147; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3302 = unuse_way == 2'h2 ? ram_0_90 : _GEN_2148; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3303 = unuse_way == 2'h2 ? ram_0_91 : _GEN_2149; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3304 = unuse_way == 2'h2 ? ram_0_92 : _GEN_2150; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3305 = unuse_way == 2'h2 ? ram_0_93 : _GEN_2151; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3306 = unuse_way == 2'h2 ? ram_0_94 : _GEN_2152; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3307 = unuse_way == 2'h2 ? ram_0_95 : _GEN_2153; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3308 = unuse_way == 2'h2 ? ram_0_96 : _GEN_2154; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3309 = unuse_way == 2'h2 ? ram_0_97 : _GEN_2155; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3310 = unuse_way == 2'h2 ? ram_0_98 : _GEN_2156; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3311 = unuse_way == 2'h2 ? ram_0_99 : _GEN_2157; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3312 = unuse_way == 2'h2 ? ram_0_100 : _GEN_2158; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3313 = unuse_way == 2'h2 ? ram_0_101 : _GEN_2159; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3314 = unuse_way == 2'h2 ? ram_0_102 : _GEN_2160; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3315 = unuse_way == 2'h2 ? ram_0_103 : _GEN_2161; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3316 = unuse_way == 2'h2 ? ram_0_104 : _GEN_2162; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3317 = unuse_way == 2'h2 ? ram_0_105 : _GEN_2163; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3318 = unuse_way == 2'h2 ? ram_0_106 : _GEN_2164; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3319 = unuse_way == 2'h2 ? ram_0_107 : _GEN_2165; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3320 = unuse_way == 2'h2 ? ram_0_108 : _GEN_2166; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3321 = unuse_way == 2'h2 ? ram_0_109 : _GEN_2167; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3322 = unuse_way == 2'h2 ? ram_0_110 : _GEN_2168; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3323 = unuse_way == 2'h2 ? ram_0_111 : _GEN_2169; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3324 = unuse_way == 2'h2 ? ram_0_112 : _GEN_2170; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3325 = unuse_way == 2'h2 ? ram_0_113 : _GEN_2171; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3326 = unuse_way == 2'h2 ? ram_0_114 : _GEN_2172; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3327 = unuse_way == 2'h2 ? ram_0_115 : _GEN_2173; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3328 = unuse_way == 2'h2 ? ram_0_116 : _GEN_2174; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3329 = unuse_way == 2'h2 ? ram_0_117 : _GEN_2175; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3330 = unuse_way == 2'h2 ? ram_0_118 : _GEN_2176; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3331 = unuse_way == 2'h2 ? ram_0_119 : _GEN_2177; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3332 = unuse_way == 2'h2 ? ram_0_120 : _GEN_2178; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3333 = unuse_way == 2'h2 ? ram_0_121 : _GEN_2179; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3334 = unuse_way == 2'h2 ? ram_0_122 : _GEN_2180; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3335 = unuse_way == 2'h2 ? ram_0_123 : _GEN_2181; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3336 = unuse_way == 2'h2 ? ram_0_124 : _GEN_2182; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3337 = unuse_way == 2'h2 ? ram_0_125 : _GEN_2183; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3338 = unuse_way == 2'h2 ? ram_0_126 : _GEN_2184; // @[i_cache.scala 17:24 91:40]
  wire [63:0] _GEN_3339 = unuse_way == 2'h2 ? ram_0_127 : _GEN_2185; // @[i_cache.scala 17:24 91:40]
  wire [31:0] _GEN_3340 = unuse_way == 2'h2 ? tag_0_0 : _GEN_2186; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3341 = unuse_way == 2'h2 ? tag_0_1 : _GEN_2187; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3342 = unuse_way == 2'h2 ? tag_0_2 : _GEN_2188; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3343 = unuse_way == 2'h2 ? tag_0_3 : _GEN_2189; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3344 = unuse_way == 2'h2 ? tag_0_4 : _GEN_2190; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3345 = unuse_way == 2'h2 ? tag_0_5 : _GEN_2191; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3346 = unuse_way == 2'h2 ? tag_0_6 : _GEN_2192; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3347 = unuse_way == 2'h2 ? tag_0_7 : _GEN_2193; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3348 = unuse_way == 2'h2 ? tag_0_8 : _GEN_2194; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3349 = unuse_way == 2'h2 ? tag_0_9 : _GEN_2195; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3350 = unuse_way == 2'h2 ? tag_0_10 : _GEN_2196; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3351 = unuse_way == 2'h2 ? tag_0_11 : _GEN_2197; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3352 = unuse_way == 2'h2 ? tag_0_12 : _GEN_2198; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3353 = unuse_way == 2'h2 ? tag_0_13 : _GEN_2199; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3354 = unuse_way == 2'h2 ? tag_0_14 : _GEN_2200; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3355 = unuse_way == 2'h2 ? tag_0_15 : _GEN_2201; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3356 = unuse_way == 2'h2 ? tag_0_16 : _GEN_2202; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3357 = unuse_way == 2'h2 ? tag_0_17 : _GEN_2203; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3358 = unuse_way == 2'h2 ? tag_0_18 : _GEN_2204; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3359 = unuse_way == 2'h2 ? tag_0_19 : _GEN_2205; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3360 = unuse_way == 2'h2 ? tag_0_20 : _GEN_2206; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3361 = unuse_way == 2'h2 ? tag_0_21 : _GEN_2207; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3362 = unuse_way == 2'h2 ? tag_0_22 : _GEN_2208; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3363 = unuse_way == 2'h2 ? tag_0_23 : _GEN_2209; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3364 = unuse_way == 2'h2 ? tag_0_24 : _GEN_2210; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3365 = unuse_way == 2'h2 ? tag_0_25 : _GEN_2211; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3366 = unuse_way == 2'h2 ? tag_0_26 : _GEN_2212; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3367 = unuse_way == 2'h2 ? tag_0_27 : _GEN_2213; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3368 = unuse_way == 2'h2 ? tag_0_28 : _GEN_2214; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3369 = unuse_way == 2'h2 ? tag_0_29 : _GEN_2215; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3370 = unuse_way == 2'h2 ? tag_0_30 : _GEN_2216; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3371 = unuse_way == 2'h2 ? tag_0_31 : _GEN_2217; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3372 = unuse_way == 2'h2 ? tag_0_32 : _GEN_2218; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3373 = unuse_way == 2'h2 ? tag_0_33 : _GEN_2219; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3374 = unuse_way == 2'h2 ? tag_0_34 : _GEN_2220; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3375 = unuse_way == 2'h2 ? tag_0_35 : _GEN_2221; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3376 = unuse_way == 2'h2 ? tag_0_36 : _GEN_2222; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3377 = unuse_way == 2'h2 ? tag_0_37 : _GEN_2223; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3378 = unuse_way == 2'h2 ? tag_0_38 : _GEN_2224; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3379 = unuse_way == 2'h2 ? tag_0_39 : _GEN_2225; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3380 = unuse_way == 2'h2 ? tag_0_40 : _GEN_2226; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3381 = unuse_way == 2'h2 ? tag_0_41 : _GEN_2227; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3382 = unuse_way == 2'h2 ? tag_0_42 : _GEN_2228; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3383 = unuse_way == 2'h2 ? tag_0_43 : _GEN_2229; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3384 = unuse_way == 2'h2 ? tag_0_44 : _GEN_2230; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3385 = unuse_way == 2'h2 ? tag_0_45 : _GEN_2231; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3386 = unuse_way == 2'h2 ? tag_0_46 : _GEN_2232; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3387 = unuse_way == 2'h2 ? tag_0_47 : _GEN_2233; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3388 = unuse_way == 2'h2 ? tag_0_48 : _GEN_2234; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3389 = unuse_way == 2'h2 ? tag_0_49 : _GEN_2235; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3390 = unuse_way == 2'h2 ? tag_0_50 : _GEN_2236; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3391 = unuse_way == 2'h2 ? tag_0_51 : _GEN_2237; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3392 = unuse_way == 2'h2 ? tag_0_52 : _GEN_2238; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3393 = unuse_way == 2'h2 ? tag_0_53 : _GEN_2239; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3394 = unuse_way == 2'h2 ? tag_0_54 : _GEN_2240; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3395 = unuse_way == 2'h2 ? tag_0_55 : _GEN_2241; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3396 = unuse_way == 2'h2 ? tag_0_56 : _GEN_2242; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3397 = unuse_way == 2'h2 ? tag_0_57 : _GEN_2243; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3398 = unuse_way == 2'h2 ? tag_0_58 : _GEN_2244; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3399 = unuse_way == 2'h2 ? tag_0_59 : _GEN_2245; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3400 = unuse_way == 2'h2 ? tag_0_60 : _GEN_2246; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3401 = unuse_way == 2'h2 ? tag_0_61 : _GEN_2247; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3402 = unuse_way == 2'h2 ? tag_0_62 : _GEN_2248; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3403 = unuse_way == 2'h2 ? tag_0_63 : _GEN_2249; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3404 = unuse_way == 2'h2 ? tag_0_64 : _GEN_2250; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3405 = unuse_way == 2'h2 ? tag_0_65 : _GEN_2251; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3406 = unuse_way == 2'h2 ? tag_0_66 : _GEN_2252; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3407 = unuse_way == 2'h2 ? tag_0_67 : _GEN_2253; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3408 = unuse_way == 2'h2 ? tag_0_68 : _GEN_2254; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3409 = unuse_way == 2'h2 ? tag_0_69 : _GEN_2255; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3410 = unuse_way == 2'h2 ? tag_0_70 : _GEN_2256; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3411 = unuse_way == 2'h2 ? tag_0_71 : _GEN_2257; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3412 = unuse_way == 2'h2 ? tag_0_72 : _GEN_2258; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3413 = unuse_way == 2'h2 ? tag_0_73 : _GEN_2259; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3414 = unuse_way == 2'h2 ? tag_0_74 : _GEN_2260; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3415 = unuse_way == 2'h2 ? tag_0_75 : _GEN_2261; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3416 = unuse_way == 2'h2 ? tag_0_76 : _GEN_2262; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3417 = unuse_way == 2'h2 ? tag_0_77 : _GEN_2263; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3418 = unuse_way == 2'h2 ? tag_0_78 : _GEN_2264; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3419 = unuse_way == 2'h2 ? tag_0_79 : _GEN_2265; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3420 = unuse_way == 2'h2 ? tag_0_80 : _GEN_2266; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3421 = unuse_way == 2'h2 ? tag_0_81 : _GEN_2267; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3422 = unuse_way == 2'h2 ? tag_0_82 : _GEN_2268; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3423 = unuse_way == 2'h2 ? tag_0_83 : _GEN_2269; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3424 = unuse_way == 2'h2 ? tag_0_84 : _GEN_2270; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3425 = unuse_way == 2'h2 ? tag_0_85 : _GEN_2271; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3426 = unuse_way == 2'h2 ? tag_0_86 : _GEN_2272; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3427 = unuse_way == 2'h2 ? tag_0_87 : _GEN_2273; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3428 = unuse_way == 2'h2 ? tag_0_88 : _GEN_2274; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3429 = unuse_way == 2'h2 ? tag_0_89 : _GEN_2275; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3430 = unuse_way == 2'h2 ? tag_0_90 : _GEN_2276; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3431 = unuse_way == 2'h2 ? tag_0_91 : _GEN_2277; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3432 = unuse_way == 2'h2 ? tag_0_92 : _GEN_2278; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3433 = unuse_way == 2'h2 ? tag_0_93 : _GEN_2279; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3434 = unuse_way == 2'h2 ? tag_0_94 : _GEN_2280; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3435 = unuse_way == 2'h2 ? tag_0_95 : _GEN_2281; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3436 = unuse_way == 2'h2 ? tag_0_96 : _GEN_2282; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3437 = unuse_way == 2'h2 ? tag_0_97 : _GEN_2283; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3438 = unuse_way == 2'h2 ? tag_0_98 : _GEN_2284; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3439 = unuse_way == 2'h2 ? tag_0_99 : _GEN_2285; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3440 = unuse_way == 2'h2 ? tag_0_100 : _GEN_2286; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3441 = unuse_way == 2'h2 ? tag_0_101 : _GEN_2287; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3442 = unuse_way == 2'h2 ? tag_0_102 : _GEN_2288; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3443 = unuse_way == 2'h2 ? tag_0_103 : _GEN_2289; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3444 = unuse_way == 2'h2 ? tag_0_104 : _GEN_2290; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3445 = unuse_way == 2'h2 ? tag_0_105 : _GEN_2291; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3446 = unuse_way == 2'h2 ? tag_0_106 : _GEN_2292; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3447 = unuse_way == 2'h2 ? tag_0_107 : _GEN_2293; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3448 = unuse_way == 2'h2 ? tag_0_108 : _GEN_2294; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3449 = unuse_way == 2'h2 ? tag_0_109 : _GEN_2295; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3450 = unuse_way == 2'h2 ? tag_0_110 : _GEN_2296; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3451 = unuse_way == 2'h2 ? tag_0_111 : _GEN_2297; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3452 = unuse_way == 2'h2 ? tag_0_112 : _GEN_2298; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3453 = unuse_way == 2'h2 ? tag_0_113 : _GEN_2299; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3454 = unuse_way == 2'h2 ? tag_0_114 : _GEN_2300; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3455 = unuse_way == 2'h2 ? tag_0_115 : _GEN_2301; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3456 = unuse_way == 2'h2 ? tag_0_116 : _GEN_2302; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3457 = unuse_way == 2'h2 ? tag_0_117 : _GEN_2303; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3458 = unuse_way == 2'h2 ? tag_0_118 : _GEN_2304; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3459 = unuse_way == 2'h2 ? tag_0_119 : _GEN_2305; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3460 = unuse_way == 2'h2 ? tag_0_120 : _GEN_2306; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3461 = unuse_way == 2'h2 ? tag_0_121 : _GEN_2307; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3462 = unuse_way == 2'h2 ? tag_0_122 : _GEN_2308; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3463 = unuse_way == 2'h2 ? tag_0_123 : _GEN_2309; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3464 = unuse_way == 2'h2 ? tag_0_124 : _GEN_2310; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3465 = unuse_way == 2'h2 ? tag_0_125 : _GEN_2311; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3466 = unuse_way == 2'h2 ? tag_0_126 : _GEN_2312; // @[i_cache.scala 19:24 91:40]
  wire [31:0] _GEN_3467 = unuse_way == 2'h2 ? tag_0_127 : _GEN_2313; // @[i_cache.scala 19:24 91:40]
  wire  _GEN_3468 = unuse_way == 2'h2 ? valid_0_0 : _GEN_2314; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3469 = unuse_way == 2'h2 ? valid_0_1 : _GEN_2315; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3470 = unuse_way == 2'h2 ? valid_0_2 : _GEN_2316; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3471 = unuse_way == 2'h2 ? valid_0_3 : _GEN_2317; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3472 = unuse_way == 2'h2 ? valid_0_4 : _GEN_2318; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3473 = unuse_way == 2'h2 ? valid_0_5 : _GEN_2319; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3474 = unuse_way == 2'h2 ? valid_0_6 : _GEN_2320; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3475 = unuse_way == 2'h2 ? valid_0_7 : _GEN_2321; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3476 = unuse_way == 2'h2 ? valid_0_8 : _GEN_2322; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3477 = unuse_way == 2'h2 ? valid_0_9 : _GEN_2323; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3478 = unuse_way == 2'h2 ? valid_0_10 : _GEN_2324; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3479 = unuse_way == 2'h2 ? valid_0_11 : _GEN_2325; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3480 = unuse_way == 2'h2 ? valid_0_12 : _GEN_2326; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3481 = unuse_way == 2'h2 ? valid_0_13 : _GEN_2327; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3482 = unuse_way == 2'h2 ? valid_0_14 : _GEN_2328; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3483 = unuse_way == 2'h2 ? valid_0_15 : _GEN_2329; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3484 = unuse_way == 2'h2 ? valid_0_16 : _GEN_2330; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3485 = unuse_way == 2'h2 ? valid_0_17 : _GEN_2331; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3486 = unuse_way == 2'h2 ? valid_0_18 : _GEN_2332; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3487 = unuse_way == 2'h2 ? valid_0_19 : _GEN_2333; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3488 = unuse_way == 2'h2 ? valid_0_20 : _GEN_2334; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3489 = unuse_way == 2'h2 ? valid_0_21 : _GEN_2335; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3490 = unuse_way == 2'h2 ? valid_0_22 : _GEN_2336; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3491 = unuse_way == 2'h2 ? valid_0_23 : _GEN_2337; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3492 = unuse_way == 2'h2 ? valid_0_24 : _GEN_2338; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3493 = unuse_way == 2'h2 ? valid_0_25 : _GEN_2339; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3494 = unuse_way == 2'h2 ? valid_0_26 : _GEN_2340; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3495 = unuse_way == 2'h2 ? valid_0_27 : _GEN_2341; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3496 = unuse_way == 2'h2 ? valid_0_28 : _GEN_2342; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3497 = unuse_way == 2'h2 ? valid_0_29 : _GEN_2343; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3498 = unuse_way == 2'h2 ? valid_0_30 : _GEN_2344; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3499 = unuse_way == 2'h2 ? valid_0_31 : _GEN_2345; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3500 = unuse_way == 2'h2 ? valid_0_32 : _GEN_2346; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3501 = unuse_way == 2'h2 ? valid_0_33 : _GEN_2347; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3502 = unuse_way == 2'h2 ? valid_0_34 : _GEN_2348; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3503 = unuse_way == 2'h2 ? valid_0_35 : _GEN_2349; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3504 = unuse_way == 2'h2 ? valid_0_36 : _GEN_2350; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3505 = unuse_way == 2'h2 ? valid_0_37 : _GEN_2351; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3506 = unuse_way == 2'h2 ? valid_0_38 : _GEN_2352; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3507 = unuse_way == 2'h2 ? valid_0_39 : _GEN_2353; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3508 = unuse_way == 2'h2 ? valid_0_40 : _GEN_2354; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3509 = unuse_way == 2'h2 ? valid_0_41 : _GEN_2355; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3510 = unuse_way == 2'h2 ? valid_0_42 : _GEN_2356; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3511 = unuse_way == 2'h2 ? valid_0_43 : _GEN_2357; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3512 = unuse_way == 2'h2 ? valid_0_44 : _GEN_2358; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3513 = unuse_way == 2'h2 ? valid_0_45 : _GEN_2359; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3514 = unuse_way == 2'h2 ? valid_0_46 : _GEN_2360; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3515 = unuse_way == 2'h2 ? valid_0_47 : _GEN_2361; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3516 = unuse_way == 2'h2 ? valid_0_48 : _GEN_2362; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3517 = unuse_way == 2'h2 ? valid_0_49 : _GEN_2363; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3518 = unuse_way == 2'h2 ? valid_0_50 : _GEN_2364; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3519 = unuse_way == 2'h2 ? valid_0_51 : _GEN_2365; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3520 = unuse_way == 2'h2 ? valid_0_52 : _GEN_2366; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3521 = unuse_way == 2'h2 ? valid_0_53 : _GEN_2367; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3522 = unuse_way == 2'h2 ? valid_0_54 : _GEN_2368; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3523 = unuse_way == 2'h2 ? valid_0_55 : _GEN_2369; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3524 = unuse_way == 2'h2 ? valid_0_56 : _GEN_2370; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3525 = unuse_way == 2'h2 ? valid_0_57 : _GEN_2371; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3526 = unuse_way == 2'h2 ? valid_0_58 : _GEN_2372; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3527 = unuse_way == 2'h2 ? valid_0_59 : _GEN_2373; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3528 = unuse_way == 2'h2 ? valid_0_60 : _GEN_2374; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3529 = unuse_way == 2'h2 ? valid_0_61 : _GEN_2375; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3530 = unuse_way == 2'h2 ? valid_0_62 : _GEN_2376; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3531 = unuse_way == 2'h2 ? valid_0_63 : _GEN_2377; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3532 = unuse_way == 2'h2 ? valid_0_64 : _GEN_2378; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3533 = unuse_way == 2'h2 ? valid_0_65 : _GEN_2379; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3534 = unuse_way == 2'h2 ? valid_0_66 : _GEN_2380; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3535 = unuse_way == 2'h2 ? valid_0_67 : _GEN_2381; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3536 = unuse_way == 2'h2 ? valid_0_68 : _GEN_2382; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3537 = unuse_way == 2'h2 ? valid_0_69 : _GEN_2383; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3538 = unuse_way == 2'h2 ? valid_0_70 : _GEN_2384; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3539 = unuse_way == 2'h2 ? valid_0_71 : _GEN_2385; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3540 = unuse_way == 2'h2 ? valid_0_72 : _GEN_2386; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3541 = unuse_way == 2'h2 ? valid_0_73 : _GEN_2387; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3542 = unuse_way == 2'h2 ? valid_0_74 : _GEN_2388; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3543 = unuse_way == 2'h2 ? valid_0_75 : _GEN_2389; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3544 = unuse_way == 2'h2 ? valid_0_76 : _GEN_2390; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3545 = unuse_way == 2'h2 ? valid_0_77 : _GEN_2391; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3546 = unuse_way == 2'h2 ? valid_0_78 : _GEN_2392; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3547 = unuse_way == 2'h2 ? valid_0_79 : _GEN_2393; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3548 = unuse_way == 2'h2 ? valid_0_80 : _GEN_2394; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3549 = unuse_way == 2'h2 ? valid_0_81 : _GEN_2395; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3550 = unuse_way == 2'h2 ? valid_0_82 : _GEN_2396; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3551 = unuse_way == 2'h2 ? valid_0_83 : _GEN_2397; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3552 = unuse_way == 2'h2 ? valid_0_84 : _GEN_2398; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3553 = unuse_way == 2'h2 ? valid_0_85 : _GEN_2399; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3554 = unuse_way == 2'h2 ? valid_0_86 : _GEN_2400; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3555 = unuse_way == 2'h2 ? valid_0_87 : _GEN_2401; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3556 = unuse_way == 2'h2 ? valid_0_88 : _GEN_2402; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3557 = unuse_way == 2'h2 ? valid_0_89 : _GEN_2403; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3558 = unuse_way == 2'h2 ? valid_0_90 : _GEN_2404; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3559 = unuse_way == 2'h2 ? valid_0_91 : _GEN_2405; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3560 = unuse_way == 2'h2 ? valid_0_92 : _GEN_2406; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3561 = unuse_way == 2'h2 ? valid_0_93 : _GEN_2407; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3562 = unuse_way == 2'h2 ? valid_0_94 : _GEN_2408; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3563 = unuse_way == 2'h2 ? valid_0_95 : _GEN_2409; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3564 = unuse_way == 2'h2 ? valid_0_96 : _GEN_2410; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3565 = unuse_way == 2'h2 ? valid_0_97 : _GEN_2411; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3566 = unuse_way == 2'h2 ? valid_0_98 : _GEN_2412; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3567 = unuse_way == 2'h2 ? valid_0_99 : _GEN_2413; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3568 = unuse_way == 2'h2 ? valid_0_100 : _GEN_2414; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3569 = unuse_way == 2'h2 ? valid_0_101 : _GEN_2415; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3570 = unuse_way == 2'h2 ? valid_0_102 : _GEN_2416; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3571 = unuse_way == 2'h2 ? valid_0_103 : _GEN_2417; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3572 = unuse_way == 2'h2 ? valid_0_104 : _GEN_2418; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3573 = unuse_way == 2'h2 ? valid_0_105 : _GEN_2419; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3574 = unuse_way == 2'h2 ? valid_0_106 : _GEN_2420; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3575 = unuse_way == 2'h2 ? valid_0_107 : _GEN_2421; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3576 = unuse_way == 2'h2 ? valid_0_108 : _GEN_2422; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3577 = unuse_way == 2'h2 ? valid_0_109 : _GEN_2423; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3578 = unuse_way == 2'h2 ? valid_0_110 : _GEN_2424; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3579 = unuse_way == 2'h2 ? valid_0_111 : _GEN_2425; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3580 = unuse_way == 2'h2 ? valid_0_112 : _GEN_2426; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3581 = unuse_way == 2'h2 ? valid_0_113 : _GEN_2427; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3582 = unuse_way == 2'h2 ? valid_0_114 : _GEN_2428; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3583 = unuse_way == 2'h2 ? valid_0_115 : _GEN_2429; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3584 = unuse_way == 2'h2 ? valid_0_116 : _GEN_2430; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3585 = unuse_way == 2'h2 ? valid_0_117 : _GEN_2431; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3586 = unuse_way == 2'h2 ? valid_0_118 : _GEN_2432; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3587 = unuse_way == 2'h2 ? valid_0_119 : _GEN_2433; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3588 = unuse_way == 2'h2 ? valid_0_120 : _GEN_2434; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3589 = unuse_way == 2'h2 ? valid_0_121 : _GEN_2435; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3590 = unuse_way == 2'h2 ? valid_0_122 : _GEN_2436; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3591 = unuse_way == 2'h2 ? valid_0_123 : _GEN_2437; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3592 = unuse_way == 2'h2 ? valid_0_124 : _GEN_2438; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3593 = unuse_way == 2'h2 ? valid_0_125 : _GEN_2439; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3594 = unuse_way == 2'h2 ? valid_0_126 : _GEN_2440; // @[i_cache.scala 21:26 91:40]
  wire  _GEN_3595 = unuse_way == 2'h2 ? valid_0_127 : _GEN_2441; // @[i_cache.scala 21:26 91:40]
  wire [63:0] _GEN_3596 = unuse_way == 2'h1 ? _GEN_522 : _GEN_3212; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3597 = unuse_way == 2'h1 ? _GEN_523 : _GEN_3213; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3598 = unuse_way == 2'h1 ? _GEN_524 : _GEN_3214; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3599 = unuse_way == 2'h1 ? _GEN_525 : _GEN_3215; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3600 = unuse_way == 2'h1 ? _GEN_526 : _GEN_3216; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3601 = unuse_way == 2'h1 ? _GEN_527 : _GEN_3217; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3602 = unuse_way == 2'h1 ? _GEN_528 : _GEN_3218; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3603 = unuse_way == 2'h1 ? _GEN_529 : _GEN_3219; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3604 = unuse_way == 2'h1 ? _GEN_530 : _GEN_3220; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3605 = unuse_way == 2'h1 ? _GEN_531 : _GEN_3221; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3606 = unuse_way == 2'h1 ? _GEN_532 : _GEN_3222; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3607 = unuse_way == 2'h1 ? _GEN_533 : _GEN_3223; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3608 = unuse_way == 2'h1 ? _GEN_534 : _GEN_3224; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3609 = unuse_way == 2'h1 ? _GEN_535 : _GEN_3225; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3610 = unuse_way == 2'h1 ? _GEN_536 : _GEN_3226; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3611 = unuse_way == 2'h1 ? _GEN_537 : _GEN_3227; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3612 = unuse_way == 2'h1 ? _GEN_538 : _GEN_3228; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3613 = unuse_way == 2'h1 ? _GEN_539 : _GEN_3229; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3614 = unuse_way == 2'h1 ? _GEN_540 : _GEN_3230; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3615 = unuse_way == 2'h1 ? _GEN_541 : _GEN_3231; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3616 = unuse_way == 2'h1 ? _GEN_542 : _GEN_3232; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3617 = unuse_way == 2'h1 ? _GEN_543 : _GEN_3233; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3618 = unuse_way == 2'h1 ? _GEN_544 : _GEN_3234; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3619 = unuse_way == 2'h1 ? _GEN_545 : _GEN_3235; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3620 = unuse_way == 2'h1 ? _GEN_546 : _GEN_3236; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3621 = unuse_way == 2'h1 ? _GEN_547 : _GEN_3237; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3622 = unuse_way == 2'h1 ? _GEN_548 : _GEN_3238; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3623 = unuse_way == 2'h1 ? _GEN_549 : _GEN_3239; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3624 = unuse_way == 2'h1 ? _GEN_550 : _GEN_3240; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3625 = unuse_way == 2'h1 ? _GEN_551 : _GEN_3241; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3626 = unuse_way == 2'h1 ? _GEN_552 : _GEN_3242; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3627 = unuse_way == 2'h1 ? _GEN_553 : _GEN_3243; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3628 = unuse_way == 2'h1 ? _GEN_554 : _GEN_3244; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3629 = unuse_way == 2'h1 ? _GEN_555 : _GEN_3245; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3630 = unuse_way == 2'h1 ? _GEN_556 : _GEN_3246; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3631 = unuse_way == 2'h1 ? _GEN_557 : _GEN_3247; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3632 = unuse_way == 2'h1 ? _GEN_558 : _GEN_3248; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3633 = unuse_way == 2'h1 ? _GEN_559 : _GEN_3249; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3634 = unuse_way == 2'h1 ? _GEN_560 : _GEN_3250; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3635 = unuse_way == 2'h1 ? _GEN_561 : _GEN_3251; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3636 = unuse_way == 2'h1 ? _GEN_562 : _GEN_3252; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3637 = unuse_way == 2'h1 ? _GEN_563 : _GEN_3253; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3638 = unuse_way == 2'h1 ? _GEN_564 : _GEN_3254; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3639 = unuse_way == 2'h1 ? _GEN_565 : _GEN_3255; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3640 = unuse_way == 2'h1 ? _GEN_566 : _GEN_3256; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3641 = unuse_way == 2'h1 ? _GEN_567 : _GEN_3257; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3642 = unuse_way == 2'h1 ? _GEN_568 : _GEN_3258; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3643 = unuse_way == 2'h1 ? _GEN_569 : _GEN_3259; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3644 = unuse_way == 2'h1 ? _GEN_570 : _GEN_3260; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3645 = unuse_way == 2'h1 ? _GEN_571 : _GEN_3261; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3646 = unuse_way == 2'h1 ? _GEN_572 : _GEN_3262; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3647 = unuse_way == 2'h1 ? _GEN_573 : _GEN_3263; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3648 = unuse_way == 2'h1 ? _GEN_574 : _GEN_3264; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3649 = unuse_way == 2'h1 ? _GEN_575 : _GEN_3265; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3650 = unuse_way == 2'h1 ? _GEN_576 : _GEN_3266; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3651 = unuse_way == 2'h1 ? _GEN_577 : _GEN_3267; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3652 = unuse_way == 2'h1 ? _GEN_578 : _GEN_3268; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3653 = unuse_way == 2'h1 ? _GEN_579 : _GEN_3269; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3654 = unuse_way == 2'h1 ? _GEN_580 : _GEN_3270; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3655 = unuse_way == 2'h1 ? _GEN_581 : _GEN_3271; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3656 = unuse_way == 2'h1 ? _GEN_582 : _GEN_3272; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3657 = unuse_way == 2'h1 ? _GEN_583 : _GEN_3273; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3658 = unuse_way == 2'h1 ? _GEN_584 : _GEN_3274; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3659 = unuse_way == 2'h1 ? _GEN_585 : _GEN_3275; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3660 = unuse_way == 2'h1 ? _GEN_586 : _GEN_3276; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3661 = unuse_way == 2'h1 ? _GEN_587 : _GEN_3277; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3662 = unuse_way == 2'h1 ? _GEN_588 : _GEN_3278; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3663 = unuse_way == 2'h1 ? _GEN_589 : _GEN_3279; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3664 = unuse_way == 2'h1 ? _GEN_590 : _GEN_3280; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3665 = unuse_way == 2'h1 ? _GEN_591 : _GEN_3281; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3666 = unuse_way == 2'h1 ? _GEN_592 : _GEN_3282; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3667 = unuse_way == 2'h1 ? _GEN_593 : _GEN_3283; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3668 = unuse_way == 2'h1 ? _GEN_594 : _GEN_3284; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3669 = unuse_way == 2'h1 ? _GEN_595 : _GEN_3285; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3670 = unuse_way == 2'h1 ? _GEN_596 : _GEN_3286; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3671 = unuse_way == 2'h1 ? _GEN_597 : _GEN_3287; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3672 = unuse_way == 2'h1 ? _GEN_598 : _GEN_3288; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3673 = unuse_way == 2'h1 ? _GEN_599 : _GEN_3289; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3674 = unuse_way == 2'h1 ? _GEN_600 : _GEN_3290; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3675 = unuse_way == 2'h1 ? _GEN_601 : _GEN_3291; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3676 = unuse_way == 2'h1 ? _GEN_602 : _GEN_3292; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3677 = unuse_way == 2'h1 ? _GEN_603 : _GEN_3293; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3678 = unuse_way == 2'h1 ? _GEN_604 : _GEN_3294; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3679 = unuse_way == 2'h1 ? _GEN_605 : _GEN_3295; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3680 = unuse_way == 2'h1 ? _GEN_606 : _GEN_3296; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3681 = unuse_way == 2'h1 ? _GEN_607 : _GEN_3297; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3682 = unuse_way == 2'h1 ? _GEN_608 : _GEN_3298; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3683 = unuse_way == 2'h1 ? _GEN_609 : _GEN_3299; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3684 = unuse_way == 2'h1 ? _GEN_610 : _GEN_3300; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3685 = unuse_way == 2'h1 ? _GEN_611 : _GEN_3301; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3686 = unuse_way == 2'h1 ? _GEN_612 : _GEN_3302; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3687 = unuse_way == 2'h1 ? _GEN_613 : _GEN_3303; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3688 = unuse_way == 2'h1 ? _GEN_614 : _GEN_3304; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3689 = unuse_way == 2'h1 ? _GEN_615 : _GEN_3305; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3690 = unuse_way == 2'h1 ? _GEN_616 : _GEN_3306; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3691 = unuse_way == 2'h1 ? _GEN_617 : _GEN_3307; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3692 = unuse_way == 2'h1 ? _GEN_618 : _GEN_3308; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3693 = unuse_way == 2'h1 ? _GEN_619 : _GEN_3309; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3694 = unuse_way == 2'h1 ? _GEN_620 : _GEN_3310; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3695 = unuse_way == 2'h1 ? _GEN_621 : _GEN_3311; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3696 = unuse_way == 2'h1 ? _GEN_622 : _GEN_3312; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3697 = unuse_way == 2'h1 ? _GEN_623 : _GEN_3313; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3698 = unuse_way == 2'h1 ? _GEN_624 : _GEN_3314; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3699 = unuse_way == 2'h1 ? _GEN_625 : _GEN_3315; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3700 = unuse_way == 2'h1 ? _GEN_626 : _GEN_3316; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3701 = unuse_way == 2'h1 ? _GEN_627 : _GEN_3317; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3702 = unuse_way == 2'h1 ? _GEN_628 : _GEN_3318; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3703 = unuse_way == 2'h1 ? _GEN_629 : _GEN_3319; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3704 = unuse_way == 2'h1 ? _GEN_630 : _GEN_3320; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3705 = unuse_way == 2'h1 ? _GEN_631 : _GEN_3321; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3706 = unuse_way == 2'h1 ? _GEN_632 : _GEN_3322; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3707 = unuse_way == 2'h1 ? _GEN_633 : _GEN_3323; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3708 = unuse_way == 2'h1 ? _GEN_634 : _GEN_3324; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3709 = unuse_way == 2'h1 ? _GEN_635 : _GEN_3325; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3710 = unuse_way == 2'h1 ? _GEN_636 : _GEN_3326; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3711 = unuse_way == 2'h1 ? _GEN_637 : _GEN_3327; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3712 = unuse_way == 2'h1 ? _GEN_638 : _GEN_3328; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3713 = unuse_way == 2'h1 ? _GEN_639 : _GEN_3329; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3714 = unuse_way == 2'h1 ? _GEN_640 : _GEN_3330; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3715 = unuse_way == 2'h1 ? _GEN_641 : _GEN_3331; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3716 = unuse_way == 2'h1 ? _GEN_642 : _GEN_3332; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3717 = unuse_way == 2'h1 ? _GEN_643 : _GEN_3333; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3718 = unuse_way == 2'h1 ? _GEN_644 : _GEN_3334; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3719 = unuse_way == 2'h1 ? _GEN_645 : _GEN_3335; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3720 = unuse_way == 2'h1 ? _GEN_646 : _GEN_3336; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3721 = unuse_way == 2'h1 ? _GEN_647 : _GEN_3337; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3722 = unuse_way == 2'h1 ? _GEN_648 : _GEN_3338; // @[i_cache.scala 86:34]
  wire [63:0] _GEN_3723 = unuse_way == 2'h1 ? _GEN_649 : _GEN_3339; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3724 = unuse_way == 2'h1 ? _GEN_650 : _GEN_3340; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3725 = unuse_way == 2'h1 ? _GEN_651 : _GEN_3341; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3726 = unuse_way == 2'h1 ? _GEN_652 : _GEN_3342; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3727 = unuse_way == 2'h1 ? _GEN_653 : _GEN_3343; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3728 = unuse_way == 2'h1 ? _GEN_654 : _GEN_3344; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3729 = unuse_way == 2'h1 ? _GEN_655 : _GEN_3345; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3730 = unuse_way == 2'h1 ? _GEN_656 : _GEN_3346; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3731 = unuse_way == 2'h1 ? _GEN_657 : _GEN_3347; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3732 = unuse_way == 2'h1 ? _GEN_658 : _GEN_3348; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3733 = unuse_way == 2'h1 ? _GEN_659 : _GEN_3349; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3734 = unuse_way == 2'h1 ? _GEN_660 : _GEN_3350; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3735 = unuse_way == 2'h1 ? _GEN_661 : _GEN_3351; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3736 = unuse_way == 2'h1 ? _GEN_662 : _GEN_3352; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3737 = unuse_way == 2'h1 ? _GEN_663 : _GEN_3353; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3738 = unuse_way == 2'h1 ? _GEN_664 : _GEN_3354; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3739 = unuse_way == 2'h1 ? _GEN_665 : _GEN_3355; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3740 = unuse_way == 2'h1 ? _GEN_666 : _GEN_3356; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3741 = unuse_way == 2'h1 ? _GEN_667 : _GEN_3357; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3742 = unuse_way == 2'h1 ? _GEN_668 : _GEN_3358; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3743 = unuse_way == 2'h1 ? _GEN_669 : _GEN_3359; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3744 = unuse_way == 2'h1 ? _GEN_670 : _GEN_3360; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3745 = unuse_way == 2'h1 ? _GEN_671 : _GEN_3361; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3746 = unuse_way == 2'h1 ? _GEN_672 : _GEN_3362; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3747 = unuse_way == 2'h1 ? _GEN_673 : _GEN_3363; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3748 = unuse_way == 2'h1 ? _GEN_674 : _GEN_3364; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3749 = unuse_way == 2'h1 ? _GEN_675 : _GEN_3365; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3750 = unuse_way == 2'h1 ? _GEN_676 : _GEN_3366; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3751 = unuse_way == 2'h1 ? _GEN_677 : _GEN_3367; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3752 = unuse_way == 2'h1 ? _GEN_678 : _GEN_3368; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3753 = unuse_way == 2'h1 ? _GEN_679 : _GEN_3369; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3754 = unuse_way == 2'h1 ? _GEN_680 : _GEN_3370; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3755 = unuse_way == 2'h1 ? _GEN_681 : _GEN_3371; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3756 = unuse_way == 2'h1 ? _GEN_682 : _GEN_3372; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3757 = unuse_way == 2'h1 ? _GEN_683 : _GEN_3373; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3758 = unuse_way == 2'h1 ? _GEN_684 : _GEN_3374; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3759 = unuse_way == 2'h1 ? _GEN_685 : _GEN_3375; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3760 = unuse_way == 2'h1 ? _GEN_686 : _GEN_3376; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3761 = unuse_way == 2'h1 ? _GEN_687 : _GEN_3377; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3762 = unuse_way == 2'h1 ? _GEN_688 : _GEN_3378; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3763 = unuse_way == 2'h1 ? _GEN_689 : _GEN_3379; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3764 = unuse_way == 2'h1 ? _GEN_690 : _GEN_3380; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3765 = unuse_way == 2'h1 ? _GEN_691 : _GEN_3381; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3766 = unuse_way == 2'h1 ? _GEN_692 : _GEN_3382; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3767 = unuse_way == 2'h1 ? _GEN_693 : _GEN_3383; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3768 = unuse_way == 2'h1 ? _GEN_694 : _GEN_3384; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3769 = unuse_way == 2'h1 ? _GEN_695 : _GEN_3385; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3770 = unuse_way == 2'h1 ? _GEN_696 : _GEN_3386; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3771 = unuse_way == 2'h1 ? _GEN_697 : _GEN_3387; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3772 = unuse_way == 2'h1 ? _GEN_698 : _GEN_3388; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3773 = unuse_way == 2'h1 ? _GEN_699 : _GEN_3389; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3774 = unuse_way == 2'h1 ? _GEN_700 : _GEN_3390; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3775 = unuse_way == 2'h1 ? _GEN_701 : _GEN_3391; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3776 = unuse_way == 2'h1 ? _GEN_702 : _GEN_3392; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3777 = unuse_way == 2'h1 ? _GEN_703 : _GEN_3393; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3778 = unuse_way == 2'h1 ? _GEN_704 : _GEN_3394; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3779 = unuse_way == 2'h1 ? _GEN_705 : _GEN_3395; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3780 = unuse_way == 2'h1 ? _GEN_706 : _GEN_3396; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3781 = unuse_way == 2'h1 ? _GEN_707 : _GEN_3397; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3782 = unuse_way == 2'h1 ? _GEN_708 : _GEN_3398; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3783 = unuse_way == 2'h1 ? _GEN_709 : _GEN_3399; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3784 = unuse_way == 2'h1 ? _GEN_710 : _GEN_3400; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3785 = unuse_way == 2'h1 ? _GEN_711 : _GEN_3401; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3786 = unuse_way == 2'h1 ? _GEN_712 : _GEN_3402; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3787 = unuse_way == 2'h1 ? _GEN_713 : _GEN_3403; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3788 = unuse_way == 2'h1 ? _GEN_714 : _GEN_3404; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3789 = unuse_way == 2'h1 ? _GEN_715 : _GEN_3405; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3790 = unuse_way == 2'h1 ? _GEN_716 : _GEN_3406; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3791 = unuse_way == 2'h1 ? _GEN_717 : _GEN_3407; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3792 = unuse_way == 2'h1 ? _GEN_718 : _GEN_3408; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3793 = unuse_way == 2'h1 ? _GEN_719 : _GEN_3409; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3794 = unuse_way == 2'h1 ? _GEN_720 : _GEN_3410; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3795 = unuse_way == 2'h1 ? _GEN_721 : _GEN_3411; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3796 = unuse_way == 2'h1 ? _GEN_722 : _GEN_3412; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3797 = unuse_way == 2'h1 ? _GEN_723 : _GEN_3413; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3798 = unuse_way == 2'h1 ? _GEN_724 : _GEN_3414; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3799 = unuse_way == 2'h1 ? _GEN_725 : _GEN_3415; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3800 = unuse_way == 2'h1 ? _GEN_726 : _GEN_3416; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3801 = unuse_way == 2'h1 ? _GEN_727 : _GEN_3417; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3802 = unuse_way == 2'h1 ? _GEN_728 : _GEN_3418; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3803 = unuse_way == 2'h1 ? _GEN_729 : _GEN_3419; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3804 = unuse_way == 2'h1 ? _GEN_730 : _GEN_3420; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3805 = unuse_way == 2'h1 ? _GEN_731 : _GEN_3421; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3806 = unuse_way == 2'h1 ? _GEN_732 : _GEN_3422; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3807 = unuse_way == 2'h1 ? _GEN_733 : _GEN_3423; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3808 = unuse_way == 2'h1 ? _GEN_734 : _GEN_3424; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3809 = unuse_way == 2'h1 ? _GEN_735 : _GEN_3425; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3810 = unuse_way == 2'h1 ? _GEN_736 : _GEN_3426; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3811 = unuse_way == 2'h1 ? _GEN_737 : _GEN_3427; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3812 = unuse_way == 2'h1 ? _GEN_738 : _GEN_3428; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3813 = unuse_way == 2'h1 ? _GEN_739 : _GEN_3429; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3814 = unuse_way == 2'h1 ? _GEN_740 : _GEN_3430; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3815 = unuse_way == 2'h1 ? _GEN_741 : _GEN_3431; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3816 = unuse_way == 2'h1 ? _GEN_742 : _GEN_3432; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3817 = unuse_way == 2'h1 ? _GEN_743 : _GEN_3433; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3818 = unuse_way == 2'h1 ? _GEN_744 : _GEN_3434; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3819 = unuse_way == 2'h1 ? _GEN_745 : _GEN_3435; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3820 = unuse_way == 2'h1 ? _GEN_746 : _GEN_3436; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3821 = unuse_way == 2'h1 ? _GEN_747 : _GEN_3437; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3822 = unuse_way == 2'h1 ? _GEN_748 : _GEN_3438; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3823 = unuse_way == 2'h1 ? _GEN_749 : _GEN_3439; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3824 = unuse_way == 2'h1 ? _GEN_750 : _GEN_3440; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3825 = unuse_way == 2'h1 ? _GEN_751 : _GEN_3441; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3826 = unuse_way == 2'h1 ? _GEN_752 : _GEN_3442; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3827 = unuse_way == 2'h1 ? _GEN_753 : _GEN_3443; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3828 = unuse_way == 2'h1 ? _GEN_754 : _GEN_3444; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3829 = unuse_way == 2'h1 ? _GEN_755 : _GEN_3445; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3830 = unuse_way == 2'h1 ? _GEN_756 : _GEN_3446; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3831 = unuse_way == 2'h1 ? _GEN_757 : _GEN_3447; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3832 = unuse_way == 2'h1 ? _GEN_758 : _GEN_3448; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3833 = unuse_way == 2'h1 ? _GEN_759 : _GEN_3449; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3834 = unuse_way == 2'h1 ? _GEN_760 : _GEN_3450; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3835 = unuse_way == 2'h1 ? _GEN_761 : _GEN_3451; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3836 = unuse_way == 2'h1 ? _GEN_762 : _GEN_3452; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3837 = unuse_way == 2'h1 ? _GEN_763 : _GEN_3453; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3838 = unuse_way == 2'h1 ? _GEN_764 : _GEN_3454; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3839 = unuse_way == 2'h1 ? _GEN_765 : _GEN_3455; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3840 = unuse_way == 2'h1 ? _GEN_766 : _GEN_3456; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3841 = unuse_way == 2'h1 ? _GEN_767 : _GEN_3457; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3842 = unuse_way == 2'h1 ? _GEN_768 : _GEN_3458; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3843 = unuse_way == 2'h1 ? _GEN_769 : _GEN_3459; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3844 = unuse_way == 2'h1 ? _GEN_770 : _GEN_3460; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3845 = unuse_way == 2'h1 ? _GEN_771 : _GEN_3461; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3846 = unuse_way == 2'h1 ? _GEN_772 : _GEN_3462; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3847 = unuse_way == 2'h1 ? _GEN_773 : _GEN_3463; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3848 = unuse_way == 2'h1 ? _GEN_774 : _GEN_3464; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3849 = unuse_way == 2'h1 ? _GEN_775 : _GEN_3465; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3850 = unuse_way == 2'h1 ? _GEN_776 : _GEN_3466; // @[i_cache.scala 86:34]
  wire [31:0] _GEN_3851 = unuse_way == 2'h1 ? _GEN_777 : _GEN_3467; // @[i_cache.scala 86:34]
  wire  _GEN_3852 = unuse_way == 2'h1 ? _GEN_778 : _GEN_3468; // @[i_cache.scala 86:34]
  wire  _GEN_3853 = unuse_way == 2'h1 ? _GEN_779 : _GEN_3469; // @[i_cache.scala 86:34]
  wire  _GEN_3854 = unuse_way == 2'h1 ? _GEN_780 : _GEN_3470; // @[i_cache.scala 86:34]
  wire  _GEN_3855 = unuse_way == 2'h1 ? _GEN_781 : _GEN_3471; // @[i_cache.scala 86:34]
  wire  _GEN_3856 = unuse_way == 2'h1 ? _GEN_782 : _GEN_3472; // @[i_cache.scala 86:34]
  wire  _GEN_3857 = unuse_way == 2'h1 ? _GEN_783 : _GEN_3473; // @[i_cache.scala 86:34]
  wire  _GEN_3858 = unuse_way == 2'h1 ? _GEN_784 : _GEN_3474; // @[i_cache.scala 86:34]
  wire  _GEN_3859 = unuse_way == 2'h1 ? _GEN_785 : _GEN_3475; // @[i_cache.scala 86:34]
  wire  _GEN_3860 = unuse_way == 2'h1 ? _GEN_786 : _GEN_3476; // @[i_cache.scala 86:34]
  wire  _GEN_3861 = unuse_way == 2'h1 ? _GEN_787 : _GEN_3477; // @[i_cache.scala 86:34]
  wire  _GEN_3862 = unuse_way == 2'h1 ? _GEN_788 : _GEN_3478; // @[i_cache.scala 86:34]
  wire  _GEN_3863 = unuse_way == 2'h1 ? _GEN_789 : _GEN_3479; // @[i_cache.scala 86:34]
  wire  _GEN_3864 = unuse_way == 2'h1 ? _GEN_790 : _GEN_3480; // @[i_cache.scala 86:34]
  wire  _GEN_3865 = unuse_way == 2'h1 ? _GEN_791 : _GEN_3481; // @[i_cache.scala 86:34]
  wire  _GEN_3866 = unuse_way == 2'h1 ? _GEN_792 : _GEN_3482; // @[i_cache.scala 86:34]
  wire  _GEN_3867 = unuse_way == 2'h1 ? _GEN_793 : _GEN_3483; // @[i_cache.scala 86:34]
  wire  _GEN_3868 = unuse_way == 2'h1 ? _GEN_794 : _GEN_3484; // @[i_cache.scala 86:34]
  wire  _GEN_3869 = unuse_way == 2'h1 ? _GEN_795 : _GEN_3485; // @[i_cache.scala 86:34]
  wire  _GEN_3870 = unuse_way == 2'h1 ? _GEN_796 : _GEN_3486; // @[i_cache.scala 86:34]
  wire  _GEN_3871 = unuse_way == 2'h1 ? _GEN_797 : _GEN_3487; // @[i_cache.scala 86:34]
  wire  _GEN_3872 = unuse_way == 2'h1 ? _GEN_798 : _GEN_3488; // @[i_cache.scala 86:34]
  wire  _GEN_3873 = unuse_way == 2'h1 ? _GEN_799 : _GEN_3489; // @[i_cache.scala 86:34]
  wire  _GEN_3874 = unuse_way == 2'h1 ? _GEN_800 : _GEN_3490; // @[i_cache.scala 86:34]
  wire  _GEN_3875 = unuse_way == 2'h1 ? _GEN_801 : _GEN_3491; // @[i_cache.scala 86:34]
  wire  _GEN_3876 = unuse_way == 2'h1 ? _GEN_802 : _GEN_3492; // @[i_cache.scala 86:34]
  wire  _GEN_3877 = unuse_way == 2'h1 ? _GEN_803 : _GEN_3493; // @[i_cache.scala 86:34]
  wire  _GEN_3878 = unuse_way == 2'h1 ? _GEN_804 : _GEN_3494; // @[i_cache.scala 86:34]
  wire  _GEN_3879 = unuse_way == 2'h1 ? _GEN_805 : _GEN_3495; // @[i_cache.scala 86:34]
  wire  _GEN_3880 = unuse_way == 2'h1 ? _GEN_806 : _GEN_3496; // @[i_cache.scala 86:34]
  wire  _GEN_3881 = unuse_way == 2'h1 ? _GEN_807 : _GEN_3497; // @[i_cache.scala 86:34]
  wire  _GEN_3882 = unuse_way == 2'h1 ? _GEN_808 : _GEN_3498; // @[i_cache.scala 86:34]
  wire  _GEN_3883 = unuse_way == 2'h1 ? _GEN_809 : _GEN_3499; // @[i_cache.scala 86:34]
  wire  _GEN_3884 = unuse_way == 2'h1 ? _GEN_810 : _GEN_3500; // @[i_cache.scala 86:34]
  wire  _GEN_3885 = unuse_way == 2'h1 ? _GEN_811 : _GEN_3501; // @[i_cache.scala 86:34]
  wire  _GEN_3886 = unuse_way == 2'h1 ? _GEN_812 : _GEN_3502; // @[i_cache.scala 86:34]
  wire  _GEN_3887 = unuse_way == 2'h1 ? _GEN_813 : _GEN_3503; // @[i_cache.scala 86:34]
  wire  _GEN_3888 = unuse_way == 2'h1 ? _GEN_814 : _GEN_3504; // @[i_cache.scala 86:34]
  wire  _GEN_3889 = unuse_way == 2'h1 ? _GEN_815 : _GEN_3505; // @[i_cache.scala 86:34]
  wire  _GEN_3890 = unuse_way == 2'h1 ? _GEN_816 : _GEN_3506; // @[i_cache.scala 86:34]
  wire  _GEN_3891 = unuse_way == 2'h1 ? _GEN_817 : _GEN_3507; // @[i_cache.scala 86:34]
  wire  _GEN_3892 = unuse_way == 2'h1 ? _GEN_818 : _GEN_3508; // @[i_cache.scala 86:34]
  wire  _GEN_3893 = unuse_way == 2'h1 ? _GEN_819 : _GEN_3509; // @[i_cache.scala 86:34]
  wire  _GEN_3894 = unuse_way == 2'h1 ? _GEN_820 : _GEN_3510; // @[i_cache.scala 86:34]
  wire  _GEN_3895 = unuse_way == 2'h1 ? _GEN_821 : _GEN_3511; // @[i_cache.scala 86:34]
  wire  _GEN_3896 = unuse_way == 2'h1 ? _GEN_822 : _GEN_3512; // @[i_cache.scala 86:34]
  wire  _GEN_3897 = unuse_way == 2'h1 ? _GEN_823 : _GEN_3513; // @[i_cache.scala 86:34]
  wire  _GEN_3898 = unuse_way == 2'h1 ? _GEN_824 : _GEN_3514; // @[i_cache.scala 86:34]
  wire  _GEN_3899 = unuse_way == 2'h1 ? _GEN_825 : _GEN_3515; // @[i_cache.scala 86:34]
  wire  _GEN_3900 = unuse_way == 2'h1 ? _GEN_826 : _GEN_3516; // @[i_cache.scala 86:34]
  wire  _GEN_3901 = unuse_way == 2'h1 ? _GEN_827 : _GEN_3517; // @[i_cache.scala 86:34]
  wire  _GEN_3902 = unuse_way == 2'h1 ? _GEN_828 : _GEN_3518; // @[i_cache.scala 86:34]
  wire  _GEN_3903 = unuse_way == 2'h1 ? _GEN_829 : _GEN_3519; // @[i_cache.scala 86:34]
  wire  _GEN_3904 = unuse_way == 2'h1 ? _GEN_830 : _GEN_3520; // @[i_cache.scala 86:34]
  wire  _GEN_3905 = unuse_way == 2'h1 ? _GEN_831 : _GEN_3521; // @[i_cache.scala 86:34]
  wire  _GEN_3906 = unuse_way == 2'h1 ? _GEN_832 : _GEN_3522; // @[i_cache.scala 86:34]
  wire  _GEN_3907 = unuse_way == 2'h1 ? _GEN_833 : _GEN_3523; // @[i_cache.scala 86:34]
  wire  _GEN_3908 = unuse_way == 2'h1 ? _GEN_834 : _GEN_3524; // @[i_cache.scala 86:34]
  wire  _GEN_3909 = unuse_way == 2'h1 ? _GEN_835 : _GEN_3525; // @[i_cache.scala 86:34]
  wire  _GEN_3910 = unuse_way == 2'h1 ? _GEN_836 : _GEN_3526; // @[i_cache.scala 86:34]
  wire  _GEN_3911 = unuse_way == 2'h1 ? _GEN_837 : _GEN_3527; // @[i_cache.scala 86:34]
  wire  _GEN_3912 = unuse_way == 2'h1 ? _GEN_838 : _GEN_3528; // @[i_cache.scala 86:34]
  wire  _GEN_3913 = unuse_way == 2'h1 ? _GEN_839 : _GEN_3529; // @[i_cache.scala 86:34]
  wire  _GEN_3914 = unuse_way == 2'h1 ? _GEN_840 : _GEN_3530; // @[i_cache.scala 86:34]
  wire  _GEN_3915 = unuse_way == 2'h1 ? _GEN_841 : _GEN_3531; // @[i_cache.scala 86:34]
  wire  _GEN_3916 = unuse_way == 2'h1 ? _GEN_842 : _GEN_3532; // @[i_cache.scala 86:34]
  wire  _GEN_3917 = unuse_way == 2'h1 ? _GEN_843 : _GEN_3533; // @[i_cache.scala 86:34]
  wire  _GEN_3918 = unuse_way == 2'h1 ? _GEN_844 : _GEN_3534; // @[i_cache.scala 86:34]
  wire  _GEN_3919 = unuse_way == 2'h1 ? _GEN_845 : _GEN_3535; // @[i_cache.scala 86:34]
  wire  _GEN_3920 = unuse_way == 2'h1 ? _GEN_846 : _GEN_3536; // @[i_cache.scala 86:34]
  wire  _GEN_3921 = unuse_way == 2'h1 ? _GEN_847 : _GEN_3537; // @[i_cache.scala 86:34]
  wire  _GEN_3922 = unuse_way == 2'h1 ? _GEN_848 : _GEN_3538; // @[i_cache.scala 86:34]
  wire  _GEN_3923 = unuse_way == 2'h1 ? _GEN_849 : _GEN_3539; // @[i_cache.scala 86:34]
  wire  _GEN_3924 = unuse_way == 2'h1 ? _GEN_850 : _GEN_3540; // @[i_cache.scala 86:34]
  wire  _GEN_3925 = unuse_way == 2'h1 ? _GEN_851 : _GEN_3541; // @[i_cache.scala 86:34]
  wire  _GEN_3926 = unuse_way == 2'h1 ? _GEN_852 : _GEN_3542; // @[i_cache.scala 86:34]
  wire  _GEN_3927 = unuse_way == 2'h1 ? _GEN_853 : _GEN_3543; // @[i_cache.scala 86:34]
  wire  _GEN_3928 = unuse_way == 2'h1 ? _GEN_854 : _GEN_3544; // @[i_cache.scala 86:34]
  wire  _GEN_3929 = unuse_way == 2'h1 ? _GEN_855 : _GEN_3545; // @[i_cache.scala 86:34]
  wire  _GEN_3930 = unuse_way == 2'h1 ? _GEN_856 : _GEN_3546; // @[i_cache.scala 86:34]
  wire  _GEN_3931 = unuse_way == 2'h1 ? _GEN_857 : _GEN_3547; // @[i_cache.scala 86:34]
  wire  _GEN_3932 = unuse_way == 2'h1 ? _GEN_858 : _GEN_3548; // @[i_cache.scala 86:34]
  wire  _GEN_3933 = unuse_way == 2'h1 ? _GEN_859 : _GEN_3549; // @[i_cache.scala 86:34]
  wire  _GEN_3934 = unuse_way == 2'h1 ? _GEN_860 : _GEN_3550; // @[i_cache.scala 86:34]
  wire  _GEN_3935 = unuse_way == 2'h1 ? _GEN_861 : _GEN_3551; // @[i_cache.scala 86:34]
  wire  _GEN_3936 = unuse_way == 2'h1 ? _GEN_862 : _GEN_3552; // @[i_cache.scala 86:34]
  wire  _GEN_3937 = unuse_way == 2'h1 ? _GEN_863 : _GEN_3553; // @[i_cache.scala 86:34]
  wire  _GEN_3938 = unuse_way == 2'h1 ? _GEN_864 : _GEN_3554; // @[i_cache.scala 86:34]
  wire  _GEN_3939 = unuse_way == 2'h1 ? _GEN_865 : _GEN_3555; // @[i_cache.scala 86:34]
  wire  _GEN_3940 = unuse_way == 2'h1 ? _GEN_866 : _GEN_3556; // @[i_cache.scala 86:34]
  wire  _GEN_3941 = unuse_way == 2'h1 ? _GEN_867 : _GEN_3557; // @[i_cache.scala 86:34]
  wire  _GEN_3942 = unuse_way == 2'h1 ? _GEN_868 : _GEN_3558; // @[i_cache.scala 86:34]
  wire  _GEN_3943 = unuse_way == 2'h1 ? _GEN_869 : _GEN_3559; // @[i_cache.scala 86:34]
  wire  _GEN_3944 = unuse_way == 2'h1 ? _GEN_870 : _GEN_3560; // @[i_cache.scala 86:34]
  wire  _GEN_3945 = unuse_way == 2'h1 ? _GEN_871 : _GEN_3561; // @[i_cache.scala 86:34]
  wire  _GEN_3946 = unuse_way == 2'h1 ? _GEN_872 : _GEN_3562; // @[i_cache.scala 86:34]
  wire  _GEN_3947 = unuse_way == 2'h1 ? _GEN_873 : _GEN_3563; // @[i_cache.scala 86:34]
  wire  _GEN_3948 = unuse_way == 2'h1 ? _GEN_874 : _GEN_3564; // @[i_cache.scala 86:34]
  wire  _GEN_3949 = unuse_way == 2'h1 ? _GEN_875 : _GEN_3565; // @[i_cache.scala 86:34]
  wire  _GEN_3950 = unuse_way == 2'h1 ? _GEN_876 : _GEN_3566; // @[i_cache.scala 86:34]
  wire  _GEN_3951 = unuse_way == 2'h1 ? _GEN_877 : _GEN_3567; // @[i_cache.scala 86:34]
  wire  _GEN_3952 = unuse_way == 2'h1 ? _GEN_878 : _GEN_3568; // @[i_cache.scala 86:34]
  wire  _GEN_3953 = unuse_way == 2'h1 ? _GEN_879 : _GEN_3569; // @[i_cache.scala 86:34]
  wire  _GEN_3954 = unuse_way == 2'h1 ? _GEN_880 : _GEN_3570; // @[i_cache.scala 86:34]
  wire  _GEN_3955 = unuse_way == 2'h1 ? _GEN_881 : _GEN_3571; // @[i_cache.scala 86:34]
  wire  _GEN_3956 = unuse_way == 2'h1 ? _GEN_882 : _GEN_3572; // @[i_cache.scala 86:34]
  wire  _GEN_3957 = unuse_way == 2'h1 ? _GEN_883 : _GEN_3573; // @[i_cache.scala 86:34]
  wire  _GEN_3958 = unuse_way == 2'h1 ? _GEN_884 : _GEN_3574; // @[i_cache.scala 86:34]
  wire  _GEN_3959 = unuse_way == 2'h1 ? _GEN_885 : _GEN_3575; // @[i_cache.scala 86:34]
  wire  _GEN_3960 = unuse_way == 2'h1 ? _GEN_886 : _GEN_3576; // @[i_cache.scala 86:34]
  wire  _GEN_3961 = unuse_way == 2'h1 ? _GEN_887 : _GEN_3577; // @[i_cache.scala 86:34]
  wire  _GEN_3962 = unuse_way == 2'h1 ? _GEN_888 : _GEN_3578; // @[i_cache.scala 86:34]
  wire  _GEN_3963 = unuse_way == 2'h1 ? _GEN_889 : _GEN_3579; // @[i_cache.scala 86:34]
  wire  _GEN_3964 = unuse_way == 2'h1 ? _GEN_890 : _GEN_3580; // @[i_cache.scala 86:34]
  wire  _GEN_3965 = unuse_way == 2'h1 ? _GEN_891 : _GEN_3581; // @[i_cache.scala 86:34]
  wire  _GEN_3966 = unuse_way == 2'h1 ? _GEN_892 : _GEN_3582; // @[i_cache.scala 86:34]
  wire  _GEN_3967 = unuse_way == 2'h1 ? _GEN_893 : _GEN_3583; // @[i_cache.scala 86:34]
  wire  _GEN_3968 = unuse_way == 2'h1 ? _GEN_894 : _GEN_3584; // @[i_cache.scala 86:34]
  wire  _GEN_3969 = unuse_way == 2'h1 ? _GEN_895 : _GEN_3585; // @[i_cache.scala 86:34]
  wire  _GEN_3970 = unuse_way == 2'h1 ? _GEN_896 : _GEN_3586; // @[i_cache.scala 86:34]
  wire  _GEN_3971 = unuse_way == 2'h1 ? _GEN_897 : _GEN_3587; // @[i_cache.scala 86:34]
  wire  _GEN_3972 = unuse_way == 2'h1 ? _GEN_898 : _GEN_3588; // @[i_cache.scala 86:34]
  wire  _GEN_3973 = unuse_way == 2'h1 ? _GEN_899 : _GEN_3589; // @[i_cache.scala 86:34]
  wire  _GEN_3974 = unuse_way == 2'h1 ? _GEN_900 : _GEN_3590; // @[i_cache.scala 86:34]
  wire  _GEN_3975 = unuse_way == 2'h1 ? _GEN_901 : _GEN_3591; // @[i_cache.scala 86:34]
  wire  _GEN_3976 = unuse_way == 2'h1 ? _GEN_902 : _GEN_3592; // @[i_cache.scala 86:34]
  wire  _GEN_3977 = unuse_way == 2'h1 ? _GEN_903 : _GEN_3593; // @[i_cache.scala 86:34]
  wire  _GEN_3978 = unuse_way == 2'h1 ? _GEN_904 : _GEN_3594; // @[i_cache.scala 86:34]
  wire  _GEN_3979 = unuse_way == 2'h1 ? _GEN_905 : _GEN_3595; // @[i_cache.scala 86:34]
  wire  _GEN_3980 = unuse_way == 2'h1 | _GEN_3211; // @[i_cache.scala 86:34 90:23]
  wire [63:0] _GEN_3981 = unuse_way == 2'h1 ? ram_1_0 : _GEN_2827; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3982 = unuse_way == 2'h1 ? ram_1_1 : _GEN_2828; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3983 = unuse_way == 2'h1 ? ram_1_2 : _GEN_2829; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3984 = unuse_way == 2'h1 ? ram_1_3 : _GEN_2830; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3985 = unuse_way == 2'h1 ? ram_1_4 : _GEN_2831; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3986 = unuse_way == 2'h1 ? ram_1_5 : _GEN_2832; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3987 = unuse_way == 2'h1 ? ram_1_6 : _GEN_2833; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3988 = unuse_way == 2'h1 ? ram_1_7 : _GEN_2834; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3989 = unuse_way == 2'h1 ? ram_1_8 : _GEN_2835; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3990 = unuse_way == 2'h1 ? ram_1_9 : _GEN_2836; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3991 = unuse_way == 2'h1 ? ram_1_10 : _GEN_2837; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3992 = unuse_way == 2'h1 ? ram_1_11 : _GEN_2838; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3993 = unuse_way == 2'h1 ? ram_1_12 : _GEN_2839; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3994 = unuse_way == 2'h1 ? ram_1_13 : _GEN_2840; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3995 = unuse_way == 2'h1 ? ram_1_14 : _GEN_2841; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3996 = unuse_way == 2'h1 ? ram_1_15 : _GEN_2842; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3997 = unuse_way == 2'h1 ? ram_1_16 : _GEN_2843; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3998 = unuse_way == 2'h1 ? ram_1_17 : _GEN_2844; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_3999 = unuse_way == 2'h1 ? ram_1_18 : _GEN_2845; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4000 = unuse_way == 2'h1 ? ram_1_19 : _GEN_2846; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4001 = unuse_way == 2'h1 ? ram_1_20 : _GEN_2847; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4002 = unuse_way == 2'h1 ? ram_1_21 : _GEN_2848; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4003 = unuse_way == 2'h1 ? ram_1_22 : _GEN_2849; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4004 = unuse_way == 2'h1 ? ram_1_23 : _GEN_2850; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4005 = unuse_way == 2'h1 ? ram_1_24 : _GEN_2851; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4006 = unuse_way == 2'h1 ? ram_1_25 : _GEN_2852; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4007 = unuse_way == 2'h1 ? ram_1_26 : _GEN_2853; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4008 = unuse_way == 2'h1 ? ram_1_27 : _GEN_2854; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4009 = unuse_way == 2'h1 ? ram_1_28 : _GEN_2855; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4010 = unuse_way == 2'h1 ? ram_1_29 : _GEN_2856; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4011 = unuse_way == 2'h1 ? ram_1_30 : _GEN_2857; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4012 = unuse_way == 2'h1 ? ram_1_31 : _GEN_2858; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4013 = unuse_way == 2'h1 ? ram_1_32 : _GEN_2859; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4014 = unuse_way == 2'h1 ? ram_1_33 : _GEN_2860; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4015 = unuse_way == 2'h1 ? ram_1_34 : _GEN_2861; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4016 = unuse_way == 2'h1 ? ram_1_35 : _GEN_2862; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4017 = unuse_way == 2'h1 ? ram_1_36 : _GEN_2863; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4018 = unuse_way == 2'h1 ? ram_1_37 : _GEN_2864; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4019 = unuse_way == 2'h1 ? ram_1_38 : _GEN_2865; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4020 = unuse_way == 2'h1 ? ram_1_39 : _GEN_2866; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4021 = unuse_way == 2'h1 ? ram_1_40 : _GEN_2867; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4022 = unuse_way == 2'h1 ? ram_1_41 : _GEN_2868; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4023 = unuse_way == 2'h1 ? ram_1_42 : _GEN_2869; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4024 = unuse_way == 2'h1 ? ram_1_43 : _GEN_2870; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4025 = unuse_way == 2'h1 ? ram_1_44 : _GEN_2871; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4026 = unuse_way == 2'h1 ? ram_1_45 : _GEN_2872; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4027 = unuse_way == 2'h1 ? ram_1_46 : _GEN_2873; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4028 = unuse_way == 2'h1 ? ram_1_47 : _GEN_2874; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4029 = unuse_way == 2'h1 ? ram_1_48 : _GEN_2875; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4030 = unuse_way == 2'h1 ? ram_1_49 : _GEN_2876; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4031 = unuse_way == 2'h1 ? ram_1_50 : _GEN_2877; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4032 = unuse_way == 2'h1 ? ram_1_51 : _GEN_2878; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4033 = unuse_way == 2'h1 ? ram_1_52 : _GEN_2879; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4034 = unuse_way == 2'h1 ? ram_1_53 : _GEN_2880; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4035 = unuse_way == 2'h1 ? ram_1_54 : _GEN_2881; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4036 = unuse_way == 2'h1 ? ram_1_55 : _GEN_2882; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4037 = unuse_way == 2'h1 ? ram_1_56 : _GEN_2883; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4038 = unuse_way == 2'h1 ? ram_1_57 : _GEN_2884; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4039 = unuse_way == 2'h1 ? ram_1_58 : _GEN_2885; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4040 = unuse_way == 2'h1 ? ram_1_59 : _GEN_2886; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4041 = unuse_way == 2'h1 ? ram_1_60 : _GEN_2887; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4042 = unuse_way == 2'h1 ? ram_1_61 : _GEN_2888; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4043 = unuse_way == 2'h1 ? ram_1_62 : _GEN_2889; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4044 = unuse_way == 2'h1 ? ram_1_63 : _GEN_2890; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4045 = unuse_way == 2'h1 ? ram_1_64 : _GEN_2891; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4046 = unuse_way == 2'h1 ? ram_1_65 : _GEN_2892; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4047 = unuse_way == 2'h1 ? ram_1_66 : _GEN_2893; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4048 = unuse_way == 2'h1 ? ram_1_67 : _GEN_2894; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4049 = unuse_way == 2'h1 ? ram_1_68 : _GEN_2895; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4050 = unuse_way == 2'h1 ? ram_1_69 : _GEN_2896; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4051 = unuse_way == 2'h1 ? ram_1_70 : _GEN_2897; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4052 = unuse_way == 2'h1 ? ram_1_71 : _GEN_2898; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4053 = unuse_way == 2'h1 ? ram_1_72 : _GEN_2899; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4054 = unuse_way == 2'h1 ? ram_1_73 : _GEN_2900; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4055 = unuse_way == 2'h1 ? ram_1_74 : _GEN_2901; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4056 = unuse_way == 2'h1 ? ram_1_75 : _GEN_2902; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4057 = unuse_way == 2'h1 ? ram_1_76 : _GEN_2903; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4058 = unuse_way == 2'h1 ? ram_1_77 : _GEN_2904; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4059 = unuse_way == 2'h1 ? ram_1_78 : _GEN_2905; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4060 = unuse_way == 2'h1 ? ram_1_79 : _GEN_2906; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4061 = unuse_way == 2'h1 ? ram_1_80 : _GEN_2907; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4062 = unuse_way == 2'h1 ? ram_1_81 : _GEN_2908; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4063 = unuse_way == 2'h1 ? ram_1_82 : _GEN_2909; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4064 = unuse_way == 2'h1 ? ram_1_83 : _GEN_2910; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4065 = unuse_way == 2'h1 ? ram_1_84 : _GEN_2911; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4066 = unuse_way == 2'h1 ? ram_1_85 : _GEN_2912; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4067 = unuse_way == 2'h1 ? ram_1_86 : _GEN_2913; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4068 = unuse_way == 2'h1 ? ram_1_87 : _GEN_2914; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4069 = unuse_way == 2'h1 ? ram_1_88 : _GEN_2915; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4070 = unuse_way == 2'h1 ? ram_1_89 : _GEN_2916; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4071 = unuse_way == 2'h1 ? ram_1_90 : _GEN_2917; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4072 = unuse_way == 2'h1 ? ram_1_91 : _GEN_2918; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4073 = unuse_way == 2'h1 ? ram_1_92 : _GEN_2919; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4074 = unuse_way == 2'h1 ? ram_1_93 : _GEN_2920; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4075 = unuse_way == 2'h1 ? ram_1_94 : _GEN_2921; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4076 = unuse_way == 2'h1 ? ram_1_95 : _GEN_2922; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4077 = unuse_way == 2'h1 ? ram_1_96 : _GEN_2923; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4078 = unuse_way == 2'h1 ? ram_1_97 : _GEN_2924; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4079 = unuse_way == 2'h1 ? ram_1_98 : _GEN_2925; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4080 = unuse_way == 2'h1 ? ram_1_99 : _GEN_2926; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4081 = unuse_way == 2'h1 ? ram_1_100 : _GEN_2927; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4082 = unuse_way == 2'h1 ? ram_1_101 : _GEN_2928; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4083 = unuse_way == 2'h1 ? ram_1_102 : _GEN_2929; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4084 = unuse_way == 2'h1 ? ram_1_103 : _GEN_2930; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4085 = unuse_way == 2'h1 ? ram_1_104 : _GEN_2931; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4086 = unuse_way == 2'h1 ? ram_1_105 : _GEN_2932; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4087 = unuse_way == 2'h1 ? ram_1_106 : _GEN_2933; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4088 = unuse_way == 2'h1 ? ram_1_107 : _GEN_2934; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4089 = unuse_way == 2'h1 ? ram_1_108 : _GEN_2935; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4090 = unuse_way == 2'h1 ? ram_1_109 : _GEN_2936; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4091 = unuse_way == 2'h1 ? ram_1_110 : _GEN_2937; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4092 = unuse_way == 2'h1 ? ram_1_111 : _GEN_2938; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4093 = unuse_way == 2'h1 ? ram_1_112 : _GEN_2939; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4094 = unuse_way == 2'h1 ? ram_1_113 : _GEN_2940; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4095 = unuse_way == 2'h1 ? ram_1_114 : _GEN_2941; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4096 = unuse_way == 2'h1 ? ram_1_115 : _GEN_2942; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4097 = unuse_way == 2'h1 ? ram_1_116 : _GEN_2943; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4098 = unuse_way == 2'h1 ? ram_1_117 : _GEN_2944; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4099 = unuse_way == 2'h1 ? ram_1_118 : _GEN_2945; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4100 = unuse_way == 2'h1 ? ram_1_119 : _GEN_2946; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4101 = unuse_way == 2'h1 ? ram_1_120 : _GEN_2947; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4102 = unuse_way == 2'h1 ? ram_1_121 : _GEN_2948; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4103 = unuse_way == 2'h1 ? ram_1_122 : _GEN_2949; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4104 = unuse_way == 2'h1 ? ram_1_123 : _GEN_2950; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4105 = unuse_way == 2'h1 ? ram_1_124 : _GEN_2951; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4106 = unuse_way == 2'h1 ? ram_1_125 : _GEN_2952; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4107 = unuse_way == 2'h1 ? ram_1_126 : _GEN_2953; // @[i_cache.scala 18:24 86:34]
  wire [63:0] _GEN_4108 = unuse_way == 2'h1 ? ram_1_127 : _GEN_2954; // @[i_cache.scala 18:24 86:34]
  wire [31:0] _GEN_4109 = unuse_way == 2'h1 ? tag_1_0 : _GEN_2955; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4110 = unuse_way == 2'h1 ? tag_1_1 : _GEN_2956; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4111 = unuse_way == 2'h1 ? tag_1_2 : _GEN_2957; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4112 = unuse_way == 2'h1 ? tag_1_3 : _GEN_2958; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4113 = unuse_way == 2'h1 ? tag_1_4 : _GEN_2959; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4114 = unuse_way == 2'h1 ? tag_1_5 : _GEN_2960; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4115 = unuse_way == 2'h1 ? tag_1_6 : _GEN_2961; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4116 = unuse_way == 2'h1 ? tag_1_7 : _GEN_2962; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4117 = unuse_way == 2'h1 ? tag_1_8 : _GEN_2963; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4118 = unuse_way == 2'h1 ? tag_1_9 : _GEN_2964; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4119 = unuse_way == 2'h1 ? tag_1_10 : _GEN_2965; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4120 = unuse_way == 2'h1 ? tag_1_11 : _GEN_2966; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4121 = unuse_way == 2'h1 ? tag_1_12 : _GEN_2967; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4122 = unuse_way == 2'h1 ? tag_1_13 : _GEN_2968; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4123 = unuse_way == 2'h1 ? tag_1_14 : _GEN_2969; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4124 = unuse_way == 2'h1 ? tag_1_15 : _GEN_2970; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4125 = unuse_way == 2'h1 ? tag_1_16 : _GEN_2971; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4126 = unuse_way == 2'h1 ? tag_1_17 : _GEN_2972; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4127 = unuse_way == 2'h1 ? tag_1_18 : _GEN_2973; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4128 = unuse_way == 2'h1 ? tag_1_19 : _GEN_2974; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4129 = unuse_way == 2'h1 ? tag_1_20 : _GEN_2975; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4130 = unuse_way == 2'h1 ? tag_1_21 : _GEN_2976; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4131 = unuse_way == 2'h1 ? tag_1_22 : _GEN_2977; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4132 = unuse_way == 2'h1 ? tag_1_23 : _GEN_2978; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4133 = unuse_way == 2'h1 ? tag_1_24 : _GEN_2979; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4134 = unuse_way == 2'h1 ? tag_1_25 : _GEN_2980; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4135 = unuse_way == 2'h1 ? tag_1_26 : _GEN_2981; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4136 = unuse_way == 2'h1 ? tag_1_27 : _GEN_2982; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4137 = unuse_way == 2'h1 ? tag_1_28 : _GEN_2983; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4138 = unuse_way == 2'h1 ? tag_1_29 : _GEN_2984; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4139 = unuse_way == 2'h1 ? tag_1_30 : _GEN_2985; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4140 = unuse_way == 2'h1 ? tag_1_31 : _GEN_2986; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4141 = unuse_way == 2'h1 ? tag_1_32 : _GEN_2987; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4142 = unuse_way == 2'h1 ? tag_1_33 : _GEN_2988; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4143 = unuse_way == 2'h1 ? tag_1_34 : _GEN_2989; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4144 = unuse_way == 2'h1 ? tag_1_35 : _GEN_2990; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4145 = unuse_way == 2'h1 ? tag_1_36 : _GEN_2991; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4146 = unuse_way == 2'h1 ? tag_1_37 : _GEN_2992; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4147 = unuse_way == 2'h1 ? tag_1_38 : _GEN_2993; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4148 = unuse_way == 2'h1 ? tag_1_39 : _GEN_2994; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4149 = unuse_way == 2'h1 ? tag_1_40 : _GEN_2995; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4150 = unuse_way == 2'h1 ? tag_1_41 : _GEN_2996; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4151 = unuse_way == 2'h1 ? tag_1_42 : _GEN_2997; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4152 = unuse_way == 2'h1 ? tag_1_43 : _GEN_2998; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4153 = unuse_way == 2'h1 ? tag_1_44 : _GEN_2999; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4154 = unuse_way == 2'h1 ? tag_1_45 : _GEN_3000; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4155 = unuse_way == 2'h1 ? tag_1_46 : _GEN_3001; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4156 = unuse_way == 2'h1 ? tag_1_47 : _GEN_3002; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4157 = unuse_way == 2'h1 ? tag_1_48 : _GEN_3003; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4158 = unuse_way == 2'h1 ? tag_1_49 : _GEN_3004; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4159 = unuse_way == 2'h1 ? tag_1_50 : _GEN_3005; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4160 = unuse_way == 2'h1 ? tag_1_51 : _GEN_3006; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4161 = unuse_way == 2'h1 ? tag_1_52 : _GEN_3007; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4162 = unuse_way == 2'h1 ? tag_1_53 : _GEN_3008; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4163 = unuse_way == 2'h1 ? tag_1_54 : _GEN_3009; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4164 = unuse_way == 2'h1 ? tag_1_55 : _GEN_3010; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4165 = unuse_way == 2'h1 ? tag_1_56 : _GEN_3011; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4166 = unuse_way == 2'h1 ? tag_1_57 : _GEN_3012; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4167 = unuse_way == 2'h1 ? tag_1_58 : _GEN_3013; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4168 = unuse_way == 2'h1 ? tag_1_59 : _GEN_3014; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4169 = unuse_way == 2'h1 ? tag_1_60 : _GEN_3015; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4170 = unuse_way == 2'h1 ? tag_1_61 : _GEN_3016; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4171 = unuse_way == 2'h1 ? tag_1_62 : _GEN_3017; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4172 = unuse_way == 2'h1 ? tag_1_63 : _GEN_3018; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4173 = unuse_way == 2'h1 ? tag_1_64 : _GEN_3019; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4174 = unuse_way == 2'h1 ? tag_1_65 : _GEN_3020; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4175 = unuse_way == 2'h1 ? tag_1_66 : _GEN_3021; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4176 = unuse_way == 2'h1 ? tag_1_67 : _GEN_3022; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4177 = unuse_way == 2'h1 ? tag_1_68 : _GEN_3023; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4178 = unuse_way == 2'h1 ? tag_1_69 : _GEN_3024; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4179 = unuse_way == 2'h1 ? tag_1_70 : _GEN_3025; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4180 = unuse_way == 2'h1 ? tag_1_71 : _GEN_3026; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4181 = unuse_way == 2'h1 ? tag_1_72 : _GEN_3027; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4182 = unuse_way == 2'h1 ? tag_1_73 : _GEN_3028; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4183 = unuse_way == 2'h1 ? tag_1_74 : _GEN_3029; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4184 = unuse_way == 2'h1 ? tag_1_75 : _GEN_3030; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4185 = unuse_way == 2'h1 ? tag_1_76 : _GEN_3031; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4186 = unuse_way == 2'h1 ? tag_1_77 : _GEN_3032; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4187 = unuse_way == 2'h1 ? tag_1_78 : _GEN_3033; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4188 = unuse_way == 2'h1 ? tag_1_79 : _GEN_3034; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4189 = unuse_way == 2'h1 ? tag_1_80 : _GEN_3035; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4190 = unuse_way == 2'h1 ? tag_1_81 : _GEN_3036; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4191 = unuse_way == 2'h1 ? tag_1_82 : _GEN_3037; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4192 = unuse_way == 2'h1 ? tag_1_83 : _GEN_3038; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4193 = unuse_way == 2'h1 ? tag_1_84 : _GEN_3039; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4194 = unuse_way == 2'h1 ? tag_1_85 : _GEN_3040; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4195 = unuse_way == 2'h1 ? tag_1_86 : _GEN_3041; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4196 = unuse_way == 2'h1 ? tag_1_87 : _GEN_3042; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4197 = unuse_way == 2'h1 ? tag_1_88 : _GEN_3043; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4198 = unuse_way == 2'h1 ? tag_1_89 : _GEN_3044; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4199 = unuse_way == 2'h1 ? tag_1_90 : _GEN_3045; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4200 = unuse_way == 2'h1 ? tag_1_91 : _GEN_3046; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4201 = unuse_way == 2'h1 ? tag_1_92 : _GEN_3047; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4202 = unuse_way == 2'h1 ? tag_1_93 : _GEN_3048; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4203 = unuse_way == 2'h1 ? tag_1_94 : _GEN_3049; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4204 = unuse_way == 2'h1 ? tag_1_95 : _GEN_3050; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4205 = unuse_way == 2'h1 ? tag_1_96 : _GEN_3051; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4206 = unuse_way == 2'h1 ? tag_1_97 : _GEN_3052; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4207 = unuse_way == 2'h1 ? tag_1_98 : _GEN_3053; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4208 = unuse_way == 2'h1 ? tag_1_99 : _GEN_3054; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4209 = unuse_way == 2'h1 ? tag_1_100 : _GEN_3055; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4210 = unuse_way == 2'h1 ? tag_1_101 : _GEN_3056; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4211 = unuse_way == 2'h1 ? tag_1_102 : _GEN_3057; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4212 = unuse_way == 2'h1 ? tag_1_103 : _GEN_3058; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4213 = unuse_way == 2'h1 ? tag_1_104 : _GEN_3059; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4214 = unuse_way == 2'h1 ? tag_1_105 : _GEN_3060; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4215 = unuse_way == 2'h1 ? tag_1_106 : _GEN_3061; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4216 = unuse_way == 2'h1 ? tag_1_107 : _GEN_3062; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4217 = unuse_way == 2'h1 ? tag_1_108 : _GEN_3063; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4218 = unuse_way == 2'h1 ? tag_1_109 : _GEN_3064; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4219 = unuse_way == 2'h1 ? tag_1_110 : _GEN_3065; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4220 = unuse_way == 2'h1 ? tag_1_111 : _GEN_3066; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4221 = unuse_way == 2'h1 ? tag_1_112 : _GEN_3067; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4222 = unuse_way == 2'h1 ? tag_1_113 : _GEN_3068; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4223 = unuse_way == 2'h1 ? tag_1_114 : _GEN_3069; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4224 = unuse_way == 2'h1 ? tag_1_115 : _GEN_3070; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4225 = unuse_way == 2'h1 ? tag_1_116 : _GEN_3071; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4226 = unuse_way == 2'h1 ? tag_1_117 : _GEN_3072; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4227 = unuse_way == 2'h1 ? tag_1_118 : _GEN_3073; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4228 = unuse_way == 2'h1 ? tag_1_119 : _GEN_3074; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4229 = unuse_way == 2'h1 ? tag_1_120 : _GEN_3075; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4230 = unuse_way == 2'h1 ? tag_1_121 : _GEN_3076; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4231 = unuse_way == 2'h1 ? tag_1_122 : _GEN_3077; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4232 = unuse_way == 2'h1 ? tag_1_123 : _GEN_3078; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4233 = unuse_way == 2'h1 ? tag_1_124 : _GEN_3079; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4234 = unuse_way == 2'h1 ? tag_1_125 : _GEN_3080; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4235 = unuse_way == 2'h1 ? tag_1_126 : _GEN_3081; // @[i_cache.scala 20:24 86:34]
  wire [31:0] _GEN_4236 = unuse_way == 2'h1 ? tag_1_127 : _GEN_3082; // @[i_cache.scala 20:24 86:34]
  wire  _GEN_4237 = unuse_way == 2'h1 ? valid_1_0 : _GEN_3083; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4238 = unuse_way == 2'h1 ? valid_1_1 : _GEN_3084; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4239 = unuse_way == 2'h1 ? valid_1_2 : _GEN_3085; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4240 = unuse_way == 2'h1 ? valid_1_3 : _GEN_3086; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4241 = unuse_way == 2'h1 ? valid_1_4 : _GEN_3087; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4242 = unuse_way == 2'h1 ? valid_1_5 : _GEN_3088; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4243 = unuse_way == 2'h1 ? valid_1_6 : _GEN_3089; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4244 = unuse_way == 2'h1 ? valid_1_7 : _GEN_3090; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4245 = unuse_way == 2'h1 ? valid_1_8 : _GEN_3091; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4246 = unuse_way == 2'h1 ? valid_1_9 : _GEN_3092; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4247 = unuse_way == 2'h1 ? valid_1_10 : _GEN_3093; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4248 = unuse_way == 2'h1 ? valid_1_11 : _GEN_3094; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4249 = unuse_way == 2'h1 ? valid_1_12 : _GEN_3095; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4250 = unuse_way == 2'h1 ? valid_1_13 : _GEN_3096; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4251 = unuse_way == 2'h1 ? valid_1_14 : _GEN_3097; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4252 = unuse_way == 2'h1 ? valid_1_15 : _GEN_3098; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4253 = unuse_way == 2'h1 ? valid_1_16 : _GEN_3099; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4254 = unuse_way == 2'h1 ? valid_1_17 : _GEN_3100; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4255 = unuse_way == 2'h1 ? valid_1_18 : _GEN_3101; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4256 = unuse_way == 2'h1 ? valid_1_19 : _GEN_3102; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4257 = unuse_way == 2'h1 ? valid_1_20 : _GEN_3103; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4258 = unuse_way == 2'h1 ? valid_1_21 : _GEN_3104; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4259 = unuse_way == 2'h1 ? valid_1_22 : _GEN_3105; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4260 = unuse_way == 2'h1 ? valid_1_23 : _GEN_3106; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4261 = unuse_way == 2'h1 ? valid_1_24 : _GEN_3107; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4262 = unuse_way == 2'h1 ? valid_1_25 : _GEN_3108; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4263 = unuse_way == 2'h1 ? valid_1_26 : _GEN_3109; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4264 = unuse_way == 2'h1 ? valid_1_27 : _GEN_3110; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4265 = unuse_way == 2'h1 ? valid_1_28 : _GEN_3111; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4266 = unuse_way == 2'h1 ? valid_1_29 : _GEN_3112; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4267 = unuse_way == 2'h1 ? valid_1_30 : _GEN_3113; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4268 = unuse_way == 2'h1 ? valid_1_31 : _GEN_3114; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4269 = unuse_way == 2'h1 ? valid_1_32 : _GEN_3115; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4270 = unuse_way == 2'h1 ? valid_1_33 : _GEN_3116; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4271 = unuse_way == 2'h1 ? valid_1_34 : _GEN_3117; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4272 = unuse_way == 2'h1 ? valid_1_35 : _GEN_3118; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4273 = unuse_way == 2'h1 ? valid_1_36 : _GEN_3119; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4274 = unuse_way == 2'h1 ? valid_1_37 : _GEN_3120; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4275 = unuse_way == 2'h1 ? valid_1_38 : _GEN_3121; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4276 = unuse_way == 2'h1 ? valid_1_39 : _GEN_3122; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4277 = unuse_way == 2'h1 ? valid_1_40 : _GEN_3123; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4278 = unuse_way == 2'h1 ? valid_1_41 : _GEN_3124; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4279 = unuse_way == 2'h1 ? valid_1_42 : _GEN_3125; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4280 = unuse_way == 2'h1 ? valid_1_43 : _GEN_3126; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4281 = unuse_way == 2'h1 ? valid_1_44 : _GEN_3127; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4282 = unuse_way == 2'h1 ? valid_1_45 : _GEN_3128; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4283 = unuse_way == 2'h1 ? valid_1_46 : _GEN_3129; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4284 = unuse_way == 2'h1 ? valid_1_47 : _GEN_3130; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4285 = unuse_way == 2'h1 ? valid_1_48 : _GEN_3131; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4286 = unuse_way == 2'h1 ? valid_1_49 : _GEN_3132; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4287 = unuse_way == 2'h1 ? valid_1_50 : _GEN_3133; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4288 = unuse_way == 2'h1 ? valid_1_51 : _GEN_3134; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4289 = unuse_way == 2'h1 ? valid_1_52 : _GEN_3135; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4290 = unuse_way == 2'h1 ? valid_1_53 : _GEN_3136; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4291 = unuse_way == 2'h1 ? valid_1_54 : _GEN_3137; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4292 = unuse_way == 2'h1 ? valid_1_55 : _GEN_3138; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4293 = unuse_way == 2'h1 ? valid_1_56 : _GEN_3139; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4294 = unuse_way == 2'h1 ? valid_1_57 : _GEN_3140; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4295 = unuse_way == 2'h1 ? valid_1_58 : _GEN_3141; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4296 = unuse_way == 2'h1 ? valid_1_59 : _GEN_3142; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4297 = unuse_way == 2'h1 ? valid_1_60 : _GEN_3143; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4298 = unuse_way == 2'h1 ? valid_1_61 : _GEN_3144; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4299 = unuse_way == 2'h1 ? valid_1_62 : _GEN_3145; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4300 = unuse_way == 2'h1 ? valid_1_63 : _GEN_3146; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4301 = unuse_way == 2'h1 ? valid_1_64 : _GEN_3147; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4302 = unuse_way == 2'h1 ? valid_1_65 : _GEN_3148; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4303 = unuse_way == 2'h1 ? valid_1_66 : _GEN_3149; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4304 = unuse_way == 2'h1 ? valid_1_67 : _GEN_3150; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4305 = unuse_way == 2'h1 ? valid_1_68 : _GEN_3151; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4306 = unuse_way == 2'h1 ? valid_1_69 : _GEN_3152; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4307 = unuse_way == 2'h1 ? valid_1_70 : _GEN_3153; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4308 = unuse_way == 2'h1 ? valid_1_71 : _GEN_3154; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4309 = unuse_way == 2'h1 ? valid_1_72 : _GEN_3155; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4310 = unuse_way == 2'h1 ? valid_1_73 : _GEN_3156; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4311 = unuse_way == 2'h1 ? valid_1_74 : _GEN_3157; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4312 = unuse_way == 2'h1 ? valid_1_75 : _GEN_3158; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4313 = unuse_way == 2'h1 ? valid_1_76 : _GEN_3159; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4314 = unuse_way == 2'h1 ? valid_1_77 : _GEN_3160; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4315 = unuse_way == 2'h1 ? valid_1_78 : _GEN_3161; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4316 = unuse_way == 2'h1 ? valid_1_79 : _GEN_3162; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4317 = unuse_way == 2'h1 ? valid_1_80 : _GEN_3163; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4318 = unuse_way == 2'h1 ? valid_1_81 : _GEN_3164; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4319 = unuse_way == 2'h1 ? valid_1_82 : _GEN_3165; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4320 = unuse_way == 2'h1 ? valid_1_83 : _GEN_3166; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4321 = unuse_way == 2'h1 ? valid_1_84 : _GEN_3167; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4322 = unuse_way == 2'h1 ? valid_1_85 : _GEN_3168; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4323 = unuse_way == 2'h1 ? valid_1_86 : _GEN_3169; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4324 = unuse_way == 2'h1 ? valid_1_87 : _GEN_3170; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4325 = unuse_way == 2'h1 ? valid_1_88 : _GEN_3171; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4326 = unuse_way == 2'h1 ? valid_1_89 : _GEN_3172; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4327 = unuse_way == 2'h1 ? valid_1_90 : _GEN_3173; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4328 = unuse_way == 2'h1 ? valid_1_91 : _GEN_3174; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4329 = unuse_way == 2'h1 ? valid_1_92 : _GEN_3175; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4330 = unuse_way == 2'h1 ? valid_1_93 : _GEN_3176; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4331 = unuse_way == 2'h1 ? valid_1_94 : _GEN_3177; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4332 = unuse_way == 2'h1 ? valid_1_95 : _GEN_3178; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4333 = unuse_way == 2'h1 ? valid_1_96 : _GEN_3179; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4334 = unuse_way == 2'h1 ? valid_1_97 : _GEN_3180; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4335 = unuse_way == 2'h1 ? valid_1_98 : _GEN_3181; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4336 = unuse_way == 2'h1 ? valid_1_99 : _GEN_3182; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4337 = unuse_way == 2'h1 ? valid_1_100 : _GEN_3183; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4338 = unuse_way == 2'h1 ? valid_1_101 : _GEN_3184; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4339 = unuse_way == 2'h1 ? valid_1_102 : _GEN_3185; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4340 = unuse_way == 2'h1 ? valid_1_103 : _GEN_3186; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4341 = unuse_way == 2'h1 ? valid_1_104 : _GEN_3187; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4342 = unuse_way == 2'h1 ? valid_1_105 : _GEN_3188; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4343 = unuse_way == 2'h1 ? valid_1_106 : _GEN_3189; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4344 = unuse_way == 2'h1 ? valid_1_107 : _GEN_3190; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4345 = unuse_way == 2'h1 ? valid_1_108 : _GEN_3191; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4346 = unuse_way == 2'h1 ? valid_1_109 : _GEN_3192; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4347 = unuse_way == 2'h1 ? valid_1_110 : _GEN_3193; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4348 = unuse_way == 2'h1 ? valid_1_111 : _GEN_3194; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4349 = unuse_way == 2'h1 ? valid_1_112 : _GEN_3195; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4350 = unuse_way == 2'h1 ? valid_1_113 : _GEN_3196; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4351 = unuse_way == 2'h1 ? valid_1_114 : _GEN_3197; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4352 = unuse_way == 2'h1 ? valid_1_115 : _GEN_3198; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4353 = unuse_way == 2'h1 ? valid_1_116 : _GEN_3199; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4354 = unuse_way == 2'h1 ? valid_1_117 : _GEN_3200; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4355 = unuse_way == 2'h1 ? valid_1_118 : _GEN_3201; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4356 = unuse_way == 2'h1 ? valid_1_119 : _GEN_3202; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4357 = unuse_way == 2'h1 ? valid_1_120 : _GEN_3203; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4358 = unuse_way == 2'h1 ? valid_1_121 : _GEN_3204; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4359 = unuse_way == 2'h1 ? valid_1_122 : _GEN_3205; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4360 = unuse_way == 2'h1 ? valid_1_123 : _GEN_3206; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4361 = unuse_way == 2'h1 ? valid_1_124 : _GEN_3207; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4362 = unuse_way == 2'h1 ? valid_1_125 : _GEN_3208; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4363 = unuse_way == 2'h1 ? valid_1_126 : _GEN_3209; // @[i_cache.scala 22:26 86:34]
  wire  _GEN_4364 = unuse_way == 2'h1 ? valid_1_127 : _GEN_3210; // @[i_cache.scala 22:26 86:34]
  wire [2:0] _GEN_4365 = 3'h4 == state ? 3'h1 : state; // @[i_cache.scala 55:18 111:19 53:24]
  wire [2:0] _GEN_4366 = 3'h3 == state ? 3'h4 : _GEN_4365; // @[i_cache.scala 55:18 85:19]
  wire [63:0] _GEN_4367 = 3'h3 == state ? _GEN_3596 : ram_0_0; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4368 = 3'h3 == state ? _GEN_3597 : ram_0_1; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4369 = 3'h3 == state ? _GEN_3598 : ram_0_2; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4370 = 3'h3 == state ? _GEN_3599 : ram_0_3; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4371 = 3'h3 == state ? _GEN_3600 : ram_0_4; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4372 = 3'h3 == state ? _GEN_3601 : ram_0_5; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4373 = 3'h3 == state ? _GEN_3602 : ram_0_6; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4374 = 3'h3 == state ? _GEN_3603 : ram_0_7; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4375 = 3'h3 == state ? _GEN_3604 : ram_0_8; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4376 = 3'h3 == state ? _GEN_3605 : ram_0_9; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4377 = 3'h3 == state ? _GEN_3606 : ram_0_10; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4378 = 3'h3 == state ? _GEN_3607 : ram_0_11; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4379 = 3'h3 == state ? _GEN_3608 : ram_0_12; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4380 = 3'h3 == state ? _GEN_3609 : ram_0_13; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4381 = 3'h3 == state ? _GEN_3610 : ram_0_14; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4382 = 3'h3 == state ? _GEN_3611 : ram_0_15; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4383 = 3'h3 == state ? _GEN_3612 : ram_0_16; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4384 = 3'h3 == state ? _GEN_3613 : ram_0_17; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4385 = 3'h3 == state ? _GEN_3614 : ram_0_18; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4386 = 3'h3 == state ? _GEN_3615 : ram_0_19; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4387 = 3'h3 == state ? _GEN_3616 : ram_0_20; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4388 = 3'h3 == state ? _GEN_3617 : ram_0_21; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4389 = 3'h3 == state ? _GEN_3618 : ram_0_22; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4390 = 3'h3 == state ? _GEN_3619 : ram_0_23; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4391 = 3'h3 == state ? _GEN_3620 : ram_0_24; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4392 = 3'h3 == state ? _GEN_3621 : ram_0_25; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4393 = 3'h3 == state ? _GEN_3622 : ram_0_26; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4394 = 3'h3 == state ? _GEN_3623 : ram_0_27; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4395 = 3'h3 == state ? _GEN_3624 : ram_0_28; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4396 = 3'h3 == state ? _GEN_3625 : ram_0_29; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4397 = 3'h3 == state ? _GEN_3626 : ram_0_30; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4398 = 3'h3 == state ? _GEN_3627 : ram_0_31; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4399 = 3'h3 == state ? _GEN_3628 : ram_0_32; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4400 = 3'h3 == state ? _GEN_3629 : ram_0_33; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4401 = 3'h3 == state ? _GEN_3630 : ram_0_34; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4402 = 3'h3 == state ? _GEN_3631 : ram_0_35; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4403 = 3'h3 == state ? _GEN_3632 : ram_0_36; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4404 = 3'h3 == state ? _GEN_3633 : ram_0_37; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4405 = 3'h3 == state ? _GEN_3634 : ram_0_38; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4406 = 3'h3 == state ? _GEN_3635 : ram_0_39; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4407 = 3'h3 == state ? _GEN_3636 : ram_0_40; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4408 = 3'h3 == state ? _GEN_3637 : ram_0_41; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4409 = 3'h3 == state ? _GEN_3638 : ram_0_42; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4410 = 3'h3 == state ? _GEN_3639 : ram_0_43; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4411 = 3'h3 == state ? _GEN_3640 : ram_0_44; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4412 = 3'h3 == state ? _GEN_3641 : ram_0_45; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4413 = 3'h3 == state ? _GEN_3642 : ram_0_46; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4414 = 3'h3 == state ? _GEN_3643 : ram_0_47; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4415 = 3'h3 == state ? _GEN_3644 : ram_0_48; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4416 = 3'h3 == state ? _GEN_3645 : ram_0_49; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4417 = 3'h3 == state ? _GEN_3646 : ram_0_50; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4418 = 3'h3 == state ? _GEN_3647 : ram_0_51; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4419 = 3'h3 == state ? _GEN_3648 : ram_0_52; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4420 = 3'h3 == state ? _GEN_3649 : ram_0_53; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4421 = 3'h3 == state ? _GEN_3650 : ram_0_54; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4422 = 3'h3 == state ? _GEN_3651 : ram_0_55; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4423 = 3'h3 == state ? _GEN_3652 : ram_0_56; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4424 = 3'h3 == state ? _GEN_3653 : ram_0_57; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4425 = 3'h3 == state ? _GEN_3654 : ram_0_58; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4426 = 3'h3 == state ? _GEN_3655 : ram_0_59; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4427 = 3'h3 == state ? _GEN_3656 : ram_0_60; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4428 = 3'h3 == state ? _GEN_3657 : ram_0_61; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4429 = 3'h3 == state ? _GEN_3658 : ram_0_62; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4430 = 3'h3 == state ? _GEN_3659 : ram_0_63; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4431 = 3'h3 == state ? _GEN_3660 : ram_0_64; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4432 = 3'h3 == state ? _GEN_3661 : ram_0_65; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4433 = 3'h3 == state ? _GEN_3662 : ram_0_66; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4434 = 3'h3 == state ? _GEN_3663 : ram_0_67; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4435 = 3'h3 == state ? _GEN_3664 : ram_0_68; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4436 = 3'h3 == state ? _GEN_3665 : ram_0_69; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4437 = 3'h3 == state ? _GEN_3666 : ram_0_70; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4438 = 3'h3 == state ? _GEN_3667 : ram_0_71; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4439 = 3'h3 == state ? _GEN_3668 : ram_0_72; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4440 = 3'h3 == state ? _GEN_3669 : ram_0_73; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4441 = 3'h3 == state ? _GEN_3670 : ram_0_74; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4442 = 3'h3 == state ? _GEN_3671 : ram_0_75; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4443 = 3'h3 == state ? _GEN_3672 : ram_0_76; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4444 = 3'h3 == state ? _GEN_3673 : ram_0_77; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4445 = 3'h3 == state ? _GEN_3674 : ram_0_78; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4446 = 3'h3 == state ? _GEN_3675 : ram_0_79; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4447 = 3'h3 == state ? _GEN_3676 : ram_0_80; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4448 = 3'h3 == state ? _GEN_3677 : ram_0_81; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4449 = 3'h3 == state ? _GEN_3678 : ram_0_82; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4450 = 3'h3 == state ? _GEN_3679 : ram_0_83; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4451 = 3'h3 == state ? _GEN_3680 : ram_0_84; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4452 = 3'h3 == state ? _GEN_3681 : ram_0_85; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4453 = 3'h3 == state ? _GEN_3682 : ram_0_86; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4454 = 3'h3 == state ? _GEN_3683 : ram_0_87; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4455 = 3'h3 == state ? _GEN_3684 : ram_0_88; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4456 = 3'h3 == state ? _GEN_3685 : ram_0_89; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4457 = 3'h3 == state ? _GEN_3686 : ram_0_90; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4458 = 3'h3 == state ? _GEN_3687 : ram_0_91; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4459 = 3'h3 == state ? _GEN_3688 : ram_0_92; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4460 = 3'h3 == state ? _GEN_3689 : ram_0_93; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4461 = 3'h3 == state ? _GEN_3690 : ram_0_94; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4462 = 3'h3 == state ? _GEN_3691 : ram_0_95; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4463 = 3'h3 == state ? _GEN_3692 : ram_0_96; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4464 = 3'h3 == state ? _GEN_3693 : ram_0_97; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4465 = 3'h3 == state ? _GEN_3694 : ram_0_98; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4466 = 3'h3 == state ? _GEN_3695 : ram_0_99; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4467 = 3'h3 == state ? _GEN_3696 : ram_0_100; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4468 = 3'h3 == state ? _GEN_3697 : ram_0_101; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4469 = 3'h3 == state ? _GEN_3698 : ram_0_102; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4470 = 3'h3 == state ? _GEN_3699 : ram_0_103; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4471 = 3'h3 == state ? _GEN_3700 : ram_0_104; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4472 = 3'h3 == state ? _GEN_3701 : ram_0_105; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4473 = 3'h3 == state ? _GEN_3702 : ram_0_106; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4474 = 3'h3 == state ? _GEN_3703 : ram_0_107; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4475 = 3'h3 == state ? _GEN_3704 : ram_0_108; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4476 = 3'h3 == state ? _GEN_3705 : ram_0_109; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4477 = 3'h3 == state ? _GEN_3706 : ram_0_110; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4478 = 3'h3 == state ? _GEN_3707 : ram_0_111; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4479 = 3'h3 == state ? _GEN_3708 : ram_0_112; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4480 = 3'h3 == state ? _GEN_3709 : ram_0_113; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4481 = 3'h3 == state ? _GEN_3710 : ram_0_114; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4482 = 3'h3 == state ? _GEN_3711 : ram_0_115; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4483 = 3'h3 == state ? _GEN_3712 : ram_0_116; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4484 = 3'h3 == state ? _GEN_3713 : ram_0_117; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4485 = 3'h3 == state ? _GEN_3714 : ram_0_118; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4486 = 3'h3 == state ? _GEN_3715 : ram_0_119; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4487 = 3'h3 == state ? _GEN_3716 : ram_0_120; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4488 = 3'h3 == state ? _GEN_3717 : ram_0_121; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4489 = 3'h3 == state ? _GEN_3718 : ram_0_122; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4490 = 3'h3 == state ? _GEN_3719 : ram_0_123; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4491 = 3'h3 == state ? _GEN_3720 : ram_0_124; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4492 = 3'h3 == state ? _GEN_3721 : ram_0_125; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4493 = 3'h3 == state ? _GEN_3722 : ram_0_126; // @[i_cache.scala 55:18 17:24]
  wire [63:0] _GEN_4494 = 3'h3 == state ? _GEN_3723 : ram_0_127; // @[i_cache.scala 55:18 17:24]
  wire [31:0] _GEN_4495 = 3'h3 == state ? _GEN_3724 : tag_0_0; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4496 = 3'h3 == state ? _GEN_3725 : tag_0_1; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4497 = 3'h3 == state ? _GEN_3726 : tag_0_2; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4498 = 3'h3 == state ? _GEN_3727 : tag_0_3; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4499 = 3'h3 == state ? _GEN_3728 : tag_0_4; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4500 = 3'h3 == state ? _GEN_3729 : tag_0_5; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4501 = 3'h3 == state ? _GEN_3730 : tag_0_6; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4502 = 3'h3 == state ? _GEN_3731 : tag_0_7; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4503 = 3'h3 == state ? _GEN_3732 : tag_0_8; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4504 = 3'h3 == state ? _GEN_3733 : tag_0_9; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4505 = 3'h3 == state ? _GEN_3734 : tag_0_10; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4506 = 3'h3 == state ? _GEN_3735 : tag_0_11; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4507 = 3'h3 == state ? _GEN_3736 : tag_0_12; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4508 = 3'h3 == state ? _GEN_3737 : tag_0_13; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4509 = 3'h3 == state ? _GEN_3738 : tag_0_14; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4510 = 3'h3 == state ? _GEN_3739 : tag_0_15; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4511 = 3'h3 == state ? _GEN_3740 : tag_0_16; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4512 = 3'h3 == state ? _GEN_3741 : tag_0_17; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4513 = 3'h3 == state ? _GEN_3742 : tag_0_18; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4514 = 3'h3 == state ? _GEN_3743 : tag_0_19; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4515 = 3'h3 == state ? _GEN_3744 : tag_0_20; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4516 = 3'h3 == state ? _GEN_3745 : tag_0_21; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4517 = 3'h3 == state ? _GEN_3746 : tag_0_22; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4518 = 3'h3 == state ? _GEN_3747 : tag_0_23; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4519 = 3'h3 == state ? _GEN_3748 : tag_0_24; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4520 = 3'h3 == state ? _GEN_3749 : tag_0_25; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4521 = 3'h3 == state ? _GEN_3750 : tag_0_26; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4522 = 3'h3 == state ? _GEN_3751 : tag_0_27; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4523 = 3'h3 == state ? _GEN_3752 : tag_0_28; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4524 = 3'h3 == state ? _GEN_3753 : tag_0_29; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4525 = 3'h3 == state ? _GEN_3754 : tag_0_30; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4526 = 3'h3 == state ? _GEN_3755 : tag_0_31; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4527 = 3'h3 == state ? _GEN_3756 : tag_0_32; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4528 = 3'h3 == state ? _GEN_3757 : tag_0_33; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4529 = 3'h3 == state ? _GEN_3758 : tag_0_34; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4530 = 3'h3 == state ? _GEN_3759 : tag_0_35; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4531 = 3'h3 == state ? _GEN_3760 : tag_0_36; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4532 = 3'h3 == state ? _GEN_3761 : tag_0_37; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4533 = 3'h3 == state ? _GEN_3762 : tag_0_38; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4534 = 3'h3 == state ? _GEN_3763 : tag_0_39; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4535 = 3'h3 == state ? _GEN_3764 : tag_0_40; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4536 = 3'h3 == state ? _GEN_3765 : tag_0_41; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4537 = 3'h3 == state ? _GEN_3766 : tag_0_42; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4538 = 3'h3 == state ? _GEN_3767 : tag_0_43; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4539 = 3'h3 == state ? _GEN_3768 : tag_0_44; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4540 = 3'h3 == state ? _GEN_3769 : tag_0_45; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4541 = 3'h3 == state ? _GEN_3770 : tag_0_46; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4542 = 3'h3 == state ? _GEN_3771 : tag_0_47; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4543 = 3'h3 == state ? _GEN_3772 : tag_0_48; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4544 = 3'h3 == state ? _GEN_3773 : tag_0_49; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4545 = 3'h3 == state ? _GEN_3774 : tag_0_50; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4546 = 3'h3 == state ? _GEN_3775 : tag_0_51; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4547 = 3'h3 == state ? _GEN_3776 : tag_0_52; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4548 = 3'h3 == state ? _GEN_3777 : tag_0_53; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4549 = 3'h3 == state ? _GEN_3778 : tag_0_54; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4550 = 3'h3 == state ? _GEN_3779 : tag_0_55; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4551 = 3'h3 == state ? _GEN_3780 : tag_0_56; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4552 = 3'h3 == state ? _GEN_3781 : tag_0_57; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4553 = 3'h3 == state ? _GEN_3782 : tag_0_58; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4554 = 3'h3 == state ? _GEN_3783 : tag_0_59; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4555 = 3'h3 == state ? _GEN_3784 : tag_0_60; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4556 = 3'h3 == state ? _GEN_3785 : tag_0_61; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4557 = 3'h3 == state ? _GEN_3786 : tag_0_62; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4558 = 3'h3 == state ? _GEN_3787 : tag_0_63; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4559 = 3'h3 == state ? _GEN_3788 : tag_0_64; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4560 = 3'h3 == state ? _GEN_3789 : tag_0_65; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4561 = 3'h3 == state ? _GEN_3790 : tag_0_66; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4562 = 3'h3 == state ? _GEN_3791 : tag_0_67; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4563 = 3'h3 == state ? _GEN_3792 : tag_0_68; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4564 = 3'h3 == state ? _GEN_3793 : tag_0_69; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4565 = 3'h3 == state ? _GEN_3794 : tag_0_70; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4566 = 3'h3 == state ? _GEN_3795 : tag_0_71; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4567 = 3'h3 == state ? _GEN_3796 : tag_0_72; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4568 = 3'h3 == state ? _GEN_3797 : tag_0_73; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4569 = 3'h3 == state ? _GEN_3798 : tag_0_74; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4570 = 3'h3 == state ? _GEN_3799 : tag_0_75; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4571 = 3'h3 == state ? _GEN_3800 : tag_0_76; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4572 = 3'h3 == state ? _GEN_3801 : tag_0_77; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4573 = 3'h3 == state ? _GEN_3802 : tag_0_78; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4574 = 3'h3 == state ? _GEN_3803 : tag_0_79; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4575 = 3'h3 == state ? _GEN_3804 : tag_0_80; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4576 = 3'h3 == state ? _GEN_3805 : tag_0_81; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4577 = 3'h3 == state ? _GEN_3806 : tag_0_82; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4578 = 3'h3 == state ? _GEN_3807 : tag_0_83; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4579 = 3'h3 == state ? _GEN_3808 : tag_0_84; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4580 = 3'h3 == state ? _GEN_3809 : tag_0_85; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4581 = 3'h3 == state ? _GEN_3810 : tag_0_86; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4582 = 3'h3 == state ? _GEN_3811 : tag_0_87; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4583 = 3'h3 == state ? _GEN_3812 : tag_0_88; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4584 = 3'h3 == state ? _GEN_3813 : tag_0_89; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4585 = 3'h3 == state ? _GEN_3814 : tag_0_90; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4586 = 3'h3 == state ? _GEN_3815 : tag_0_91; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4587 = 3'h3 == state ? _GEN_3816 : tag_0_92; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4588 = 3'h3 == state ? _GEN_3817 : tag_0_93; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4589 = 3'h3 == state ? _GEN_3818 : tag_0_94; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4590 = 3'h3 == state ? _GEN_3819 : tag_0_95; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4591 = 3'h3 == state ? _GEN_3820 : tag_0_96; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4592 = 3'h3 == state ? _GEN_3821 : tag_0_97; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4593 = 3'h3 == state ? _GEN_3822 : tag_0_98; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4594 = 3'h3 == state ? _GEN_3823 : tag_0_99; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4595 = 3'h3 == state ? _GEN_3824 : tag_0_100; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4596 = 3'h3 == state ? _GEN_3825 : tag_0_101; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4597 = 3'h3 == state ? _GEN_3826 : tag_0_102; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4598 = 3'h3 == state ? _GEN_3827 : tag_0_103; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4599 = 3'h3 == state ? _GEN_3828 : tag_0_104; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4600 = 3'h3 == state ? _GEN_3829 : tag_0_105; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4601 = 3'h3 == state ? _GEN_3830 : tag_0_106; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4602 = 3'h3 == state ? _GEN_3831 : tag_0_107; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4603 = 3'h3 == state ? _GEN_3832 : tag_0_108; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4604 = 3'h3 == state ? _GEN_3833 : tag_0_109; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4605 = 3'h3 == state ? _GEN_3834 : tag_0_110; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4606 = 3'h3 == state ? _GEN_3835 : tag_0_111; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4607 = 3'h3 == state ? _GEN_3836 : tag_0_112; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4608 = 3'h3 == state ? _GEN_3837 : tag_0_113; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4609 = 3'h3 == state ? _GEN_3838 : tag_0_114; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4610 = 3'h3 == state ? _GEN_3839 : tag_0_115; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4611 = 3'h3 == state ? _GEN_3840 : tag_0_116; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4612 = 3'h3 == state ? _GEN_3841 : tag_0_117; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4613 = 3'h3 == state ? _GEN_3842 : tag_0_118; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4614 = 3'h3 == state ? _GEN_3843 : tag_0_119; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4615 = 3'h3 == state ? _GEN_3844 : tag_0_120; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4616 = 3'h3 == state ? _GEN_3845 : tag_0_121; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4617 = 3'h3 == state ? _GEN_3846 : tag_0_122; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4618 = 3'h3 == state ? _GEN_3847 : tag_0_123; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4619 = 3'h3 == state ? _GEN_3848 : tag_0_124; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4620 = 3'h3 == state ? _GEN_3849 : tag_0_125; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4621 = 3'h3 == state ? _GEN_3850 : tag_0_126; // @[i_cache.scala 55:18 19:24]
  wire [31:0] _GEN_4622 = 3'h3 == state ? _GEN_3851 : tag_0_127; // @[i_cache.scala 55:18 19:24]
  wire  _GEN_4623 = 3'h3 == state ? _GEN_3852 : valid_0_0; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4624 = 3'h3 == state ? _GEN_3853 : valid_0_1; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4625 = 3'h3 == state ? _GEN_3854 : valid_0_2; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4626 = 3'h3 == state ? _GEN_3855 : valid_0_3; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4627 = 3'h3 == state ? _GEN_3856 : valid_0_4; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4628 = 3'h3 == state ? _GEN_3857 : valid_0_5; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4629 = 3'h3 == state ? _GEN_3858 : valid_0_6; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4630 = 3'h3 == state ? _GEN_3859 : valid_0_7; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4631 = 3'h3 == state ? _GEN_3860 : valid_0_8; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4632 = 3'h3 == state ? _GEN_3861 : valid_0_9; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4633 = 3'h3 == state ? _GEN_3862 : valid_0_10; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4634 = 3'h3 == state ? _GEN_3863 : valid_0_11; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4635 = 3'h3 == state ? _GEN_3864 : valid_0_12; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4636 = 3'h3 == state ? _GEN_3865 : valid_0_13; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4637 = 3'h3 == state ? _GEN_3866 : valid_0_14; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4638 = 3'h3 == state ? _GEN_3867 : valid_0_15; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4639 = 3'h3 == state ? _GEN_3868 : valid_0_16; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4640 = 3'h3 == state ? _GEN_3869 : valid_0_17; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4641 = 3'h3 == state ? _GEN_3870 : valid_0_18; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4642 = 3'h3 == state ? _GEN_3871 : valid_0_19; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4643 = 3'h3 == state ? _GEN_3872 : valid_0_20; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4644 = 3'h3 == state ? _GEN_3873 : valid_0_21; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4645 = 3'h3 == state ? _GEN_3874 : valid_0_22; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4646 = 3'h3 == state ? _GEN_3875 : valid_0_23; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4647 = 3'h3 == state ? _GEN_3876 : valid_0_24; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4648 = 3'h3 == state ? _GEN_3877 : valid_0_25; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4649 = 3'h3 == state ? _GEN_3878 : valid_0_26; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4650 = 3'h3 == state ? _GEN_3879 : valid_0_27; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4651 = 3'h3 == state ? _GEN_3880 : valid_0_28; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4652 = 3'h3 == state ? _GEN_3881 : valid_0_29; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4653 = 3'h3 == state ? _GEN_3882 : valid_0_30; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4654 = 3'h3 == state ? _GEN_3883 : valid_0_31; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4655 = 3'h3 == state ? _GEN_3884 : valid_0_32; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4656 = 3'h3 == state ? _GEN_3885 : valid_0_33; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4657 = 3'h3 == state ? _GEN_3886 : valid_0_34; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4658 = 3'h3 == state ? _GEN_3887 : valid_0_35; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4659 = 3'h3 == state ? _GEN_3888 : valid_0_36; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4660 = 3'h3 == state ? _GEN_3889 : valid_0_37; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4661 = 3'h3 == state ? _GEN_3890 : valid_0_38; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4662 = 3'h3 == state ? _GEN_3891 : valid_0_39; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4663 = 3'h3 == state ? _GEN_3892 : valid_0_40; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4664 = 3'h3 == state ? _GEN_3893 : valid_0_41; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4665 = 3'h3 == state ? _GEN_3894 : valid_0_42; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4666 = 3'h3 == state ? _GEN_3895 : valid_0_43; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4667 = 3'h3 == state ? _GEN_3896 : valid_0_44; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4668 = 3'h3 == state ? _GEN_3897 : valid_0_45; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4669 = 3'h3 == state ? _GEN_3898 : valid_0_46; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4670 = 3'h3 == state ? _GEN_3899 : valid_0_47; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4671 = 3'h3 == state ? _GEN_3900 : valid_0_48; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4672 = 3'h3 == state ? _GEN_3901 : valid_0_49; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4673 = 3'h3 == state ? _GEN_3902 : valid_0_50; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4674 = 3'h3 == state ? _GEN_3903 : valid_0_51; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4675 = 3'h3 == state ? _GEN_3904 : valid_0_52; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4676 = 3'h3 == state ? _GEN_3905 : valid_0_53; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4677 = 3'h3 == state ? _GEN_3906 : valid_0_54; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4678 = 3'h3 == state ? _GEN_3907 : valid_0_55; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4679 = 3'h3 == state ? _GEN_3908 : valid_0_56; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4680 = 3'h3 == state ? _GEN_3909 : valid_0_57; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4681 = 3'h3 == state ? _GEN_3910 : valid_0_58; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4682 = 3'h3 == state ? _GEN_3911 : valid_0_59; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4683 = 3'h3 == state ? _GEN_3912 : valid_0_60; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4684 = 3'h3 == state ? _GEN_3913 : valid_0_61; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4685 = 3'h3 == state ? _GEN_3914 : valid_0_62; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4686 = 3'h3 == state ? _GEN_3915 : valid_0_63; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4687 = 3'h3 == state ? _GEN_3916 : valid_0_64; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4688 = 3'h3 == state ? _GEN_3917 : valid_0_65; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4689 = 3'h3 == state ? _GEN_3918 : valid_0_66; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4690 = 3'h3 == state ? _GEN_3919 : valid_0_67; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4691 = 3'h3 == state ? _GEN_3920 : valid_0_68; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4692 = 3'h3 == state ? _GEN_3921 : valid_0_69; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4693 = 3'h3 == state ? _GEN_3922 : valid_0_70; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4694 = 3'h3 == state ? _GEN_3923 : valid_0_71; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4695 = 3'h3 == state ? _GEN_3924 : valid_0_72; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4696 = 3'h3 == state ? _GEN_3925 : valid_0_73; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4697 = 3'h3 == state ? _GEN_3926 : valid_0_74; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4698 = 3'h3 == state ? _GEN_3927 : valid_0_75; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4699 = 3'h3 == state ? _GEN_3928 : valid_0_76; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4700 = 3'h3 == state ? _GEN_3929 : valid_0_77; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4701 = 3'h3 == state ? _GEN_3930 : valid_0_78; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4702 = 3'h3 == state ? _GEN_3931 : valid_0_79; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4703 = 3'h3 == state ? _GEN_3932 : valid_0_80; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4704 = 3'h3 == state ? _GEN_3933 : valid_0_81; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4705 = 3'h3 == state ? _GEN_3934 : valid_0_82; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4706 = 3'h3 == state ? _GEN_3935 : valid_0_83; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4707 = 3'h3 == state ? _GEN_3936 : valid_0_84; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4708 = 3'h3 == state ? _GEN_3937 : valid_0_85; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4709 = 3'h3 == state ? _GEN_3938 : valid_0_86; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4710 = 3'h3 == state ? _GEN_3939 : valid_0_87; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4711 = 3'h3 == state ? _GEN_3940 : valid_0_88; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4712 = 3'h3 == state ? _GEN_3941 : valid_0_89; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4713 = 3'h3 == state ? _GEN_3942 : valid_0_90; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4714 = 3'h3 == state ? _GEN_3943 : valid_0_91; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4715 = 3'h3 == state ? _GEN_3944 : valid_0_92; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4716 = 3'h3 == state ? _GEN_3945 : valid_0_93; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4717 = 3'h3 == state ? _GEN_3946 : valid_0_94; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4718 = 3'h3 == state ? _GEN_3947 : valid_0_95; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4719 = 3'h3 == state ? _GEN_3948 : valid_0_96; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4720 = 3'h3 == state ? _GEN_3949 : valid_0_97; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4721 = 3'h3 == state ? _GEN_3950 : valid_0_98; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4722 = 3'h3 == state ? _GEN_3951 : valid_0_99; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4723 = 3'h3 == state ? _GEN_3952 : valid_0_100; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4724 = 3'h3 == state ? _GEN_3953 : valid_0_101; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4725 = 3'h3 == state ? _GEN_3954 : valid_0_102; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4726 = 3'h3 == state ? _GEN_3955 : valid_0_103; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4727 = 3'h3 == state ? _GEN_3956 : valid_0_104; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4728 = 3'h3 == state ? _GEN_3957 : valid_0_105; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4729 = 3'h3 == state ? _GEN_3958 : valid_0_106; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4730 = 3'h3 == state ? _GEN_3959 : valid_0_107; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4731 = 3'h3 == state ? _GEN_3960 : valid_0_108; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4732 = 3'h3 == state ? _GEN_3961 : valid_0_109; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4733 = 3'h3 == state ? _GEN_3962 : valid_0_110; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4734 = 3'h3 == state ? _GEN_3963 : valid_0_111; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4735 = 3'h3 == state ? _GEN_3964 : valid_0_112; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4736 = 3'h3 == state ? _GEN_3965 : valid_0_113; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4737 = 3'h3 == state ? _GEN_3966 : valid_0_114; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4738 = 3'h3 == state ? _GEN_3967 : valid_0_115; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4739 = 3'h3 == state ? _GEN_3968 : valid_0_116; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4740 = 3'h3 == state ? _GEN_3969 : valid_0_117; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4741 = 3'h3 == state ? _GEN_3970 : valid_0_118; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4742 = 3'h3 == state ? _GEN_3971 : valid_0_119; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4743 = 3'h3 == state ? _GEN_3972 : valid_0_120; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4744 = 3'h3 == state ? _GEN_3973 : valid_0_121; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4745 = 3'h3 == state ? _GEN_3974 : valid_0_122; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4746 = 3'h3 == state ? _GEN_3975 : valid_0_123; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4747 = 3'h3 == state ? _GEN_3976 : valid_0_124; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4748 = 3'h3 == state ? _GEN_3977 : valid_0_125; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4749 = 3'h3 == state ? _GEN_3978 : valid_0_126; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4750 = 3'h3 == state ? _GEN_3979 : valid_0_127; // @[i_cache.scala 55:18 21:26]
  wire  _GEN_4751 = 3'h3 == state ? _GEN_3980 : quene; // @[i_cache.scala 55:18 28:24]
  wire [63:0] _GEN_4752 = 3'h3 == state ? _GEN_3981 : ram_1_0; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4753 = 3'h3 == state ? _GEN_3982 : ram_1_1; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4754 = 3'h3 == state ? _GEN_3983 : ram_1_2; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4755 = 3'h3 == state ? _GEN_3984 : ram_1_3; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4756 = 3'h3 == state ? _GEN_3985 : ram_1_4; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4757 = 3'h3 == state ? _GEN_3986 : ram_1_5; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4758 = 3'h3 == state ? _GEN_3987 : ram_1_6; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4759 = 3'h3 == state ? _GEN_3988 : ram_1_7; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4760 = 3'h3 == state ? _GEN_3989 : ram_1_8; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4761 = 3'h3 == state ? _GEN_3990 : ram_1_9; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4762 = 3'h3 == state ? _GEN_3991 : ram_1_10; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4763 = 3'h3 == state ? _GEN_3992 : ram_1_11; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4764 = 3'h3 == state ? _GEN_3993 : ram_1_12; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4765 = 3'h3 == state ? _GEN_3994 : ram_1_13; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4766 = 3'h3 == state ? _GEN_3995 : ram_1_14; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4767 = 3'h3 == state ? _GEN_3996 : ram_1_15; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4768 = 3'h3 == state ? _GEN_3997 : ram_1_16; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4769 = 3'h3 == state ? _GEN_3998 : ram_1_17; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4770 = 3'h3 == state ? _GEN_3999 : ram_1_18; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4771 = 3'h3 == state ? _GEN_4000 : ram_1_19; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4772 = 3'h3 == state ? _GEN_4001 : ram_1_20; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4773 = 3'h3 == state ? _GEN_4002 : ram_1_21; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4774 = 3'h3 == state ? _GEN_4003 : ram_1_22; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4775 = 3'h3 == state ? _GEN_4004 : ram_1_23; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4776 = 3'h3 == state ? _GEN_4005 : ram_1_24; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4777 = 3'h3 == state ? _GEN_4006 : ram_1_25; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4778 = 3'h3 == state ? _GEN_4007 : ram_1_26; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4779 = 3'h3 == state ? _GEN_4008 : ram_1_27; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4780 = 3'h3 == state ? _GEN_4009 : ram_1_28; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4781 = 3'h3 == state ? _GEN_4010 : ram_1_29; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4782 = 3'h3 == state ? _GEN_4011 : ram_1_30; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4783 = 3'h3 == state ? _GEN_4012 : ram_1_31; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4784 = 3'h3 == state ? _GEN_4013 : ram_1_32; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4785 = 3'h3 == state ? _GEN_4014 : ram_1_33; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4786 = 3'h3 == state ? _GEN_4015 : ram_1_34; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4787 = 3'h3 == state ? _GEN_4016 : ram_1_35; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4788 = 3'h3 == state ? _GEN_4017 : ram_1_36; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4789 = 3'h3 == state ? _GEN_4018 : ram_1_37; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4790 = 3'h3 == state ? _GEN_4019 : ram_1_38; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4791 = 3'h3 == state ? _GEN_4020 : ram_1_39; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4792 = 3'h3 == state ? _GEN_4021 : ram_1_40; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4793 = 3'h3 == state ? _GEN_4022 : ram_1_41; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4794 = 3'h3 == state ? _GEN_4023 : ram_1_42; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4795 = 3'h3 == state ? _GEN_4024 : ram_1_43; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4796 = 3'h3 == state ? _GEN_4025 : ram_1_44; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4797 = 3'h3 == state ? _GEN_4026 : ram_1_45; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4798 = 3'h3 == state ? _GEN_4027 : ram_1_46; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4799 = 3'h3 == state ? _GEN_4028 : ram_1_47; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4800 = 3'h3 == state ? _GEN_4029 : ram_1_48; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4801 = 3'h3 == state ? _GEN_4030 : ram_1_49; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4802 = 3'h3 == state ? _GEN_4031 : ram_1_50; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4803 = 3'h3 == state ? _GEN_4032 : ram_1_51; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4804 = 3'h3 == state ? _GEN_4033 : ram_1_52; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4805 = 3'h3 == state ? _GEN_4034 : ram_1_53; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4806 = 3'h3 == state ? _GEN_4035 : ram_1_54; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4807 = 3'h3 == state ? _GEN_4036 : ram_1_55; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4808 = 3'h3 == state ? _GEN_4037 : ram_1_56; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4809 = 3'h3 == state ? _GEN_4038 : ram_1_57; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4810 = 3'h3 == state ? _GEN_4039 : ram_1_58; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4811 = 3'h3 == state ? _GEN_4040 : ram_1_59; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4812 = 3'h3 == state ? _GEN_4041 : ram_1_60; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4813 = 3'h3 == state ? _GEN_4042 : ram_1_61; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4814 = 3'h3 == state ? _GEN_4043 : ram_1_62; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4815 = 3'h3 == state ? _GEN_4044 : ram_1_63; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4816 = 3'h3 == state ? _GEN_4045 : ram_1_64; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4817 = 3'h3 == state ? _GEN_4046 : ram_1_65; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4818 = 3'h3 == state ? _GEN_4047 : ram_1_66; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4819 = 3'h3 == state ? _GEN_4048 : ram_1_67; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4820 = 3'h3 == state ? _GEN_4049 : ram_1_68; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4821 = 3'h3 == state ? _GEN_4050 : ram_1_69; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4822 = 3'h3 == state ? _GEN_4051 : ram_1_70; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4823 = 3'h3 == state ? _GEN_4052 : ram_1_71; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4824 = 3'h3 == state ? _GEN_4053 : ram_1_72; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4825 = 3'h3 == state ? _GEN_4054 : ram_1_73; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4826 = 3'h3 == state ? _GEN_4055 : ram_1_74; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4827 = 3'h3 == state ? _GEN_4056 : ram_1_75; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4828 = 3'h3 == state ? _GEN_4057 : ram_1_76; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4829 = 3'h3 == state ? _GEN_4058 : ram_1_77; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4830 = 3'h3 == state ? _GEN_4059 : ram_1_78; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4831 = 3'h3 == state ? _GEN_4060 : ram_1_79; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4832 = 3'h3 == state ? _GEN_4061 : ram_1_80; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4833 = 3'h3 == state ? _GEN_4062 : ram_1_81; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4834 = 3'h3 == state ? _GEN_4063 : ram_1_82; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4835 = 3'h3 == state ? _GEN_4064 : ram_1_83; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4836 = 3'h3 == state ? _GEN_4065 : ram_1_84; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4837 = 3'h3 == state ? _GEN_4066 : ram_1_85; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4838 = 3'h3 == state ? _GEN_4067 : ram_1_86; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4839 = 3'h3 == state ? _GEN_4068 : ram_1_87; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4840 = 3'h3 == state ? _GEN_4069 : ram_1_88; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4841 = 3'h3 == state ? _GEN_4070 : ram_1_89; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4842 = 3'h3 == state ? _GEN_4071 : ram_1_90; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4843 = 3'h3 == state ? _GEN_4072 : ram_1_91; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4844 = 3'h3 == state ? _GEN_4073 : ram_1_92; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4845 = 3'h3 == state ? _GEN_4074 : ram_1_93; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4846 = 3'h3 == state ? _GEN_4075 : ram_1_94; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4847 = 3'h3 == state ? _GEN_4076 : ram_1_95; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4848 = 3'h3 == state ? _GEN_4077 : ram_1_96; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4849 = 3'h3 == state ? _GEN_4078 : ram_1_97; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4850 = 3'h3 == state ? _GEN_4079 : ram_1_98; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4851 = 3'h3 == state ? _GEN_4080 : ram_1_99; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4852 = 3'h3 == state ? _GEN_4081 : ram_1_100; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4853 = 3'h3 == state ? _GEN_4082 : ram_1_101; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4854 = 3'h3 == state ? _GEN_4083 : ram_1_102; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4855 = 3'h3 == state ? _GEN_4084 : ram_1_103; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4856 = 3'h3 == state ? _GEN_4085 : ram_1_104; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4857 = 3'h3 == state ? _GEN_4086 : ram_1_105; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4858 = 3'h3 == state ? _GEN_4087 : ram_1_106; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4859 = 3'h3 == state ? _GEN_4088 : ram_1_107; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4860 = 3'h3 == state ? _GEN_4089 : ram_1_108; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4861 = 3'h3 == state ? _GEN_4090 : ram_1_109; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4862 = 3'h3 == state ? _GEN_4091 : ram_1_110; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4863 = 3'h3 == state ? _GEN_4092 : ram_1_111; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4864 = 3'h3 == state ? _GEN_4093 : ram_1_112; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4865 = 3'h3 == state ? _GEN_4094 : ram_1_113; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4866 = 3'h3 == state ? _GEN_4095 : ram_1_114; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4867 = 3'h3 == state ? _GEN_4096 : ram_1_115; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4868 = 3'h3 == state ? _GEN_4097 : ram_1_116; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4869 = 3'h3 == state ? _GEN_4098 : ram_1_117; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4870 = 3'h3 == state ? _GEN_4099 : ram_1_118; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4871 = 3'h3 == state ? _GEN_4100 : ram_1_119; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4872 = 3'h3 == state ? _GEN_4101 : ram_1_120; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4873 = 3'h3 == state ? _GEN_4102 : ram_1_121; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4874 = 3'h3 == state ? _GEN_4103 : ram_1_122; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4875 = 3'h3 == state ? _GEN_4104 : ram_1_123; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4876 = 3'h3 == state ? _GEN_4105 : ram_1_124; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4877 = 3'h3 == state ? _GEN_4106 : ram_1_125; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4878 = 3'h3 == state ? _GEN_4107 : ram_1_126; // @[i_cache.scala 55:18 18:24]
  wire [63:0] _GEN_4879 = 3'h3 == state ? _GEN_4108 : ram_1_127; // @[i_cache.scala 55:18 18:24]
  wire [31:0] _GEN_4880 = 3'h3 == state ? _GEN_4109 : tag_1_0; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4881 = 3'h3 == state ? _GEN_4110 : tag_1_1; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4882 = 3'h3 == state ? _GEN_4111 : tag_1_2; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4883 = 3'h3 == state ? _GEN_4112 : tag_1_3; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4884 = 3'h3 == state ? _GEN_4113 : tag_1_4; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4885 = 3'h3 == state ? _GEN_4114 : tag_1_5; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4886 = 3'h3 == state ? _GEN_4115 : tag_1_6; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4887 = 3'h3 == state ? _GEN_4116 : tag_1_7; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4888 = 3'h3 == state ? _GEN_4117 : tag_1_8; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4889 = 3'h3 == state ? _GEN_4118 : tag_1_9; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4890 = 3'h3 == state ? _GEN_4119 : tag_1_10; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4891 = 3'h3 == state ? _GEN_4120 : tag_1_11; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4892 = 3'h3 == state ? _GEN_4121 : tag_1_12; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4893 = 3'h3 == state ? _GEN_4122 : tag_1_13; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4894 = 3'h3 == state ? _GEN_4123 : tag_1_14; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4895 = 3'h3 == state ? _GEN_4124 : tag_1_15; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4896 = 3'h3 == state ? _GEN_4125 : tag_1_16; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4897 = 3'h3 == state ? _GEN_4126 : tag_1_17; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4898 = 3'h3 == state ? _GEN_4127 : tag_1_18; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4899 = 3'h3 == state ? _GEN_4128 : tag_1_19; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4900 = 3'h3 == state ? _GEN_4129 : tag_1_20; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4901 = 3'h3 == state ? _GEN_4130 : tag_1_21; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4902 = 3'h3 == state ? _GEN_4131 : tag_1_22; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4903 = 3'h3 == state ? _GEN_4132 : tag_1_23; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4904 = 3'h3 == state ? _GEN_4133 : tag_1_24; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4905 = 3'h3 == state ? _GEN_4134 : tag_1_25; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4906 = 3'h3 == state ? _GEN_4135 : tag_1_26; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4907 = 3'h3 == state ? _GEN_4136 : tag_1_27; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4908 = 3'h3 == state ? _GEN_4137 : tag_1_28; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4909 = 3'h3 == state ? _GEN_4138 : tag_1_29; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4910 = 3'h3 == state ? _GEN_4139 : tag_1_30; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4911 = 3'h3 == state ? _GEN_4140 : tag_1_31; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4912 = 3'h3 == state ? _GEN_4141 : tag_1_32; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4913 = 3'h3 == state ? _GEN_4142 : tag_1_33; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4914 = 3'h3 == state ? _GEN_4143 : tag_1_34; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4915 = 3'h3 == state ? _GEN_4144 : tag_1_35; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4916 = 3'h3 == state ? _GEN_4145 : tag_1_36; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4917 = 3'h3 == state ? _GEN_4146 : tag_1_37; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4918 = 3'h3 == state ? _GEN_4147 : tag_1_38; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4919 = 3'h3 == state ? _GEN_4148 : tag_1_39; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4920 = 3'h3 == state ? _GEN_4149 : tag_1_40; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4921 = 3'h3 == state ? _GEN_4150 : tag_1_41; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4922 = 3'h3 == state ? _GEN_4151 : tag_1_42; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4923 = 3'h3 == state ? _GEN_4152 : tag_1_43; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4924 = 3'h3 == state ? _GEN_4153 : tag_1_44; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4925 = 3'h3 == state ? _GEN_4154 : tag_1_45; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4926 = 3'h3 == state ? _GEN_4155 : tag_1_46; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4927 = 3'h3 == state ? _GEN_4156 : tag_1_47; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4928 = 3'h3 == state ? _GEN_4157 : tag_1_48; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4929 = 3'h3 == state ? _GEN_4158 : tag_1_49; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4930 = 3'h3 == state ? _GEN_4159 : tag_1_50; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4931 = 3'h3 == state ? _GEN_4160 : tag_1_51; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4932 = 3'h3 == state ? _GEN_4161 : tag_1_52; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4933 = 3'h3 == state ? _GEN_4162 : tag_1_53; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4934 = 3'h3 == state ? _GEN_4163 : tag_1_54; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4935 = 3'h3 == state ? _GEN_4164 : tag_1_55; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4936 = 3'h3 == state ? _GEN_4165 : tag_1_56; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4937 = 3'h3 == state ? _GEN_4166 : tag_1_57; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4938 = 3'h3 == state ? _GEN_4167 : tag_1_58; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4939 = 3'h3 == state ? _GEN_4168 : tag_1_59; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4940 = 3'h3 == state ? _GEN_4169 : tag_1_60; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4941 = 3'h3 == state ? _GEN_4170 : tag_1_61; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4942 = 3'h3 == state ? _GEN_4171 : tag_1_62; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4943 = 3'h3 == state ? _GEN_4172 : tag_1_63; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4944 = 3'h3 == state ? _GEN_4173 : tag_1_64; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4945 = 3'h3 == state ? _GEN_4174 : tag_1_65; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4946 = 3'h3 == state ? _GEN_4175 : tag_1_66; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4947 = 3'h3 == state ? _GEN_4176 : tag_1_67; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4948 = 3'h3 == state ? _GEN_4177 : tag_1_68; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4949 = 3'h3 == state ? _GEN_4178 : tag_1_69; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4950 = 3'h3 == state ? _GEN_4179 : tag_1_70; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4951 = 3'h3 == state ? _GEN_4180 : tag_1_71; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4952 = 3'h3 == state ? _GEN_4181 : tag_1_72; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4953 = 3'h3 == state ? _GEN_4182 : tag_1_73; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4954 = 3'h3 == state ? _GEN_4183 : tag_1_74; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4955 = 3'h3 == state ? _GEN_4184 : tag_1_75; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4956 = 3'h3 == state ? _GEN_4185 : tag_1_76; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4957 = 3'h3 == state ? _GEN_4186 : tag_1_77; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4958 = 3'h3 == state ? _GEN_4187 : tag_1_78; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4959 = 3'h3 == state ? _GEN_4188 : tag_1_79; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4960 = 3'h3 == state ? _GEN_4189 : tag_1_80; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4961 = 3'h3 == state ? _GEN_4190 : tag_1_81; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4962 = 3'h3 == state ? _GEN_4191 : tag_1_82; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4963 = 3'h3 == state ? _GEN_4192 : tag_1_83; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4964 = 3'h3 == state ? _GEN_4193 : tag_1_84; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4965 = 3'h3 == state ? _GEN_4194 : tag_1_85; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4966 = 3'h3 == state ? _GEN_4195 : tag_1_86; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4967 = 3'h3 == state ? _GEN_4196 : tag_1_87; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4968 = 3'h3 == state ? _GEN_4197 : tag_1_88; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4969 = 3'h3 == state ? _GEN_4198 : tag_1_89; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4970 = 3'h3 == state ? _GEN_4199 : tag_1_90; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4971 = 3'h3 == state ? _GEN_4200 : tag_1_91; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4972 = 3'h3 == state ? _GEN_4201 : tag_1_92; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4973 = 3'h3 == state ? _GEN_4202 : tag_1_93; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4974 = 3'h3 == state ? _GEN_4203 : tag_1_94; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4975 = 3'h3 == state ? _GEN_4204 : tag_1_95; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4976 = 3'h3 == state ? _GEN_4205 : tag_1_96; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4977 = 3'h3 == state ? _GEN_4206 : tag_1_97; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4978 = 3'h3 == state ? _GEN_4207 : tag_1_98; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4979 = 3'h3 == state ? _GEN_4208 : tag_1_99; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4980 = 3'h3 == state ? _GEN_4209 : tag_1_100; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4981 = 3'h3 == state ? _GEN_4210 : tag_1_101; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4982 = 3'h3 == state ? _GEN_4211 : tag_1_102; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4983 = 3'h3 == state ? _GEN_4212 : tag_1_103; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4984 = 3'h3 == state ? _GEN_4213 : tag_1_104; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4985 = 3'h3 == state ? _GEN_4214 : tag_1_105; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4986 = 3'h3 == state ? _GEN_4215 : tag_1_106; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4987 = 3'h3 == state ? _GEN_4216 : tag_1_107; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4988 = 3'h3 == state ? _GEN_4217 : tag_1_108; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4989 = 3'h3 == state ? _GEN_4218 : tag_1_109; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4990 = 3'h3 == state ? _GEN_4219 : tag_1_110; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4991 = 3'h3 == state ? _GEN_4220 : tag_1_111; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4992 = 3'h3 == state ? _GEN_4221 : tag_1_112; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4993 = 3'h3 == state ? _GEN_4222 : tag_1_113; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4994 = 3'h3 == state ? _GEN_4223 : tag_1_114; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4995 = 3'h3 == state ? _GEN_4224 : tag_1_115; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4996 = 3'h3 == state ? _GEN_4225 : tag_1_116; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4997 = 3'h3 == state ? _GEN_4226 : tag_1_117; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4998 = 3'h3 == state ? _GEN_4227 : tag_1_118; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_4999 = 3'h3 == state ? _GEN_4228 : tag_1_119; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5000 = 3'h3 == state ? _GEN_4229 : tag_1_120; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5001 = 3'h3 == state ? _GEN_4230 : tag_1_121; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5002 = 3'h3 == state ? _GEN_4231 : tag_1_122; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5003 = 3'h3 == state ? _GEN_4232 : tag_1_123; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5004 = 3'h3 == state ? _GEN_4233 : tag_1_124; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5005 = 3'h3 == state ? _GEN_4234 : tag_1_125; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5006 = 3'h3 == state ? _GEN_4235 : tag_1_126; // @[i_cache.scala 55:18 20:24]
  wire [31:0] _GEN_5007 = 3'h3 == state ? _GEN_4236 : tag_1_127; // @[i_cache.scala 55:18 20:24]
  wire  _GEN_5008 = 3'h3 == state ? _GEN_4237 : valid_1_0; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5009 = 3'h3 == state ? _GEN_4238 : valid_1_1; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5010 = 3'h3 == state ? _GEN_4239 : valid_1_2; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5011 = 3'h3 == state ? _GEN_4240 : valid_1_3; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5012 = 3'h3 == state ? _GEN_4241 : valid_1_4; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5013 = 3'h3 == state ? _GEN_4242 : valid_1_5; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5014 = 3'h3 == state ? _GEN_4243 : valid_1_6; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5015 = 3'h3 == state ? _GEN_4244 : valid_1_7; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5016 = 3'h3 == state ? _GEN_4245 : valid_1_8; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5017 = 3'h3 == state ? _GEN_4246 : valid_1_9; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5018 = 3'h3 == state ? _GEN_4247 : valid_1_10; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5019 = 3'h3 == state ? _GEN_4248 : valid_1_11; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5020 = 3'h3 == state ? _GEN_4249 : valid_1_12; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5021 = 3'h3 == state ? _GEN_4250 : valid_1_13; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5022 = 3'h3 == state ? _GEN_4251 : valid_1_14; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5023 = 3'h3 == state ? _GEN_4252 : valid_1_15; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5024 = 3'h3 == state ? _GEN_4253 : valid_1_16; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5025 = 3'h3 == state ? _GEN_4254 : valid_1_17; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5026 = 3'h3 == state ? _GEN_4255 : valid_1_18; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5027 = 3'h3 == state ? _GEN_4256 : valid_1_19; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5028 = 3'h3 == state ? _GEN_4257 : valid_1_20; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5029 = 3'h3 == state ? _GEN_4258 : valid_1_21; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5030 = 3'h3 == state ? _GEN_4259 : valid_1_22; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5031 = 3'h3 == state ? _GEN_4260 : valid_1_23; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5032 = 3'h3 == state ? _GEN_4261 : valid_1_24; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5033 = 3'h3 == state ? _GEN_4262 : valid_1_25; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5034 = 3'h3 == state ? _GEN_4263 : valid_1_26; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5035 = 3'h3 == state ? _GEN_4264 : valid_1_27; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5036 = 3'h3 == state ? _GEN_4265 : valid_1_28; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5037 = 3'h3 == state ? _GEN_4266 : valid_1_29; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5038 = 3'h3 == state ? _GEN_4267 : valid_1_30; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5039 = 3'h3 == state ? _GEN_4268 : valid_1_31; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5040 = 3'h3 == state ? _GEN_4269 : valid_1_32; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5041 = 3'h3 == state ? _GEN_4270 : valid_1_33; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5042 = 3'h3 == state ? _GEN_4271 : valid_1_34; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5043 = 3'h3 == state ? _GEN_4272 : valid_1_35; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5044 = 3'h3 == state ? _GEN_4273 : valid_1_36; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5045 = 3'h3 == state ? _GEN_4274 : valid_1_37; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5046 = 3'h3 == state ? _GEN_4275 : valid_1_38; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5047 = 3'h3 == state ? _GEN_4276 : valid_1_39; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5048 = 3'h3 == state ? _GEN_4277 : valid_1_40; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5049 = 3'h3 == state ? _GEN_4278 : valid_1_41; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5050 = 3'h3 == state ? _GEN_4279 : valid_1_42; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5051 = 3'h3 == state ? _GEN_4280 : valid_1_43; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5052 = 3'h3 == state ? _GEN_4281 : valid_1_44; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5053 = 3'h3 == state ? _GEN_4282 : valid_1_45; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5054 = 3'h3 == state ? _GEN_4283 : valid_1_46; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5055 = 3'h3 == state ? _GEN_4284 : valid_1_47; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5056 = 3'h3 == state ? _GEN_4285 : valid_1_48; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5057 = 3'h3 == state ? _GEN_4286 : valid_1_49; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5058 = 3'h3 == state ? _GEN_4287 : valid_1_50; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5059 = 3'h3 == state ? _GEN_4288 : valid_1_51; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5060 = 3'h3 == state ? _GEN_4289 : valid_1_52; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5061 = 3'h3 == state ? _GEN_4290 : valid_1_53; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5062 = 3'h3 == state ? _GEN_4291 : valid_1_54; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5063 = 3'h3 == state ? _GEN_4292 : valid_1_55; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5064 = 3'h3 == state ? _GEN_4293 : valid_1_56; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5065 = 3'h3 == state ? _GEN_4294 : valid_1_57; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5066 = 3'h3 == state ? _GEN_4295 : valid_1_58; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5067 = 3'h3 == state ? _GEN_4296 : valid_1_59; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5068 = 3'h3 == state ? _GEN_4297 : valid_1_60; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5069 = 3'h3 == state ? _GEN_4298 : valid_1_61; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5070 = 3'h3 == state ? _GEN_4299 : valid_1_62; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5071 = 3'h3 == state ? _GEN_4300 : valid_1_63; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5072 = 3'h3 == state ? _GEN_4301 : valid_1_64; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5073 = 3'h3 == state ? _GEN_4302 : valid_1_65; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5074 = 3'h3 == state ? _GEN_4303 : valid_1_66; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5075 = 3'h3 == state ? _GEN_4304 : valid_1_67; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5076 = 3'h3 == state ? _GEN_4305 : valid_1_68; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5077 = 3'h3 == state ? _GEN_4306 : valid_1_69; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5078 = 3'h3 == state ? _GEN_4307 : valid_1_70; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5079 = 3'h3 == state ? _GEN_4308 : valid_1_71; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5080 = 3'h3 == state ? _GEN_4309 : valid_1_72; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5081 = 3'h3 == state ? _GEN_4310 : valid_1_73; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5082 = 3'h3 == state ? _GEN_4311 : valid_1_74; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5083 = 3'h3 == state ? _GEN_4312 : valid_1_75; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5084 = 3'h3 == state ? _GEN_4313 : valid_1_76; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5085 = 3'h3 == state ? _GEN_4314 : valid_1_77; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5086 = 3'h3 == state ? _GEN_4315 : valid_1_78; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5087 = 3'h3 == state ? _GEN_4316 : valid_1_79; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5088 = 3'h3 == state ? _GEN_4317 : valid_1_80; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5089 = 3'h3 == state ? _GEN_4318 : valid_1_81; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5090 = 3'h3 == state ? _GEN_4319 : valid_1_82; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5091 = 3'h3 == state ? _GEN_4320 : valid_1_83; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5092 = 3'h3 == state ? _GEN_4321 : valid_1_84; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5093 = 3'h3 == state ? _GEN_4322 : valid_1_85; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5094 = 3'h3 == state ? _GEN_4323 : valid_1_86; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5095 = 3'h3 == state ? _GEN_4324 : valid_1_87; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5096 = 3'h3 == state ? _GEN_4325 : valid_1_88; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5097 = 3'h3 == state ? _GEN_4326 : valid_1_89; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5098 = 3'h3 == state ? _GEN_4327 : valid_1_90; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5099 = 3'h3 == state ? _GEN_4328 : valid_1_91; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5100 = 3'h3 == state ? _GEN_4329 : valid_1_92; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5101 = 3'h3 == state ? _GEN_4330 : valid_1_93; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5102 = 3'h3 == state ? _GEN_4331 : valid_1_94; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5103 = 3'h3 == state ? _GEN_4332 : valid_1_95; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5104 = 3'h3 == state ? _GEN_4333 : valid_1_96; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5105 = 3'h3 == state ? _GEN_4334 : valid_1_97; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5106 = 3'h3 == state ? _GEN_4335 : valid_1_98; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5107 = 3'h3 == state ? _GEN_4336 : valid_1_99; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5108 = 3'h3 == state ? _GEN_4337 : valid_1_100; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5109 = 3'h3 == state ? _GEN_4338 : valid_1_101; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5110 = 3'h3 == state ? _GEN_4339 : valid_1_102; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5111 = 3'h3 == state ? _GEN_4340 : valid_1_103; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5112 = 3'h3 == state ? _GEN_4341 : valid_1_104; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5113 = 3'h3 == state ? _GEN_4342 : valid_1_105; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5114 = 3'h3 == state ? _GEN_4343 : valid_1_106; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5115 = 3'h3 == state ? _GEN_4344 : valid_1_107; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5116 = 3'h3 == state ? _GEN_4345 : valid_1_108; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5117 = 3'h3 == state ? _GEN_4346 : valid_1_109; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5118 = 3'h3 == state ? _GEN_4347 : valid_1_110; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5119 = 3'h3 == state ? _GEN_4348 : valid_1_111; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5120 = 3'h3 == state ? _GEN_4349 : valid_1_112; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5121 = 3'h3 == state ? _GEN_4350 : valid_1_113; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5122 = 3'h3 == state ? _GEN_4351 : valid_1_114; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5123 = 3'h3 == state ? _GEN_4352 : valid_1_115; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5124 = 3'h3 == state ? _GEN_4353 : valid_1_116; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5125 = 3'h3 == state ? _GEN_4354 : valid_1_117; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5126 = 3'h3 == state ? _GEN_4355 : valid_1_118; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5127 = 3'h3 == state ? _GEN_4356 : valid_1_119; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5128 = 3'h3 == state ? _GEN_4357 : valid_1_120; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5129 = 3'h3 == state ? _GEN_4358 : valid_1_121; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5130 = 3'h3 == state ? _GEN_4359 : valid_1_122; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5131 = 3'h3 == state ? _GEN_4360 : valid_1_123; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5132 = 3'h3 == state ? _GEN_4361 : valid_1_124; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5133 = 3'h3 == state ? _GEN_4362 : valid_1_125; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5134 = 3'h3 == state ? _GEN_4363 : valid_1_126; // @[i_cache.scala 55:18 22:26]
  wire  _GEN_5135 = 3'h3 == state ? _GEN_4364 : valid_1_127; // @[i_cache.scala 55:18 22:26]
  wire [63:0] _GEN_7450 = 7'h1 == index ? ram_0_1 : ram_0_0; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7451 = 7'h2 == index ? ram_0_2 : _GEN_7450; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7452 = 7'h3 == index ? ram_0_3 : _GEN_7451; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7453 = 7'h4 == index ? ram_0_4 : _GEN_7452; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7454 = 7'h5 == index ? ram_0_5 : _GEN_7453; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7455 = 7'h6 == index ? ram_0_6 : _GEN_7454; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7456 = 7'h7 == index ? ram_0_7 : _GEN_7455; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7457 = 7'h8 == index ? ram_0_8 : _GEN_7456; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7458 = 7'h9 == index ? ram_0_9 : _GEN_7457; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7459 = 7'ha == index ? ram_0_10 : _GEN_7458; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7460 = 7'hb == index ? ram_0_11 : _GEN_7459; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7461 = 7'hc == index ? ram_0_12 : _GEN_7460; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7462 = 7'hd == index ? ram_0_13 : _GEN_7461; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7463 = 7'he == index ? ram_0_14 : _GEN_7462; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7464 = 7'hf == index ? ram_0_15 : _GEN_7463; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7465 = 7'h10 == index ? ram_0_16 : _GEN_7464; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7466 = 7'h11 == index ? ram_0_17 : _GEN_7465; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7467 = 7'h12 == index ? ram_0_18 : _GEN_7466; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7468 = 7'h13 == index ? ram_0_19 : _GEN_7467; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7469 = 7'h14 == index ? ram_0_20 : _GEN_7468; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7470 = 7'h15 == index ? ram_0_21 : _GEN_7469; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7471 = 7'h16 == index ? ram_0_22 : _GEN_7470; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7472 = 7'h17 == index ? ram_0_23 : _GEN_7471; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7473 = 7'h18 == index ? ram_0_24 : _GEN_7472; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7474 = 7'h19 == index ? ram_0_25 : _GEN_7473; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7475 = 7'h1a == index ? ram_0_26 : _GEN_7474; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7476 = 7'h1b == index ? ram_0_27 : _GEN_7475; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7477 = 7'h1c == index ? ram_0_28 : _GEN_7476; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7478 = 7'h1d == index ? ram_0_29 : _GEN_7477; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7479 = 7'h1e == index ? ram_0_30 : _GEN_7478; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7480 = 7'h1f == index ? ram_0_31 : _GEN_7479; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7481 = 7'h20 == index ? ram_0_32 : _GEN_7480; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7482 = 7'h21 == index ? ram_0_33 : _GEN_7481; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7483 = 7'h22 == index ? ram_0_34 : _GEN_7482; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7484 = 7'h23 == index ? ram_0_35 : _GEN_7483; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7485 = 7'h24 == index ? ram_0_36 : _GEN_7484; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7486 = 7'h25 == index ? ram_0_37 : _GEN_7485; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7487 = 7'h26 == index ? ram_0_38 : _GEN_7486; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7488 = 7'h27 == index ? ram_0_39 : _GEN_7487; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7489 = 7'h28 == index ? ram_0_40 : _GEN_7488; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7490 = 7'h29 == index ? ram_0_41 : _GEN_7489; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7491 = 7'h2a == index ? ram_0_42 : _GEN_7490; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7492 = 7'h2b == index ? ram_0_43 : _GEN_7491; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7493 = 7'h2c == index ? ram_0_44 : _GEN_7492; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7494 = 7'h2d == index ? ram_0_45 : _GEN_7493; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7495 = 7'h2e == index ? ram_0_46 : _GEN_7494; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7496 = 7'h2f == index ? ram_0_47 : _GEN_7495; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7497 = 7'h30 == index ? ram_0_48 : _GEN_7496; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7498 = 7'h31 == index ? ram_0_49 : _GEN_7497; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7499 = 7'h32 == index ? ram_0_50 : _GEN_7498; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7500 = 7'h33 == index ? ram_0_51 : _GEN_7499; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7501 = 7'h34 == index ? ram_0_52 : _GEN_7500; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7502 = 7'h35 == index ? ram_0_53 : _GEN_7501; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7503 = 7'h36 == index ? ram_0_54 : _GEN_7502; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7504 = 7'h37 == index ? ram_0_55 : _GEN_7503; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7505 = 7'h38 == index ? ram_0_56 : _GEN_7504; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7506 = 7'h39 == index ? ram_0_57 : _GEN_7505; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7507 = 7'h3a == index ? ram_0_58 : _GEN_7506; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7508 = 7'h3b == index ? ram_0_59 : _GEN_7507; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7509 = 7'h3c == index ? ram_0_60 : _GEN_7508; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7510 = 7'h3d == index ? ram_0_61 : _GEN_7509; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7511 = 7'h3e == index ? ram_0_62 : _GEN_7510; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7512 = 7'h3f == index ? ram_0_63 : _GEN_7511; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7513 = 7'h40 == index ? ram_0_64 : _GEN_7512; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7514 = 7'h41 == index ? ram_0_65 : _GEN_7513; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7515 = 7'h42 == index ? ram_0_66 : _GEN_7514; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7516 = 7'h43 == index ? ram_0_67 : _GEN_7515; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7517 = 7'h44 == index ? ram_0_68 : _GEN_7516; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7518 = 7'h45 == index ? ram_0_69 : _GEN_7517; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7519 = 7'h46 == index ? ram_0_70 : _GEN_7518; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7520 = 7'h47 == index ? ram_0_71 : _GEN_7519; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7521 = 7'h48 == index ? ram_0_72 : _GEN_7520; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7522 = 7'h49 == index ? ram_0_73 : _GEN_7521; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7523 = 7'h4a == index ? ram_0_74 : _GEN_7522; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7524 = 7'h4b == index ? ram_0_75 : _GEN_7523; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7525 = 7'h4c == index ? ram_0_76 : _GEN_7524; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7526 = 7'h4d == index ? ram_0_77 : _GEN_7525; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7527 = 7'h4e == index ? ram_0_78 : _GEN_7526; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7528 = 7'h4f == index ? ram_0_79 : _GEN_7527; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7529 = 7'h50 == index ? ram_0_80 : _GEN_7528; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7530 = 7'h51 == index ? ram_0_81 : _GEN_7529; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7531 = 7'h52 == index ? ram_0_82 : _GEN_7530; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7532 = 7'h53 == index ? ram_0_83 : _GEN_7531; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7533 = 7'h54 == index ? ram_0_84 : _GEN_7532; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7534 = 7'h55 == index ? ram_0_85 : _GEN_7533; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7535 = 7'h56 == index ? ram_0_86 : _GEN_7534; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7536 = 7'h57 == index ? ram_0_87 : _GEN_7535; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7537 = 7'h58 == index ? ram_0_88 : _GEN_7536; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7538 = 7'h59 == index ? ram_0_89 : _GEN_7537; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7539 = 7'h5a == index ? ram_0_90 : _GEN_7538; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7540 = 7'h5b == index ? ram_0_91 : _GEN_7539; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7541 = 7'h5c == index ? ram_0_92 : _GEN_7540; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7542 = 7'h5d == index ? ram_0_93 : _GEN_7541; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7543 = 7'h5e == index ? ram_0_94 : _GEN_7542; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7544 = 7'h5f == index ? ram_0_95 : _GEN_7543; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7545 = 7'h60 == index ? ram_0_96 : _GEN_7544; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7546 = 7'h61 == index ? ram_0_97 : _GEN_7545; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7547 = 7'h62 == index ? ram_0_98 : _GEN_7546; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7548 = 7'h63 == index ? ram_0_99 : _GEN_7547; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7549 = 7'h64 == index ? ram_0_100 : _GEN_7548; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7550 = 7'h65 == index ? ram_0_101 : _GEN_7549; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7551 = 7'h66 == index ? ram_0_102 : _GEN_7550; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7552 = 7'h67 == index ? ram_0_103 : _GEN_7551; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7553 = 7'h68 == index ? ram_0_104 : _GEN_7552; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7554 = 7'h69 == index ? ram_0_105 : _GEN_7553; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7555 = 7'h6a == index ? ram_0_106 : _GEN_7554; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7556 = 7'h6b == index ? ram_0_107 : _GEN_7555; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7557 = 7'h6c == index ? ram_0_108 : _GEN_7556; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7558 = 7'h6d == index ? ram_0_109 : _GEN_7557; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7559 = 7'h6e == index ? ram_0_110 : _GEN_7558; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7560 = 7'h6f == index ? ram_0_111 : _GEN_7559; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7561 = 7'h70 == index ? ram_0_112 : _GEN_7560; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7562 = 7'h71 == index ? ram_0_113 : _GEN_7561; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7563 = 7'h72 == index ? ram_0_114 : _GEN_7562; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7564 = 7'h73 == index ? ram_0_115 : _GEN_7563; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7565 = 7'h74 == index ? ram_0_116 : _GEN_7564; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7566 = 7'h75 == index ? ram_0_117 : _GEN_7565; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7567 = 7'h76 == index ? ram_0_118 : _GEN_7566; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7568 = 7'h77 == index ? ram_0_119 : _GEN_7567; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7569 = 7'h78 == index ? ram_0_120 : _GEN_7568; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7570 = 7'h79 == index ? ram_0_121 : _GEN_7569; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7571 = 7'h7a == index ? ram_0_122 : _GEN_7570; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7572 = 7'h7b == index ? ram_0_123 : _GEN_7571; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7573 = 7'h7c == index ? ram_0_124 : _GEN_7572; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7574 = 7'h7d == index ? ram_0_125 : _GEN_7573; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7575 = 7'h7e == index ? ram_0_126 : _GEN_7574; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7576 = 7'h7f == index ? ram_0_127 : _GEN_7575; // @[i_cache.scala 141:{33,33}]
  wire [63:0] _GEN_7578 = 7'h1 == index ? ram_1_1 : ram_1_0; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7579 = 7'h2 == index ? ram_1_2 : _GEN_7578; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7580 = 7'h3 == index ? ram_1_3 : _GEN_7579; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7581 = 7'h4 == index ? ram_1_4 : _GEN_7580; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7582 = 7'h5 == index ? ram_1_5 : _GEN_7581; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7583 = 7'h6 == index ? ram_1_6 : _GEN_7582; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7584 = 7'h7 == index ? ram_1_7 : _GEN_7583; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7585 = 7'h8 == index ? ram_1_8 : _GEN_7584; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7586 = 7'h9 == index ? ram_1_9 : _GEN_7585; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7587 = 7'ha == index ? ram_1_10 : _GEN_7586; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7588 = 7'hb == index ? ram_1_11 : _GEN_7587; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7589 = 7'hc == index ? ram_1_12 : _GEN_7588; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7590 = 7'hd == index ? ram_1_13 : _GEN_7589; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7591 = 7'he == index ? ram_1_14 : _GEN_7590; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7592 = 7'hf == index ? ram_1_15 : _GEN_7591; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7593 = 7'h10 == index ? ram_1_16 : _GEN_7592; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7594 = 7'h11 == index ? ram_1_17 : _GEN_7593; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7595 = 7'h12 == index ? ram_1_18 : _GEN_7594; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7596 = 7'h13 == index ? ram_1_19 : _GEN_7595; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7597 = 7'h14 == index ? ram_1_20 : _GEN_7596; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7598 = 7'h15 == index ? ram_1_21 : _GEN_7597; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7599 = 7'h16 == index ? ram_1_22 : _GEN_7598; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7600 = 7'h17 == index ? ram_1_23 : _GEN_7599; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7601 = 7'h18 == index ? ram_1_24 : _GEN_7600; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7602 = 7'h19 == index ? ram_1_25 : _GEN_7601; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7603 = 7'h1a == index ? ram_1_26 : _GEN_7602; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7604 = 7'h1b == index ? ram_1_27 : _GEN_7603; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7605 = 7'h1c == index ? ram_1_28 : _GEN_7604; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7606 = 7'h1d == index ? ram_1_29 : _GEN_7605; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7607 = 7'h1e == index ? ram_1_30 : _GEN_7606; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7608 = 7'h1f == index ? ram_1_31 : _GEN_7607; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7609 = 7'h20 == index ? ram_1_32 : _GEN_7608; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7610 = 7'h21 == index ? ram_1_33 : _GEN_7609; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7611 = 7'h22 == index ? ram_1_34 : _GEN_7610; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7612 = 7'h23 == index ? ram_1_35 : _GEN_7611; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7613 = 7'h24 == index ? ram_1_36 : _GEN_7612; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7614 = 7'h25 == index ? ram_1_37 : _GEN_7613; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7615 = 7'h26 == index ? ram_1_38 : _GEN_7614; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7616 = 7'h27 == index ? ram_1_39 : _GEN_7615; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7617 = 7'h28 == index ? ram_1_40 : _GEN_7616; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7618 = 7'h29 == index ? ram_1_41 : _GEN_7617; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7619 = 7'h2a == index ? ram_1_42 : _GEN_7618; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7620 = 7'h2b == index ? ram_1_43 : _GEN_7619; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7621 = 7'h2c == index ? ram_1_44 : _GEN_7620; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7622 = 7'h2d == index ? ram_1_45 : _GEN_7621; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7623 = 7'h2e == index ? ram_1_46 : _GEN_7622; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7624 = 7'h2f == index ? ram_1_47 : _GEN_7623; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7625 = 7'h30 == index ? ram_1_48 : _GEN_7624; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7626 = 7'h31 == index ? ram_1_49 : _GEN_7625; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7627 = 7'h32 == index ? ram_1_50 : _GEN_7626; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7628 = 7'h33 == index ? ram_1_51 : _GEN_7627; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7629 = 7'h34 == index ? ram_1_52 : _GEN_7628; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7630 = 7'h35 == index ? ram_1_53 : _GEN_7629; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7631 = 7'h36 == index ? ram_1_54 : _GEN_7630; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7632 = 7'h37 == index ? ram_1_55 : _GEN_7631; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7633 = 7'h38 == index ? ram_1_56 : _GEN_7632; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7634 = 7'h39 == index ? ram_1_57 : _GEN_7633; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7635 = 7'h3a == index ? ram_1_58 : _GEN_7634; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7636 = 7'h3b == index ? ram_1_59 : _GEN_7635; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7637 = 7'h3c == index ? ram_1_60 : _GEN_7636; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7638 = 7'h3d == index ? ram_1_61 : _GEN_7637; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7639 = 7'h3e == index ? ram_1_62 : _GEN_7638; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7640 = 7'h3f == index ? ram_1_63 : _GEN_7639; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7641 = 7'h40 == index ? ram_1_64 : _GEN_7640; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7642 = 7'h41 == index ? ram_1_65 : _GEN_7641; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7643 = 7'h42 == index ? ram_1_66 : _GEN_7642; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7644 = 7'h43 == index ? ram_1_67 : _GEN_7643; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7645 = 7'h44 == index ? ram_1_68 : _GEN_7644; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7646 = 7'h45 == index ? ram_1_69 : _GEN_7645; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7647 = 7'h46 == index ? ram_1_70 : _GEN_7646; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7648 = 7'h47 == index ? ram_1_71 : _GEN_7647; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7649 = 7'h48 == index ? ram_1_72 : _GEN_7648; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7650 = 7'h49 == index ? ram_1_73 : _GEN_7649; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7651 = 7'h4a == index ? ram_1_74 : _GEN_7650; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7652 = 7'h4b == index ? ram_1_75 : _GEN_7651; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7653 = 7'h4c == index ? ram_1_76 : _GEN_7652; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7654 = 7'h4d == index ? ram_1_77 : _GEN_7653; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7655 = 7'h4e == index ? ram_1_78 : _GEN_7654; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7656 = 7'h4f == index ? ram_1_79 : _GEN_7655; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7657 = 7'h50 == index ? ram_1_80 : _GEN_7656; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7658 = 7'h51 == index ? ram_1_81 : _GEN_7657; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7659 = 7'h52 == index ? ram_1_82 : _GEN_7658; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7660 = 7'h53 == index ? ram_1_83 : _GEN_7659; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7661 = 7'h54 == index ? ram_1_84 : _GEN_7660; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7662 = 7'h55 == index ? ram_1_85 : _GEN_7661; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7663 = 7'h56 == index ? ram_1_86 : _GEN_7662; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7664 = 7'h57 == index ? ram_1_87 : _GEN_7663; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7665 = 7'h58 == index ? ram_1_88 : _GEN_7664; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7666 = 7'h59 == index ? ram_1_89 : _GEN_7665; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7667 = 7'h5a == index ? ram_1_90 : _GEN_7666; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7668 = 7'h5b == index ? ram_1_91 : _GEN_7667; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7669 = 7'h5c == index ? ram_1_92 : _GEN_7668; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7670 = 7'h5d == index ? ram_1_93 : _GEN_7669; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7671 = 7'h5e == index ? ram_1_94 : _GEN_7670; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7672 = 7'h5f == index ? ram_1_95 : _GEN_7671; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7673 = 7'h60 == index ? ram_1_96 : _GEN_7672; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7674 = 7'h61 == index ? ram_1_97 : _GEN_7673; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7675 = 7'h62 == index ? ram_1_98 : _GEN_7674; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7676 = 7'h63 == index ? ram_1_99 : _GEN_7675; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7677 = 7'h64 == index ? ram_1_100 : _GEN_7676; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7678 = 7'h65 == index ? ram_1_101 : _GEN_7677; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7679 = 7'h66 == index ? ram_1_102 : _GEN_7678; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7680 = 7'h67 == index ? ram_1_103 : _GEN_7679; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7681 = 7'h68 == index ? ram_1_104 : _GEN_7680; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7682 = 7'h69 == index ? ram_1_105 : _GEN_7681; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7683 = 7'h6a == index ? ram_1_106 : _GEN_7682; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7684 = 7'h6b == index ? ram_1_107 : _GEN_7683; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7685 = 7'h6c == index ? ram_1_108 : _GEN_7684; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7686 = 7'h6d == index ? ram_1_109 : _GEN_7685; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7687 = 7'h6e == index ? ram_1_110 : _GEN_7686; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7688 = 7'h6f == index ? ram_1_111 : _GEN_7687; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7689 = 7'h70 == index ? ram_1_112 : _GEN_7688; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7690 = 7'h71 == index ? ram_1_113 : _GEN_7689; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7691 = 7'h72 == index ? ram_1_114 : _GEN_7690; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7692 = 7'h73 == index ? ram_1_115 : _GEN_7691; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7693 = 7'h74 == index ? ram_1_116 : _GEN_7692; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7694 = 7'h75 == index ? ram_1_117 : _GEN_7693; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7695 = 7'h76 == index ? ram_1_118 : _GEN_7694; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7696 = 7'h77 == index ? ram_1_119 : _GEN_7695; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7697 = 7'h78 == index ? ram_1_120 : _GEN_7696; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7698 = 7'h79 == index ? ram_1_121 : _GEN_7697; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7699 = 7'h7a == index ? ram_1_122 : _GEN_7698; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7700 = 7'h7b == index ? ram_1_123 : _GEN_7699; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7701 = 7'h7c == index ? ram_1_124 : _GEN_7700; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7702 = 7'h7d == index ? ram_1_125 : _GEN_7701; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7703 = 7'h7e == index ? ram_1_126 : _GEN_7702; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7704 = 7'h7f == index ? ram_1_127 : _GEN_7703; // @[i_cache.scala 149:{33,33}]
  wire [63:0] _GEN_7705 = way1_hit ? _GEN_7704 : 64'h0; // @[i_cache.scala 148:33 149:33 156:33]
  wire [63:0] _GEN_7709 = way0_hit ? _GEN_7576 : _GEN_7705; // @[i_cache.scala 140:23 141:33]
  wire  _GEN_7711 = way0_hit | way1_hit; // @[i_cache.scala 140:23 143:34]
  wire  _T_18 = state == 3'h2; // @[i_cache.scala 163:21]
  wire  _GEN_7722 = state == 3'h1 ? 1'h0 : _T_18; // @[i_cache.scala 130:31 131:27]
  wire  _GEN_7724 = state == 3'h1 ? 1'h0 : io_from_ifu_rready; // @[i_cache.scala 130:31 133:26]
  wire [63:0] _GEN_7726 = state == 3'h1 ? _GEN_7709 : 64'h0; // @[i_cache.scala 130:31]
  wire  _GEN_7728 = state == 3'h1 & _GEN_7711; // @[i_cache.scala 130:31]
  assign io_to_ifu_rdata = state == 3'h0 ? 64'h0 : _GEN_7726; // @[i_cache.scala 114:23 115:25]
  assign io_to_ifu_rvalid = state == 3'h0 ? 1'h0 : _GEN_7728; // @[i_cache.scala 114:23 117:26]
  assign io_to_axi_araddr = io_from_ifu_araddr; // @[i_cache.scala 114:23 122:26]
  assign io_to_axi_arvalid = state == 3'h0 ? 1'h0 : _GEN_7722; // @[i_cache.scala 114:23 121:27]
  assign io_to_axi_rready = state == 3'h0 ? io_from_ifu_rready : _GEN_7724; // @[i_cache.scala 114:23 123:26]
  always @(posedge clock) begin
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_0 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_0 <= _GEN_4367;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_1 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_1 <= _GEN_4368;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_2 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_2 <= _GEN_4369;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_3 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_3 <= _GEN_4370;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_4 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_4 <= _GEN_4371;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_5 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_5 <= _GEN_4372;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_6 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_6 <= _GEN_4373;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_7 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_7 <= _GEN_4374;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_8 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_8 <= _GEN_4375;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_9 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_9 <= _GEN_4376;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_10 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_10 <= _GEN_4377;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_11 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_11 <= _GEN_4378;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_12 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_12 <= _GEN_4379;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_13 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_13 <= _GEN_4380;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_14 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_14 <= _GEN_4381;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_15 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_15 <= _GEN_4382;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_16 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_16 <= _GEN_4383;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_17 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_17 <= _GEN_4384;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_18 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_18 <= _GEN_4385;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_19 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_19 <= _GEN_4386;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_20 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_20 <= _GEN_4387;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_21 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_21 <= _GEN_4388;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_22 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_22 <= _GEN_4389;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_23 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_23 <= _GEN_4390;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_24 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_24 <= _GEN_4391;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_25 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_25 <= _GEN_4392;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_26 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_26 <= _GEN_4393;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_27 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_27 <= _GEN_4394;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_28 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_28 <= _GEN_4395;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_29 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_29 <= _GEN_4396;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_30 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_30 <= _GEN_4397;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_31 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_31 <= _GEN_4398;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_32 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_32 <= _GEN_4399;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_33 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_33 <= _GEN_4400;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_34 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_34 <= _GEN_4401;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_35 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_35 <= _GEN_4402;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_36 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_36 <= _GEN_4403;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_37 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_37 <= _GEN_4404;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_38 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_38 <= _GEN_4405;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_39 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_39 <= _GEN_4406;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_40 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_40 <= _GEN_4407;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_41 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_41 <= _GEN_4408;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_42 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_42 <= _GEN_4409;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_43 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_43 <= _GEN_4410;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_44 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_44 <= _GEN_4411;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_45 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_45 <= _GEN_4412;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_46 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_46 <= _GEN_4413;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_47 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_47 <= _GEN_4414;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_48 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_48 <= _GEN_4415;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_49 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_49 <= _GEN_4416;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_50 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_50 <= _GEN_4417;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_51 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_51 <= _GEN_4418;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_52 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_52 <= _GEN_4419;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_53 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_53 <= _GEN_4420;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_54 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_54 <= _GEN_4421;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_55 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_55 <= _GEN_4422;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_56 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_56 <= _GEN_4423;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_57 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_57 <= _GEN_4424;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_58 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_58 <= _GEN_4425;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_59 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_59 <= _GEN_4426;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_60 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_60 <= _GEN_4427;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_61 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_61 <= _GEN_4428;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_62 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_62 <= _GEN_4429;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_63 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_63 <= _GEN_4430;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_64 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_64 <= _GEN_4431;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_65 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_65 <= _GEN_4432;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_66 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_66 <= _GEN_4433;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_67 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_67 <= _GEN_4434;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_68 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_68 <= _GEN_4435;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_69 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_69 <= _GEN_4436;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_70 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_70 <= _GEN_4437;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_71 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_71 <= _GEN_4438;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_72 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_72 <= _GEN_4439;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_73 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_73 <= _GEN_4440;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_74 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_74 <= _GEN_4441;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_75 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_75 <= _GEN_4442;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_76 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_76 <= _GEN_4443;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_77 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_77 <= _GEN_4444;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_78 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_78 <= _GEN_4445;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_79 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_79 <= _GEN_4446;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_80 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_80 <= _GEN_4447;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_81 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_81 <= _GEN_4448;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_82 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_82 <= _GEN_4449;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_83 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_83 <= _GEN_4450;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_84 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_84 <= _GEN_4451;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_85 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_85 <= _GEN_4452;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_86 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_86 <= _GEN_4453;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_87 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_87 <= _GEN_4454;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_88 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_88 <= _GEN_4455;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_89 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_89 <= _GEN_4456;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_90 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_90 <= _GEN_4457;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_91 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_91 <= _GEN_4458;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_92 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_92 <= _GEN_4459;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_93 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_93 <= _GEN_4460;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_94 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_94 <= _GEN_4461;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_95 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_95 <= _GEN_4462;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_96 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_96 <= _GEN_4463;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_97 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_97 <= _GEN_4464;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_98 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_98 <= _GEN_4465;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_99 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_99 <= _GEN_4466;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_100 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_100 <= _GEN_4467;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_101 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_101 <= _GEN_4468;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_102 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_102 <= _GEN_4469;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_103 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_103 <= _GEN_4470;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_104 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_104 <= _GEN_4471;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_105 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_105 <= _GEN_4472;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_106 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_106 <= _GEN_4473;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_107 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_107 <= _GEN_4474;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_108 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_108 <= _GEN_4475;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_109 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_109 <= _GEN_4476;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_110 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_110 <= _GEN_4477;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_111 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_111 <= _GEN_4478;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_112 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_112 <= _GEN_4479;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_113 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_113 <= _GEN_4480;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_114 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_114 <= _GEN_4481;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_115 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_115 <= _GEN_4482;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_116 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_116 <= _GEN_4483;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_117 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_117 <= _GEN_4484;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_118 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_118 <= _GEN_4485;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_119 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_119 <= _GEN_4486;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_120 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_120 <= _GEN_4487;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_121 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_121 <= _GEN_4488;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_122 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_122 <= _GEN_4489;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_123 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_123 <= _GEN_4490;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_124 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_124 <= _GEN_4491;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_125 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_125 <= _GEN_4492;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_126 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_126 <= _GEN_4493;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 17:24]
      ram_0_127 <= 64'h0; // @[i_cache.scala 17:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_0_127 <= _GEN_4494;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_0 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_0 <= _GEN_4752;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_1 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_1 <= _GEN_4753;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_2 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_2 <= _GEN_4754;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_3 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_3 <= _GEN_4755;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_4 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_4 <= _GEN_4756;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_5 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_5 <= _GEN_4757;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_6 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_6 <= _GEN_4758;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_7 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_7 <= _GEN_4759;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_8 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_8 <= _GEN_4760;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_9 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_9 <= _GEN_4761;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_10 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_10 <= _GEN_4762;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_11 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_11 <= _GEN_4763;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_12 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_12 <= _GEN_4764;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_13 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_13 <= _GEN_4765;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_14 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_14 <= _GEN_4766;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_15 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_15 <= _GEN_4767;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_16 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_16 <= _GEN_4768;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_17 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_17 <= _GEN_4769;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_18 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_18 <= _GEN_4770;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_19 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_19 <= _GEN_4771;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_20 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_20 <= _GEN_4772;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_21 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_21 <= _GEN_4773;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_22 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_22 <= _GEN_4774;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_23 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_23 <= _GEN_4775;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_24 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_24 <= _GEN_4776;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_25 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_25 <= _GEN_4777;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_26 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_26 <= _GEN_4778;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_27 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_27 <= _GEN_4779;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_28 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_28 <= _GEN_4780;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_29 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_29 <= _GEN_4781;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_30 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_30 <= _GEN_4782;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_31 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_31 <= _GEN_4783;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_32 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_32 <= _GEN_4784;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_33 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_33 <= _GEN_4785;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_34 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_34 <= _GEN_4786;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_35 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_35 <= _GEN_4787;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_36 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_36 <= _GEN_4788;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_37 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_37 <= _GEN_4789;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_38 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_38 <= _GEN_4790;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_39 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_39 <= _GEN_4791;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_40 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_40 <= _GEN_4792;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_41 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_41 <= _GEN_4793;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_42 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_42 <= _GEN_4794;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_43 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_43 <= _GEN_4795;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_44 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_44 <= _GEN_4796;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_45 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_45 <= _GEN_4797;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_46 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_46 <= _GEN_4798;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_47 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_47 <= _GEN_4799;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_48 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_48 <= _GEN_4800;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_49 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_49 <= _GEN_4801;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_50 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_50 <= _GEN_4802;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_51 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_51 <= _GEN_4803;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_52 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_52 <= _GEN_4804;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_53 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_53 <= _GEN_4805;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_54 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_54 <= _GEN_4806;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_55 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_55 <= _GEN_4807;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_56 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_56 <= _GEN_4808;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_57 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_57 <= _GEN_4809;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_58 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_58 <= _GEN_4810;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_59 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_59 <= _GEN_4811;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_60 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_60 <= _GEN_4812;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_61 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_61 <= _GEN_4813;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_62 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_62 <= _GEN_4814;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_63 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_63 <= _GEN_4815;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_64 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_64 <= _GEN_4816;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_65 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_65 <= _GEN_4817;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_66 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_66 <= _GEN_4818;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_67 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_67 <= _GEN_4819;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_68 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_68 <= _GEN_4820;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_69 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_69 <= _GEN_4821;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_70 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_70 <= _GEN_4822;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_71 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_71 <= _GEN_4823;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_72 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_72 <= _GEN_4824;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_73 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_73 <= _GEN_4825;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_74 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_74 <= _GEN_4826;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_75 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_75 <= _GEN_4827;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_76 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_76 <= _GEN_4828;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_77 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_77 <= _GEN_4829;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_78 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_78 <= _GEN_4830;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_79 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_79 <= _GEN_4831;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_80 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_80 <= _GEN_4832;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_81 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_81 <= _GEN_4833;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_82 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_82 <= _GEN_4834;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_83 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_83 <= _GEN_4835;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_84 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_84 <= _GEN_4836;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_85 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_85 <= _GEN_4837;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_86 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_86 <= _GEN_4838;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_87 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_87 <= _GEN_4839;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_88 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_88 <= _GEN_4840;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_89 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_89 <= _GEN_4841;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_90 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_90 <= _GEN_4842;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_91 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_91 <= _GEN_4843;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_92 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_92 <= _GEN_4844;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_93 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_93 <= _GEN_4845;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_94 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_94 <= _GEN_4846;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_95 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_95 <= _GEN_4847;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_96 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_96 <= _GEN_4848;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_97 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_97 <= _GEN_4849;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_98 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_98 <= _GEN_4850;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_99 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_99 <= _GEN_4851;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_100 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_100 <= _GEN_4852;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_101 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_101 <= _GEN_4853;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_102 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_102 <= _GEN_4854;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_103 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_103 <= _GEN_4855;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_104 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_104 <= _GEN_4856;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_105 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_105 <= _GEN_4857;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_106 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_106 <= _GEN_4858;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_107 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_107 <= _GEN_4859;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_108 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_108 <= _GEN_4860;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_109 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_109 <= _GEN_4861;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_110 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_110 <= _GEN_4862;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_111 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_111 <= _GEN_4863;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_112 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_112 <= _GEN_4864;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_113 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_113 <= _GEN_4865;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_114 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_114 <= _GEN_4866;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_115 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_115 <= _GEN_4867;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_116 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_116 <= _GEN_4868;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_117 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_117 <= _GEN_4869;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_118 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_118 <= _GEN_4870;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_119 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_119 <= _GEN_4871;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_120 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_120 <= _GEN_4872;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_121 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_121 <= _GEN_4873;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_122 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_122 <= _GEN_4874;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_123 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_123 <= _GEN_4875;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_124 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_124 <= _GEN_4876;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_125 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_125 <= _GEN_4877;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_126 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_126 <= _GEN_4878;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 18:24]
      ram_1_127 <= 64'h0; // @[i_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          ram_1_127 <= _GEN_4879;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_0 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_0 <= _GEN_4495;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_1 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_1 <= _GEN_4496;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_2 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_2 <= _GEN_4497;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_3 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_3 <= _GEN_4498;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_4 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_4 <= _GEN_4499;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_5 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_5 <= _GEN_4500;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_6 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_6 <= _GEN_4501;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_7 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_7 <= _GEN_4502;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_8 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_8 <= _GEN_4503;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_9 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_9 <= _GEN_4504;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_10 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_10 <= _GEN_4505;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_11 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_11 <= _GEN_4506;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_12 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_12 <= _GEN_4507;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_13 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_13 <= _GEN_4508;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_14 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_14 <= _GEN_4509;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_15 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_15 <= _GEN_4510;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_16 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_16 <= _GEN_4511;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_17 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_17 <= _GEN_4512;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_18 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_18 <= _GEN_4513;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_19 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_19 <= _GEN_4514;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_20 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_20 <= _GEN_4515;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_21 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_21 <= _GEN_4516;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_22 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_22 <= _GEN_4517;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_23 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_23 <= _GEN_4518;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_24 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_24 <= _GEN_4519;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_25 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_25 <= _GEN_4520;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_26 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_26 <= _GEN_4521;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_27 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_27 <= _GEN_4522;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_28 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_28 <= _GEN_4523;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_29 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_29 <= _GEN_4524;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_30 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_30 <= _GEN_4525;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_31 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_31 <= _GEN_4526;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_32 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_32 <= _GEN_4527;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_33 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_33 <= _GEN_4528;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_34 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_34 <= _GEN_4529;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_35 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_35 <= _GEN_4530;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_36 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_36 <= _GEN_4531;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_37 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_37 <= _GEN_4532;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_38 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_38 <= _GEN_4533;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_39 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_39 <= _GEN_4534;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_40 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_40 <= _GEN_4535;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_41 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_41 <= _GEN_4536;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_42 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_42 <= _GEN_4537;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_43 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_43 <= _GEN_4538;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_44 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_44 <= _GEN_4539;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_45 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_45 <= _GEN_4540;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_46 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_46 <= _GEN_4541;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_47 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_47 <= _GEN_4542;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_48 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_48 <= _GEN_4543;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_49 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_49 <= _GEN_4544;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_50 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_50 <= _GEN_4545;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_51 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_51 <= _GEN_4546;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_52 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_52 <= _GEN_4547;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_53 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_53 <= _GEN_4548;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_54 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_54 <= _GEN_4549;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_55 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_55 <= _GEN_4550;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_56 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_56 <= _GEN_4551;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_57 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_57 <= _GEN_4552;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_58 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_58 <= _GEN_4553;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_59 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_59 <= _GEN_4554;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_60 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_60 <= _GEN_4555;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_61 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_61 <= _GEN_4556;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_62 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_62 <= _GEN_4557;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_63 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_63 <= _GEN_4558;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_64 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_64 <= _GEN_4559;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_65 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_65 <= _GEN_4560;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_66 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_66 <= _GEN_4561;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_67 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_67 <= _GEN_4562;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_68 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_68 <= _GEN_4563;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_69 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_69 <= _GEN_4564;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_70 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_70 <= _GEN_4565;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_71 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_71 <= _GEN_4566;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_72 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_72 <= _GEN_4567;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_73 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_73 <= _GEN_4568;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_74 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_74 <= _GEN_4569;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_75 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_75 <= _GEN_4570;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_76 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_76 <= _GEN_4571;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_77 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_77 <= _GEN_4572;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_78 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_78 <= _GEN_4573;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_79 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_79 <= _GEN_4574;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_80 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_80 <= _GEN_4575;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_81 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_81 <= _GEN_4576;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_82 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_82 <= _GEN_4577;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_83 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_83 <= _GEN_4578;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_84 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_84 <= _GEN_4579;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_85 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_85 <= _GEN_4580;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_86 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_86 <= _GEN_4581;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_87 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_87 <= _GEN_4582;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_88 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_88 <= _GEN_4583;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_89 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_89 <= _GEN_4584;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_90 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_90 <= _GEN_4585;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_91 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_91 <= _GEN_4586;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_92 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_92 <= _GEN_4587;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_93 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_93 <= _GEN_4588;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_94 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_94 <= _GEN_4589;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_95 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_95 <= _GEN_4590;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_96 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_96 <= _GEN_4591;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_97 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_97 <= _GEN_4592;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_98 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_98 <= _GEN_4593;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_99 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_99 <= _GEN_4594;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_100 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_100 <= _GEN_4595;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_101 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_101 <= _GEN_4596;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_102 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_102 <= _GEN_4597;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_103 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_103 <= _GEN_4598;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_104 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_104 <= _GEN_4599;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_105 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_105 <= _GEN_4600;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_106 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_106 <= _GEN_4601;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_107 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_107 <= _GEN_4602;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_108 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_108 <= _GEN_4603;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_109 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_109 <= _GEN_4604;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_110 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_110 <= _GEN_4605;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_111 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_111 <= _GEN_4606;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_112 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_112 <= _GEN_4607;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_113 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_113 <= _GEN_4608;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_114 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_114 <= _GEN_4609;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_115 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_115 <= _GEN_4610;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_116 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_116 <= _GEN_4611;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_117 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_117 <= _GEN_4612;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_118 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_118 <= _GEN_4613;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_119 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_119 <= _GEN_4614;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_120 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_120 <= _GEN_4615;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_121 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_121 <= _GEN_4616;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_122 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_122 <= _GEN_4617;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_123 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_123 <= _GEN_4618;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_124 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_124 <= _GEN_4619;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_125 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_125 <= _GEN_4620;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_126 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_126 <= _GEN_4621;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      tag_0_127 <= 32'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_0_127 <= _GEN_4622;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_0 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_0 <= _GEN_4880;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_1 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_1 <= _GEN_4881;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_2 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_2 <= _GEN_4882;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_3 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_3 <= _GEN_4883;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_4 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_4 <= _GEN_4884;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_5 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_5 <= _GEN_4885;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_6 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_6 <= _GEN_4886;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_7 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_7 <= _GEN_4887;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_8 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_8 <= _GEN_4888;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_9 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_9 <= _GEN_4889;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_10 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_10 <= _GEN_4890;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_11 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_11 <= _GEN_4891;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_12 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_12 <= _GEN_4892;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_13 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_13 <= _GEN_4893;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_14 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_14 <= _GEN_4894;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_15 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_15 <= _GEN_4895;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_16 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_16 <= _GEN_4896;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_17 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_17 <= _GEN_4897;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_18 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_18 <= _GEN_4898;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_19 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_19 <= _GEN_4899;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_20 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_20 <= _GEN_4900;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_21 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_21 <= _GEN_4901;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_22 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_22 <= _GEN_4902;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_23 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_23 <= _GEN_4903;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_24 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_24 <= _GEN_4904;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_25 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_25 <= _GEN_4905;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_26 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_26 <= _GEN_4906;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_27 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_27 <= _GEN_4907;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_28 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_28 <= _GEN_4908;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_29 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_29 <= _GEN_4909;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_30 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_30 <= _GEN_4910;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_31 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_31 <= _GEN_4911;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_32 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_32 <= _GEN_4912;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_33 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_33 <= _GEN_4913;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_34 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_34 <= _GEN_4914;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_35 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_35 <= _GEN_4915;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_36 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_36 <= _GEN_4916;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_37 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_37 <= _GEN_4917;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_38 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_38 <= _GEN_4918;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_39 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_39 <= _GEN_4919;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_40 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_40 <= _GEN_4920;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_41 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_41 <= _GEN_4921;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_42 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_42 <= _GEN_4922;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_43 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_43 <= _GEN_4923;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_44 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_44 <= _GEN_4924;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_45 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_45 <= _GEN_4925;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_46 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_46 <= _GEN_4926;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_47 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_47 <= _GEN_4927;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_48 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_48 <= _GEN_4928;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_49 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_49 <= _GEN_4929;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_50 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_50 <= _GEN_4930;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_51 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_51 <= _GEN_4931;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_52 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_52 <= _GEN_4932;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_53 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_53 <= _GEN_4933;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_54 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_54 <= _GEN_4934;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_55 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_55 <= _GEN_4935;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_56 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_56 <= _GEN_4936;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_57 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_57 <= _GEN_4937;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_58 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_58 <= _GEN_4938;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_59 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_59 <= _GEN_4939;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_60 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_60 <= _GEN_4940;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_61 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_61 <= _GEN_4941;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_62 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_62 <= _GEN_4942;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_63 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_63 <= _GEN_4943;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_64 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_64 <= _GEN_4944;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_65 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_65 <= _GEN_4945;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_66 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_66 <= _GEN_4946;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_67 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_67 <= _GEN_4947;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_68 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_68 <= _GEN_4948;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_69 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_69 <= _GEN_4949;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_70 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_70 <= _GEN_4950;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_71 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_71 <= _GEN_4951;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_72 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_72 <= _GEN_4952;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_73 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_73 <= _GEN_4953;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_74 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_74 <= _GEN_4954;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_75 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_75 <= _GEN_4955;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_76 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_76 <= _GEN_4956;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_77 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_77 <= _GEN_4957;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_78 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_78 <= _GEN_4958;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_79 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_79 <= _GEN_4959;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_80 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_80 <= _GEN_4960;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_81 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_81 <= _GEN_4961;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_82 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_82 <= _GEN_4962;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_83 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_83 <= _GEN_4963;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_84 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_84 <= _GEN_4964;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_85 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_85 <= _GEN_4965;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_86 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_86 <= _GEN_4966;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_87 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_87 <= _GEN_4967;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_88 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_88 <= _GEN_4968;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_89 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_89 <= _GEN_4969;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_90 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_90 <= _GEN_4970;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_91 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_91 <= _GEN_4971;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_92 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_92 <= _GEN_4972;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_93 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_93 <= _GEN_4973;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_94 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_94 <= _GEN_4974;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_95 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_95 <= _GEN_4975;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_96 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_96 <= _GEN_4976;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_97 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_97 <= _GEN_4977;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_98 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_98 <= _GEN_4978;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_99 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_99 <= _GEN_4979;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_100 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_100 <= _GEN_4980;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_101 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_101 <= _GEN_4981;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_102 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_102 <= _GEN_4982;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_103 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_103 <= _GEN_4983;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_104 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_104 <= _GEN_4984;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_105 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_105 <= _GEN_4985;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_106 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_106 <= _GEN_4986;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_107 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_107 <= _GEN_4987;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_108 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_108 <= _GEN_4988;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_109 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_109 <= _GEN_4989;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_110 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_110 <= _GEN_4990;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_111 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_111 <= _GEN_4991;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_112 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_112 <= _GEN_4992;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_113 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_113 <= _GEN_4993;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_114 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_114 <= _GEN_4994;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_115 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_115 <= _GEN_4995;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_116 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_116 <= _GEN_4996;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_117 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_117 <= _GEN_4997;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_118 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_118 <= _GEN_4998;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_119 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_119 <= _GEN_4999;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_120 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_120 <= _GEN_5000;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_121 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_121 <= _GEN_5001;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_122 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_122 <= _GEN_5002;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_123 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_123 <= _GEN_5003;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_124 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_124 <= _GEN_5004;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_125 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_125 <= _GEN_5005;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_126 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_126 <= _GEN_5006;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      tag_1_127 <= 32'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          tag_1_127 <= _GEN_5007;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_0 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_0 <= _GEN_4623;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_1 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_1 <= _GEN_4624;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_2 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_2 <= _GEN_4625;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_3 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_3 <= _GEN_4626;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_4 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_4 <= _GEN_4627;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_5 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_5 <= _GEN_4628;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_6 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_6 <= _GEN_4629;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_7 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_7 <= _GEN_4630;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_8 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_8 <= _GEN_4631;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_9 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_9 <= _GEN_4632;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_10 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_10 <= _GEN_4633;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_11 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_11 <= _GEN_4634;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_12 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_12 <= _GEN_4635;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_13 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_13 <= _GEN_4636;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_14 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_14 <= _GEN_4637;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_15 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_15 <= _GEN_4638;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_16 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_16 <= _GEN_4639;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_17 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_17 <= _GEN_4640;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_18 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_18 <= _GEN_4641;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_19 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_19 <= _GEN_4642;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_20 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_20 <= _GEN_4643;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_21 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_21 <= _GEN_4644;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_22 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_22 <= _GEN_4645;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_23 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_23 <= _GEN_4646;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_24 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_24 <= _GEN_4647;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_25 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_25 <= _GEN_4648;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_26 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_26 <= _GEN_4649;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_27 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_27 <= _GEN_4650;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_28 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_28 <= _GEN_4651;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_29 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_29 <= _GEN_4652;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_30 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_30 <= _GEN_4653;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_31 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_31 <= _GEN_4654;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_32 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_32 <= _GEN_4655;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_33 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_33 <= _GEN_4656;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_34 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_34 <= _GEN_4657;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_35 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_35 <= _GEN_4658;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_36 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_36 <= _GEN_4659;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_37 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_37 <= _GEN_4660;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_38 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_38 <= _GEN_4661;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_39 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_39 <= _GEN_4662;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_40 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_40 <= _GEN_4663;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_41 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_41 <= _GEN_4664;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_42 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_42 <= _GEN_4665;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_43 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_43 <= _GEN_4666;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_44 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_44 <= _GEN_4667;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_45 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_45 <= _GEN_4668;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_46 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_46 <= _GEN_4669;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_47 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_47 <= _GEN_4670;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_48 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_48 <= _GEN_4671;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_49 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_49 <= _GEN_4672;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_50 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_50 <= _GEN_4673;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_51 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_51 <= _GEN_4674;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_52 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_52 <= _GEN_4675;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_53 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_53 <= _GEN_4676;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_54 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_54 <= _GEN_4677;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_55 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_55 <= _GEN_4678;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_56 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_56 <= _GEN_4679;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_57 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_57 <= _GEN_4680;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_58 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_58 <= _GEN_4681;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_59 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_59 <= _GEN_4682;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_60 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_60 <= _GEN_4683;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_61 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_61 <= _GEN_4684;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_62 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_62 <= _GEN_4685;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_63 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_63 <= _GEN_4686;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_64 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_64 <= _GEN_4687;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_65 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_65 <= _GEN_4688;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_66 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_66 <= _GEN_4689;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_67 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_67 <= _GEN_4690;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_68 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_68 <= _GEN_4691;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_69 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_69 <= _GEN_4692;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_70 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_70 <= _GEN_4693;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_71 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_71 <= _GEN_4694;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_72 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_72 <= _GEN_4695;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_73 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_73 <= _GEN_4696;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_74 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_74 <= _GEN_4697;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_75 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_75 <= _GEN_4698;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_76 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_76 <= _GEN_4699;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_77 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_77 <= _GEN_4700;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_78 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_78 <= _GEN_4701;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_79 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_79 <= _GEN_4702;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_80 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_80 <= _GEN_4703;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_81 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_81 <= _GEN_4704;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_82 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_82 <= _GEN_4705;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_83 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_83 <= _GEN_4706;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_84 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_84 <= _GEN_4707;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_85 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_85 <= _GEN_4708;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_86 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_86 <= _GEN_4709;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_87 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_87 <= _GEN_4710;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_88 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_88 <= _GEN_4711;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_89 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_89 <= _GEN_4712;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_90 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_90 <= _GEN_4713;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_91 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_91 <= _GEN_4714;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_92 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_92 <= _GEN_4715;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_93 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_93 <= _GEN_4716;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_94 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_94 <= _GEN_4717;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_95 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_95 <= _GEN_4718;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_96 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_96 <= _GEN_4719;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_97 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_97 <= _GEN_4720;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_98 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_98 <= _GEN_4721;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_99 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_99 <= _GEN_4722;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_100 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_100 <= _GEN_4723;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_101 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_101 <= _GEN_4724;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_102 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_102 <= _GEN_4725;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_103 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_103 <= _GEN_4726;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_104 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_104 <= _GEN_4727;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_105 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_105 <= _GEN_4728;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_106 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_106 <= _GEN_4729;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_107 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_107 <= _GEN_4730;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_108 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_108 <= _GEN_4731;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_109 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_109 <= _GEN_4732;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_110 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_110 <= _GEN_4733;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_111 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_111 <= _GEN_4734;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_112 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_112 <= _GEN_4735;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_113 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_113 <= _GEN_4736;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_114 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_114 <= _GEN_4737;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_115 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_115 <= _GEN_4738;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_116 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_116 <= _GEN_4739;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_117 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_117 <= _GEN_4740;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_118 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_118 <= _GEN_4741;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_119 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_119 <= _GEN_4742;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_120 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_120 <= _GEN_4743;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_121 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_121 <= _GEN_4744;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_122 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_122 <= _GEN_4745;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_123 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_123 <= _GEN_4746;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_124 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_124 <= _GEN_4747;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_125 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_125 <= _GEN_4748;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_126 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_126 <= _GEN_4749;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:26]
      valid_0_127 <= 1'h0; // @[i_cache.scala 21:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_0_127 <= _GEN_4750;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_0 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_0 <= _GEN_5008;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_1 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_1 <= _GEN_5009;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_2 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_2 <= _GEN_5010;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_3 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_3 <= _GEN_5011;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_4 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_4 <= _GEN_5012;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_5 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_5 <= _GEN_5013;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_6 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_6 <= _GEN_5014;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_7 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_7 <= _GEN_5015;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_8 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_8 <= _GEN_5016;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_9 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_9 <= _GEN_5017;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_10 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_10 <= _GEN_5018;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_11 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_11 <= _GEN_5019;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_12 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_12 <= _GEN_5020;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_13 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_13 <= _GEN_5021;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_14 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_14 <= _GEN_5022;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_15 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_15 <= _GEN_5023;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_16 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_16 <= _GEN_5024;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_17 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_17 <= _GEN_5025;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_18 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_18 <= _GEN_5026;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_19 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_19 <= _GEN_5027;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_20 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_20 <= _GEN_5028;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_21 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_21 <= _GEN_5029;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_22 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_22 <= _GEN_5030;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_23 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_23 <= _GEN_5031;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_24 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_24 <= _GEN_5032;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_25 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_25 <= _GEN_5033;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_26 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_26 <= _GEN_5034;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_27 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_27 <= _GEN_5035;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_28 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_28 <= _GEN_5036;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_29 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_29 <= _GEN_5037;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_30 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_30 <= _GEN_5038;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_31 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_31 <= _GEN_5039;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_32 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_32 <= _GEN_5040;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_33 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_33 <= _GEN_5041;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_34 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_34 <= _GEN_5042;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_35 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_35 <= _GEN_5043;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_36 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_36 <= _GEN_5044;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_37 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_37 <= _GEN_5045;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_38 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_38 <= _GEN_5046;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_39 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_39 <= _GEN_5047;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_40 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_40 <= _GEN_5048;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_41 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_41 <= _GEN_5049;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_42 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_42 <= _GEN_5050;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_43 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_43 <= _GEN_5051;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_44 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_44 <= _GEN_5052;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_45 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_45 <= _GEN_5053;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_46 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_46 <= _GEN_5054;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_47 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_47 <= _GEN_5055;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_48 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_48 <= _GEN_5056;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_49 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_49 <= _GEN_5057;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_50 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_50 <= _GEN_5058;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_51 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_51 <= _GEN_5059;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_52 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_52 <= _GEN_5060;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_53 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_53 <= _GEN_5061;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_54 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_54 <= _GEN_5062;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_55 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_55 <= _GEN_5063;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_56 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_56 <= _GEN_5064;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_57 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_57 <= _GEN_5065;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_58 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_58 <= _GEN_5066;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_59 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_59 <= _GEN_5067;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_60 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_60 <= _GEN_5068;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_61 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_61 <= _GEN_5069;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_62 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_62 <= _GEN_5070;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_63 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_63 <= _GEN_5071;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_64 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_64 <= _GEN_5072;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_65 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_65 <= _GEN_5073;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_66 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_66 <= _GEN_5074;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_67 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_67 <= _GEN_5075;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_68 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_68 <= _GEN_5076;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_69 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_69 <= _GEN_5077;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_70 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_70 <= _GEN_5078;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_71 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_71 <= _GEN_5079;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_72 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_72 <= _GEN_5080;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_73 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_73 <= _GEN_5081;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_74 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_74 <= _GEN_5082;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_75 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_75 <= _GEN_5083;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_76 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_76 <= _GEN_5084;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_77 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_77 <= _GEN_5085;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_78 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_78 <= _GEN_5086;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_79 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_79 <= _GEN_5087;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_80 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_80 <= _GEN_5088;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_81 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_81 <= _GEN_5089;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_82 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_82 <= _GEN_5090;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_83 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_83 <= _GEN_5091;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_84 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_84 <= _GEN_5092;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_85 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_85 <= _GEN_5093;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_86 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_86 <= _GEN_5094;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_87 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_87 <= _GEN_5095;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_88 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_88 <= _GEN_5096;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_89 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_89 <= _GEN_5097;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_90 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_90 <= _GEN_5098;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_91 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_91 <= _GEN_5099;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_92 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_92 <= _GEN_5100;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_93 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_93 <= _GEN_5101;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_94 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_94 <= _GEN_5102;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_95 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_95 <= _GEN_5103;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_96 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_96 <= _GEN_5104;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_97 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_97 <= _GEN_5105;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_98 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_98 <= _GEN_5106;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_99 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_99 <= _GEN_5107;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_100 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_100 <= _GEN_5108;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_101 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_101 <= _GEN_5109;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_102 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_102 <= _GEN_5110;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_103 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_103 <= _GEN_5111;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_104 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_104 <= _GEN_5112;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_105 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_105 <= _GEN_5113;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_106 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_106 <= _GEN_5114;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_107 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_107 <= _GEN_5115;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_108 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_108 <= _GEN_5116;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_109 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_109 <= _GEN_5117;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_110 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_110 <= _GEN_5118;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_111 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_111 <= _GEN_5119;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_112 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_112 <= _GEN_5120;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_113 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_113 <= _GEN_5121;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_114 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_114 <= _GEN_5122;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_115 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_115 <= _GEN_5123;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_116 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_116 <= _GEN_5124;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_117 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_117 <= _GEN_5125;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_118 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_118 <= _GEN_5126;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_119 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_119 <= _GEN_5127;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_120 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_120 <= _GEN_5128;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_121 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_121 <= _GEN_5129;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_122 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_122 <= _GEN_5130;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_123 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_123 <= _GEN_5131;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_124 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_124 <= _GEN_5132;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_125 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_125 <= _GEN_5133;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_126 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_126 <= _GEN_5134;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:26]
      valid_1_127 <= 1'h0; // @[i_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          valid_1_127 <= _GEN_5135;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:27]
      way0_hit <= 1'h0; // @[i_cache.scala 23:27]
    end else begin
      way0_hit <= _T_2;
    end
    if (reset) begin // @[i_cache.scala 24:27]
      way1_hit <= 1'h0; // @[i_cache.scala 24:27]
    end else begin
      way1_hit <= _T_5;
    end
    if (reset) begin // @[i_cache.scala 26:28]
      unuse_way <= 2'h0; // @[i_cache.scala 26:28]
    end else if (~_GEN_255) begin // @[i_cache.scala 45:31]
      unuse_way <= 2'h1; // @[i_cache.scala 46:19]
    end else if (~_GEN_512) begin // @[i_cache.scala 47:37]
      unuse_way <= 2'h2; // @[i_cache.scala 48:19]
    end else begin
      unuse_way <= 2'h0; // @[i_cache.scala 50:19]
    end
    if (reset) begin // @[i_cache.scala 27:31]
      receive_data <= 64'h0; // @[i_cache.scala 27:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (3'h2 == state) begin // @[i_cache.scala 55:18]
          receive_data <= _GEN_521;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:24]
      quene <= 1'h0; // @[i_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 55:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 55:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 55:18]
          quene <= _GEN_4751;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 53:24]
      state <= 3'h0; // @[i_cache.scala 53:24]
    end else if (3'h0 == state) begin // @[i_cache.scala 55:18]
      if (io_from_ifu_arvalid) begin // @[i_cache.scala 57:38]
        state <= 3'h1; // @[i_cache.scala 58:23]
      end
    end else if (3'h1 == state) begin // @[i_cache.scala 55:18]
      if (way0_hit) begin // @[i_cache.scala 63:27]
        state <= _GEN_517;
      end else begin
        state <= _GEN_518;
      end
    end else if (3'h2 == state) begin // @[i_cache.scala 55:18]
      state <= _GEN_520;
    end else begin
      state <= _GEN_4366;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ram_0_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ram_0_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ram_0_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ram_0_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ram_0_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ram_0_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ram_0_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ram_0_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  ram_0_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  ram_0_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  ram_0_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  ram_0_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  ram_0_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  ram_0_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  ram_0_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  ram_0_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  ram_0_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  ram_0_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  ram_0_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  ram_0_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  ram_0_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  ram_0_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  ram_0_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  ram_0_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  ram_0_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  ram_0_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  ram_0_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  ram_0_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  ram_0_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  ram_0_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  ram_0_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  ram_0_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  ram_0_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  ram_0_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  ram_0_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  ram_0_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  ram_0_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  ram_0_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  ram_0_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  ram_0_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  ram_0_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  ram_0_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  ram_0_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  ram_0_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  ram_0_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  ram_0_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  ram_0_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  ram_0_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  ram_0_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  ram_0_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  ram_0_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  ram_0_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  ram_0_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  ram_0_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  ram_0_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  ram_0_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  ram_0_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  ram_0_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  ram_0_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  ram_0_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  ram_0_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  ram_0_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  ram_0_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  ram_0_63 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  ram_0_64 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  ram_0_65 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  ram_0_66 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  ram_0_67 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  ram_0_68 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  ram_0_69 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  ram_0_70 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  ram_0_71 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  ram_0_72 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  ram_0_73 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  ram_0_74 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  ram_0_75 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  ram_0_76 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  ram_0_77 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  ram_0_78 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  ram_0_79 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  ram_0_80 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  ram_0_81 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  ram_0_82 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  ram_0_83 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  ram_0_84 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  ram_0_85 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  ram_0_86 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  ram_0_87 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  ram_0_88 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  ram_0_89 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  ram_0_90 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  ram_0_91 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  ram_0_92 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  ram_0_93 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  ram_0_94 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  ram_0_95 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  ram_0_96 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  ram_0_97 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  ram_0_98 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  ram_0_99 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  ram_0_100 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  ram_0_101 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  ram_0_102 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  ram_0_103 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  ram_0_104 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  ram_0_105 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  ram_0_106 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  ram_0_107 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  ram_0_108 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  ram_0_109 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  ram_0_110 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  ram_0_111 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  ram_0_112 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  ram_0_113 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  ram_0_114 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  ram_0_115 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  ram_0_116 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  ram_0_117 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  ram_0_118 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  ram_0_119 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  ram_0_120 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  ram_0_121 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  ram_0_122 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  ram_0_123 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  ram_0_124 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  ram_0_125 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  ram_0_126 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  ram_0_127 = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  ram_1_0 = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  ram_1_1 = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  ram_1_2 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  ram_1_3 = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  ram_1_4 = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  ram_1_5 = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  ram_1_6 = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  ram_1_7 = _RAND_135[63:0];
  _RAND_136 = {2{`RANDOM}};
  ram_1_8 = _RAND_136[63:0];
  _RAND_137 = {2{`RANDOM}};
  ram_1_9 = _RAND_137[63:0];
  _RAND_138 = {2{`RANDOM}};
  ram_1_10 = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  ram_1_11 = _RAND_139[63:0];
  _RAND_140 = {2{`RANDOM}};
  ram_1_12 = _RAND_140[63:0];
  _RAND_141 = {2{`RANDOM}};
  ram_1_13 = _RAND_141[63:0];
  _RAND_142 = {2{`RANDOM}};
  ram_1_14 = _RAND_142[63:0];
  _RAND_143 = {2{`RANDOM}};
  ram_1_15 = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  ram_1_16 = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  ram_1_17 = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  ram_1_18 = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  ram_1_19 = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  ram_1_20 = _RAND_148[63:0];
  _RAND_149 = {2{`RANDOM}};
  ram_1_21 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  ram_1_22 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  ram_1_23 = _RAND_151[63:0];
  _RAND_152 = {2{`RANDOM}};
  ram_1_24 = _RAND_152[63:0];
  _RAND_153 = {2{`RANDOM}};
  ram_1_25 = _RAND_153[63:0];
  _RAND_154 = {2{`RANDOM}};
  ram_1_26 = _RAND_154[63:0];
  _RAND_155 = {2{`RANDOM}};
  ram_1_27 = _RAND_155[63:0];
  _RAND_156 = {2{`RANDOM}};
  ram_1_28 = _RAND_156[63:0];
  _RAND_157 = {2{`RANDOM}};
  ram_1_29 = _RAND_157[63:0];
  _RAND_158 = {2{`RANDOM}};
  ram_1_30 = _RAND_158[63:0];
  _RAND_159 = {2{`RANDOM}};
  ram_1_31 = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  ram_1_32 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  ram_1_33 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  ram_1_34 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  ram_1_35 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  ram_1_36 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  ram_1_37 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  ram_1_38 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  ram_1_39 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  ram_1_40 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  ram_1_41 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  ram_1_42 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  ram_1_43 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  ram_1_44 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  ram_1_45 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  ram_1_46 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  ram_1_47 = _RAND_175[63:0];
  _RAND_176 = {2{`RANDOM}};
  ram_1_48 = _RAND_176[63:0];
  _RAND_177 = {2{`RANDOM}};
  ram_1_49 = _RAND_177[63:0];
  _RAND_178 = {2{`RANDOM}};
  ram_1_50 = _RAND_178[63:0];
  _RAND_179 = {2{`RANDOM}};
  ram_1_51 = _RAND_179[63:0];
  _RAND_180 = {2{`RANDOM}};
  ram_1_52 = _RAND_180[63:0];
  _RAND_181 = {2{`RANDOM}};
  ram_1_53 = _RAND_181[63:0];
  _RAND_182 = {2{`RANDOM}};
  ram_1_54 = _RAND_182[63:0];
  _RAND_183 = {2{`RANDOM}};
  ram_1_55 = _RAND_183[63:0];
  _RAND_184 = {2{`RANDOM}};
  ram_1_56 = _RAND_184[63:0];
  _RAND_185 = {2{`RANDOM}};
  ram_1_57 = _RAND_185[63:0];
  _RAND_186 = {2{`RANDOM}};
  ram_1_58 = _RAND_186[63:0];
  _RAND_187 = {2{`RANDOM}};
  ram_1_59 = _RAND_187[63:0];
  _RAND_188 = {2{`RANDOM}};
  ram_1_60 = _RAND_188[63:0];
  _RAND_189 = {2{`RANDOM}};
  ram_1_61 = _RAND_189[63:0];
  _RAND_190 = {2{`RANDOM}};
  ram_1_62 = _RAND_190[63:0];
  _RAND_191 = {2{`RANDOM}};
  ram_1_63 = _RAND_191[63:0];
  _RAND_192 = {2{`RANDOM}};
  ram_1_64 = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  ram_1_65 = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  ram_1_66 = _RAND_194[63:0];
  _RAND_195 = {2{`RANDOM}};
  ram_1_67 = _RAND_195[63:0];
  _RAND_196 = {2{`RANDOM}};
  ram_1_68 = _RAND_196[63:0];
  _RAND_197 = {2{`RANDOM}};
  ram_1_69 = _RAND_197[63:0];
  _RAND_198 = {2{`RANDOM}};
  ram_1_70 = _RAND_198[63:0];
  _RAND_199 = {2{`RANDOM}};
  ram_1_71 = _RAND_199[63:0];
  _RAND_200 = {2{`RANDOM}};
  ram_1_72 = _RAND_200[63:0];
  _RAND_201 = {2{`RANDOM}};
  ram_1_73 = _RAND_201[63:0];
  _RAND_202 = {2{`RANDOM}};
  ram_1_74 = _RAND_202[63:0];
  _RAND_203 = {2{`RANDOM}};
  ram_1_75 = _RAND_203[63:0];
  _RAND_204 = {2{`RANDOM}};
  ram_1_76 = _RAND_204[63:0];
  _RAND_205 = {2{`RANDOM}};
  ram_1_77 = _RAND_205[63:0];
  _RAND_206 = {2{`RANDOM}};
  ram_1_78 = _RAND_206[63:0];
  _RAND_207 = {2{`RANDOM}};
  ram_1_79 = _RAND_207[63:0];
  _RAND_208 = {2{`RANDOM}};
  ram_1_80 = _RAND_208[63:0];
  _RAND_209 = {2{`RANDOM}};
  ram_1_81 = _RAND_209[63:0];
  _RAND_210 = {2{`RANDOM}};
  ram_1_82 = _RAND_210[63:0];
  _RAND_211 = {2{`RANDOM}};
  ram_1_83 = _RAND_211[63:0];
  _RAND_212 = {2{`RANDOM}};
  ram_1_84 = _RAND_212[63:0];
  _RAND_213 = {2{`RANDOM}};
  ram_1_85 = _RAND_213[63:0];
  _RAND_214 = {2{`RANDOM}};
  ram_1_86 = _RAND_214[63:0];
  _RAND_215 = {2{`RANDOM}};
  ram_1_87 = _RAND_215[63:0];
  _RAND_216 = {2{`RANDOM}};
  ram_1_88 = _RAND_216[63:0];
  _RAND_217 = {2{`RANDOM}};
  ram_1_89 = _RAND_217[63:0];
  _RAND_218 = {2{`RANDOM}};
  ram_1_90 = _RAND_218[63:0];
  _RAND_219 = {2{`RANDOM}};
  ram_1_91 = _RAND_219[63:0];
  _RAND_220 = {2{`RANDOM}};
  ram_1_92 = _RAND_220[63:0];
  _RAND_221 = {2{`RANDOM}};
  ram_1_93 = _RAND_221[63:0];
  _RAND_222 = {2{`RANDOM}};
  ram_1_94 = _RAND_222[63:0];
  _RAND_223 = {2{`RANDOM}};
  ram_1_95 = _RAND_223[63:0];
  _RAND_224 = {2{`RANDOM}};
  ram_1_96 = _RAND_224[63:0];
  _RAND_225 = {2{`RANDOM}};
  ram_1_97 = _RAND_225[63:0];
  _RAND_226 = {2{`RANDOM}};
  ram_1_98 = _RAND_226[63:0];
  _RAND_227 = {2{`RANDOM}};
  ram_1_99 = _RAND_227[63:0];
  _RAND_228 = {2{`RANDOM}};
  ram_1_100 = _RAND_228[63:0];
  _RAND_229 = {2{`RANDOM}};
  ram_1_101 = _RAND_229[63:0];
  _RAND_230 = {2{`RANDOM}};
  ram_1_102 = _RAND_230[63:0];
  _RAND_231 = {2{`RANDOM}};
  ram_1_103 = _RAND_231[63:0];
  _RAND_232 = {2{`RANDOM}};
  ram_1_104 = _RAND_232[63:0];
  _RAND_233 = {2{`RANDOM}};
  ram_1_105 = _RAND_233[63:0];
  _RAND_234 = {2{`RANDOM}};
  ram_1_106 = _RAND_234[63:0];
  _RAND_235 = {2{`RANDOM}};
  ram_1_107 = _RAND_235[63:0];
  _RAND_236 = {2{`RANDOM}};
  ram_1_108 = _RAND_236[63:0];
  _RAND_237 = {2{`RANDOM}};
  ram_1_109 = _RAND_237[63:0];
  _RAND_238 = {2{`RANDOM}};
  ram_1_110 = _RAND_238[63:0];
  _RAND_239 = {2{`RANDOM}};
  ram_1_111 = _RAND_239[63:0];
  _RAND_240 = {2{`RANDOM}};
  ram_1_112 = _RAND_240[63:0];
  _RAND_241 = {2{`RANDOM}};
  ram_1_113 = _RAND_241[63:0];
  _RAND_242 = {2{`RANDOM}};
  ram_1_114 = _RAND_242[63:0];
  _RAND_243 = {2{`RANDOM}};
  ram_1_115 = _RAND_243[63:0];
  _RAND_244 = {2{`RANDOM}};
  ram_1_116 = _RAND_244[63:0];
  _RAND_245 = {2{`RANDOM}};
  ram_1_117 = _RAND_245[63:0];
  _RAND_246 = {2{`RANDOM}};
  ram_1_118 = _RAND_246[63:0];
  _RAND_247 = {2{`RANDOM}};
  ram_1_119 = _RAND_247[63:0];
  _RAND_248 = {2{`RANDOM}};
  ram_1_120 = _RAND_248[63:0];
  _RAND_249 = {2{`RANDOM}};
  ram_1_121 = _RAND_249[63:0];
  _RAND_250 = {2{`RANDOM}};
  ram_1_122 = _RAND_250[63:0];
  _RAND_251 = {2{`RANDOM}};
  ram_1_123 = _RAND_251[63:0];
  _RAND_252 = {2{`RANDOM}};
  ram_1_124 = _RAND_252[63:0];
  _RAND_253 = {2{`RANDOM}};
  ram_1_125 = _RAND_253[63:0];
  _RAND_254 = {2{`RANDOM}};
  ram_1_126 = _RAND_254[63:0];
  _RAND_255 = {2{`RANDOM}};
  ram_1_127 = _RAND_255[63:0];
  _RAND_256 = {1{`RANDOM}};
  tag_0_0 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  tag_0_1 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  tag_0_2 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  tag_0_3 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  tag_0_4 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  tag_0_5 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  tag_0_6 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  tag_0_7 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  tag_0_8 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  tag_0_9 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  tag_0_10 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  tag_0_11 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  tag_0_12 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  tag_0_13 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  tag_0_14 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  tag_0_15 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  tag_0_16 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  tag_0_17 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  tag_0_18 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  tag_0_19 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  tag_0_20 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  tag_0_21 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  tag_0_22 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  tag_0_23 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  tag_0_24 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  tag_0_25 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  tag_0_26 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  tag_0_27 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  tag_0_28 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  tag_0_29 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  tag_0_30 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  tag_0_31 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  tag_0_32 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  tag_0_33 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  tag_0_34 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  tag_0_35 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  tag_0_36 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  tag_0_37 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  tag_0_38 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  tag_0_39 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  tag_0_40 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  tag_0_41 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  tag_0_42 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  tag_0_43 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  tag_0_44 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  tag_0_45 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  tag_0_46 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  tag_0_47 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  tag_0_48 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  tag_0_49 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  tag_0_50 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  tag_0_51 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  tag_0_52 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  tag_0_53 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  tag_0_54 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  tag_0_55 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  tag_0_56 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  tag_0_57 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  tag_0_58 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  tag_0_59 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  tag_0_60 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  tag_0_61 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  tag_0_62 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  tag_0_63 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  tag_0_64 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  tag_0_65 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  tag_0_66 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  tag_0_67 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  tag_0_68 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  tag_0_69 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  tag_0_70 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  tag_0_71 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  tag_0_72 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  tag_0_73 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  tag_0_74 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  tag_0_75 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  tag_0_76 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  tag_0_77 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  tag_0_78 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  tag_0_79 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  tag_0_80 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  tag_0_81 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  tag_0_82 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  tag_0_83 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  tag_0_84 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  tag_0_85 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  tag_0_86 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  tag_0_87 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  tag_0_88 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  tag_0_89 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  tag_0_90 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  tag_0_91 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  tag_0_92 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  tag_0_93 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  tag_0_94 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  tag_0_95 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  tag_0_96 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  tag_0_97 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  tag_0_98 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  tag_0_99 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  tag_0_100 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  tag_0_101 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  tag_0_102 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  tag_0_103 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  tag_0_104 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  tag_0_105 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  tag_0_106 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  tag_0_107 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  tag_0_108 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  tag_0_109 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  tag_0_110 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  tag_0_111 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  tag_0_112 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  tag_0_113 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  tag_0_114 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  tag_0_115 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  tag_0_116 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  tag_0_117 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  tag_0_118 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  tag_0_119 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  tag_0_120 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  tag_0_121 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  tag_0_122 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  tag_0_123 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  tag_0_124 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  tag_0_125 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  tag_0_126 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  tag_0_127 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  tag_1_0 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  tag_1_1 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  tag_1_2 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  tag_1_3 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  tag_1_4 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  tag_1_5 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  tag_1_6 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  tag_1_7 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  tag_1_8 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  tag_1_9 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  tag_1_10 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  tag_1_11 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  tag_1_12 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  tag_1_13 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  tag_1_14 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  tag_1_15 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  tag_1_16 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  tag_1_17 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  tag_1_18 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  tag_1_19 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  tag_1_20 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  tag_1_21 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  tag_1_22 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  tag_1_23 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  tag_1_24 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  tag_1_25 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  tag_1_26 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  tag_1_27 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  tag_1_28 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  tag_1_29 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  tag_1_30 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  tag_1_31 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  tag_1_32 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  tag_1_33 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  tag_1_34 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  tag_1_35 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  tag_1_36 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  tag_1_37 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  tag_1_38 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  tag_1_39 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  tag_1_40 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  tag_1_41 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  tag_1_42 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  tag_1_43 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  tag_1_44 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  tag_1_45 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  tag_1_46 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  tag_1_47 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  tag_1_48 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  tag_1_49 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  tag_1_50 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  tag_1_51 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  tag_1_52 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  tag_1_53 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  tag_1_54 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  tag_1_55 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  tag_1_56 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  tag_1_57 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  tag_1_58 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  tag_1_59 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  tag_1_60 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  tag_1_61 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  tag_1_62 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  tag_1_63 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  tag_1_64 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  tag_1_65 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  tag_1_66 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  tag_1_67 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  tag_1_68 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  tag_1_69 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  tag_1_70 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  tag_1_71 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  tag_1_72 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  tag_1_73 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  tag_1_74 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  tag_1_75 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  tag_1_76 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  tag_1_77 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  tag_1_78 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  tag_1_79 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  tag_1_80 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  tag_1_81 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  tag_1_82 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  tag_1_83 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  tag_1_84 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  tag_1_85 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  tag_1_86 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  tag_1_87 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  tag_1_88 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  tag_1_89 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  tag_1_90 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  tag_1_91 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  tag_1_92 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  tag_1_93 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  tag_1_94 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  tag_1_95 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  tag_1_96 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  tag_1_97 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  tag_1_98 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  tag_1_99 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  tag_1_100 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  tag_1_101 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  tag_1_102 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  tag_1_103 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  tag_1_104 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  tag_1_105 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  tag_1_106 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  tag_1_107 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  tag_1_108 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  tag_1_109 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  tag_1_110 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  tag_1_111 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  tag_1_112 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  tag_1_113 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  tag_1_114 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  tag_1_115 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  tag_1_116 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  tag_1_117 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  tag_1_118 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  tag_1_119 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  tag_1_120 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  tag_1_121 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  tag_1_122 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  tag_1_123 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  tag_1_124 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  tag_1_125 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  tag_1_126 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  tag_1_127 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  valid_0_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid_0_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  valid_0_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  valid_0_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  valid_0_4 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  valid_0_5 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  valid_0_6 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  valid_0_7 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  valid_0_8 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  valid_0_9 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  valid_0_10 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  valid_0_11 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  valid_0_12 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  valid_0_13 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  valid_0_14 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  valid_0_15 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  valid_0_16 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  valid_0_17 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  valid_0_18 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  valid_0_19 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  valid_0_20 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  valid_0_21 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  valid_0_22 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  valid_0_23 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  valid_0_24 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  valid_0_25 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  valid_0_26 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  valid_0_27 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  valid_0_28 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  valid_0_29 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  valid_0_30 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  valid_0_31 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  valid_0_32 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  valid_0_33 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  valid_0_34 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  valid_0_35 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  valid_0_36 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  valid_0_37 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  valid_0_38 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  valid_0_39 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  valid_0_40 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  valid_0_41 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  valid_0_42 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  valid_0_43 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  valid_0_44 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  valid_0_45 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  valid_0_46 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  valid_0_47 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  valid_0_48 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  valid_0_49 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  valid_0_50 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  valid_0_51 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  valid_0_52 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  valid_0_53 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  valid_0_54 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  valid_0_55 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  valid_0_56 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  valid_0_57 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  valid_0_58 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  valid_0_59 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  valid_0_60 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  valid_0_61 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  valid_0_62 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  valid_0_63 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  valid_0_64 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  valid_0_65 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  valid_0_66 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  valid_0_67 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  valid_0_68 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  valid_0_69 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  valid_0_70 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  valid_0_71 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  valid_0_72 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  valid_0_73 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  valid_0_74 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  valid_0_75 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  valid_0_76 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  valid_0_77 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  valid_0_78 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  valid_0_79 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  valid_0_80 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  valid_0_81 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  valid_0_82 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  valid_0_83 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  valid_0_84 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  valid_0_85 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  valid_0_86 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  valid_0_87 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  valid_0_88 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  valid_0_89 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  valid_0_90 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  valid_0_91 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  valid_0_92 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  valid_0_93 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  valid_0_94 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  valid_0_95 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  valid_0_96 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  valid_0_97 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  valid_0_98 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  valid_0_99 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  valid_0_100 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  valid_0_101 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  valid_0_102 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  valid_0_103 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  valid_0_104 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  valid_0_105 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  valid_0_106 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  valid_0_107 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  valid_0_108 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  valid_0_109 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  valid_0_110 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  valid_0_111 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  valid_0_112 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  valid_0_113 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  valid_0_114 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  valid_0_115 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  valid_0_116 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  valid_0_117 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  valid_0_118 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  valid_0_119 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  valid_0_120 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  valid_0_121 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  valid_0_122 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  valid_0_123 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  valid_0_124 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  valid_0_125 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  valid_0_126 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  valid_0_127 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  valid_1_0 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  valid_1_1 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  valid_1_2 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  valid_1_3 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  valid_1_4 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  valid_1_5 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  valid_1_6 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  valid_1_7 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  valid_1_8 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  valid_1_9 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  valid_1_10 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  valid_1_11 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  valid_1_12 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  valid_1_13 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  valid_1_14 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  valid_1_15 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  valid_1_16 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  valid_1_17 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  valid_1_18 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  valid_1_19 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  valid_1_20 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  valid_1_21 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  valid_1_22 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  valid_1_23 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  valid_1_24 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  valid_1_25 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  valid_1_26 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  valid_1_27 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  valid_1_28 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  valid_1_29 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  valid_1_30 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  valid_1_31 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  valid_1_32 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  valid_1_33 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  valid_1_34 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  valid_1_35 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  valid_1_36 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  valid_1_37 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  valid_1_38 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  valid_1_39 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  valid_1_40 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  valid_1_41 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  valid_1_42 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  valid_1_43 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  valid_1_44 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  valid_1_45 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  valid_1_46 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  valid_1_47 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  valid_1_48 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  valid_1_49 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  valid_1_50 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  valid_1_51 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  valid_1_52 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  valid_1_53 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  valid_1_54 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  valid_1_55 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  valid_1_56 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  valid_1_57 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  valid_1_58 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  valid_1_59 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  valid_1_60 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  valid_1_61 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  valid_1_62 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  valid_1_63 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  valid_1_64 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  valid_1_65 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  valid_1_66 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  valid_1_67 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  valid_1_68 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  valid_1_69 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  valid_1_70 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  valid_1_71 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  valid_1_72 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  valid_1_73 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  valid_1_74 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  valid_1_75 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  valid_1_76 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  valid_1_77 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  valid_1_78 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  valid_1_79 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  valid_1_80 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  valid_1_81 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  valid_1_82 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  valid_1_83 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  valid_1_84 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  valid_1_85 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  valid_1_86 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  valid_1_87 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  valid_1_88 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  valid_1_89 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  valid_1_90 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  valid_1_91 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  valid_1_92 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  valid_1_93 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  valid_1_94 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  valid_1_95 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  valid_1_96 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  valid_1_97 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  valid_1_98 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  valid_1_99 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  valid_1_100 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  valid_1_101 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  valid_1_102 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  valid_1_103 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  valid_1_104 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  valid_1_105 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  valid_1_106 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  valid_1_107 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  valid_1_108 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  valid_1_109 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  valid_1_110 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  valid_1_111 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  valid_1_112 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  valid_1_113 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  valid_1_114 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  valid_1_115 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  valid_1_116 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  valid_1_117 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  valid_1_118 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  valid_1_119 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  valid_1_120 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  valid_1_121 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  valid_1_122 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  valid_1_123 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  valid_1_124 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  valid_1_125 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  valid_1_126 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  valid_1_127 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  way0_hit = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  way1_hit = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  unuse_way = _RAND_770[1:0];
  _RAND_771 = {2{`RANDOM}};
  receive_data = _RAND_771[63:0];
  _RAND_772 = {1{`RANDOM}};
  quene = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  state = _RAND_773[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module D_CACHE(
  input         clock,
  input         reset,
  input  [63:0] io_pc_now,
  input  [31:0] io_from_lsu_araddr,
  input         io_from_lsu_arvalid,
  input         io_from_lsu_rready,
  input  [31:0] io_from_lsu_awaddr,
  input         io_from_lsu_awvalid,
  input  [63:0] io_from_lsu_wdata,
  input  [7:0]  io_from_lsu_wstrb,
  input         io_from_lsu_wvalid,
  input         io_from_lsu_bready,
  output        io_to_lsu_arready,
  output [63:0] io_to_lsu_rdata,
  output        io_to_lsu_rvalid,
  output        io_to_lsu_awready,
  output        io_to_lsu_wready,
  output        io_to_lsu_bvalid,
  output [31:0] io_to_axi_araddr,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  output [31:0] io_to_axi_awaddr,
  output        io_to_axi_awvalid,
  output [63:0] io_to_axi_wdata,
  output [7:0]  io_to_axi_wstrb,
  output        io_to_axi_wvalid,
  output        io_to_axi_bready,
  input         io_from_axi_arready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rvalid,
  input         io_from_axi_awready,
  input         io_from_axi_wready,
  input         io_from_axi_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [63:0] _RAND_256;
  reg [63:0] _RAND_257;
  reg [63:0] _RAND_258;
  reg [63:0] _RAND_259;
  reg [63:0] _RAND_260;
  reg [63:0] _RAND_261;
  reg [63:0] _RAND_262;
  reg [63:0] _RAND_263;
  reg [63:0] _RAND_264;
  reg [63:0] _RAND_265;
  reg [63:0] _RAND_266;
  reg [63:0] _RAND_267;
  reg [63:0] _RAND_268;
  reg [63:0] _RAND_269;
  reg [63:0] _RAND_270;
  reg [63:0] _RAND_271;
  reg [63:0] _RAND_272;
  reg [63:0] _RAND_273;
  reg [63:0] _RAND_274;
  reg [63:0] _RAND_275;
  reg [63:0] _RAND_276;
  reg [63:0] _RAND_277;
  reg [63:0] _RAND_278;
  reg [63:0] _RAND_279;
  reg [63:0] _RAND_280;
  reg [63:0] _RAND_281;
  reg [63:0] _RAND_282;
  reg [63:0] _RAND_283;
  reg [63:0] _RAND_284;
  reg [63:0] _RAND_285;
  reg [63:0] _RAND_286;
  reg [63:0] _RAND_287;
  reg [63:0] _RAND_288;
  reg [63:0] _RAND_289;
  reg [63:0] _RAND_290;
  reg [63:0] _RAND_291;
  reg [63:0] _RAND_292;
  reg [63:0] _RAND_293;
  reg [63:0] _RAND_294;
  reg [63:0] _RAND_295;
  reg [63:0] _RAND_296;
  reg [63:0] _RAND_297;
  reg [63:0] _RAND_298;
  reg [63:0] _RAND_299;
  reg [63:0] _RAND_300;
  reg [63:0] _RAND_301;
  reg [63:0] _RAND_302;
  reg [63:0] _RAND_303;
  reg [63:0] _RAND_304;
  reg [63:0] _RAND_305;
  reg [63:0] _RAND_306;
  reg [63:0] _RAND_307;
  reg [63:0] _RAND_308;
  reg [63:0] _RAND_309;
  reg [63:0] _RAND_310;
  reg [63:0] _RAND_311;
  reg [63:0] _RAND_312;
  reg [63:0] _RAND_313;
  reg [63:0] _RAND_314;
  reg [63:0] _RAND_315;
  reg [63:0] _RAND_316;
  reg [63:0] _RAND_317;
  reg [63:0] _RAND_318;
  reg [63:0] _RAND_319;
  reg [63:0] _RAND_320;
  reg [63:0] _RAND_321;
  reg [63:0] _RAND_322;
  reg [63:0] _RAND_323;
  reg [63:0] _RAND_324;
  reg [63:0] _RAND_325;
  reg [63:0] _RAND_326;
  reg [63:0] _RAND_327;
  reg [63:0] _RAND_328;
  reg [63:0] _RAND_329;
  reg [63:0] _RAND_330;
  reg [63:0] _RAND_331;
  reg [63:0] _RAND_332;
  reg [63:0] _RAND_333;
  reg [63:0] _RAND_334;
  reg [63:0] _RAND_335;
  reg [63:0] _RAND_336;
  reg [63:0] _RAND_337;
  reg [63:0] _RAND_338;
  reg [63:0] _RAND_339;
  reg [63:0] _RAND_340;
  reg [63:0] _RAND_341;
  reg [63:0] _RAND_342;
  reg [63:0] _RAND_343;
  reg [63:0] _RAND_344;
  reg [63:0] _RAND_345;
  reg [63:0] _RAND_346;
  reg [63:0] _RAND_347;
  reg [63:0] _RAND_348;
  reg [63:0] _RAND_349;
  reg [63:0] _RAND_350;
  reg [63:0] _RAND_351;
  reg [63:0] _RAND_352;
  reg [63:0] _RAND_353;
  reg [63:0] _RAND_354;
  reg [63:0] _RAND_355;
  reg [63:0] _RAND_356;
  reg [63:0] _RAND_357;
  reg [63:0] _RAND_358;
  reg [63:0] _RAND_359;
  reg [63:0] _RAND_360;
  reg [63:0] _RAND_361;
  reg [63:0] _RAND_362;
  reg [63:0] _RAND_363;
  reg [63:0] _RAND_364;
  reg [63:0] _RAND_365;
  reg [63:0] _RAND_366;
  reg [63:0] _RAND_367;
  reg [63:0] _RAND_368;
  reg [63:0] _RAND_369;
  reg [63:0] _RAND_370;
  reg [63:0] _RAND_371;
  reg [63:0] _RAND_372;
  reg [63:0] _RAND_373;
  reg [63:0] _RAND_374;
  reg [63:0] _RAND_375;
  reg [63:0] _RAND_376;
  reg [63:0] _RAND_377;
  reg [63:0] _RAND_378;
  reg [63:0] _RAND_379;
  reg [63:0] _RAND_380;
  reg [63:0] _RAND_381;
  reg [63:0] _RAND_382;
  reg [63:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [63:0] _RAND_512;
  reg [63:0] _RAND_513;
  reg [63:0] _RAND_514;
  reg [63:0] _RAND_515;
  reg [63:0] _RAND_516;
  reg [63:0] _RAND_517;
  reg [63:0] _RAND_518;
  reg [63:0] _RAND_519;
  reg [63:0] _RAND_520;
  reg [63:0] _RAND_521;
  reg [63:0] _RAND_522;
  reg [63:0] _RAND_523;
  reg [63:0] _RAND_524;
  reg [63:0] _RAND_525;
  reg [63:0] _RAND_526;
  reg [63:0] _RAND_527;
  reg [63:0] _RAND_528;
  reg [63:0] _RAND_529;
  reg [63:0] _RAND_530;
  reg [63:0] _RAND_531;
  reg [63:0] _RAND_532;
  reg [63:0] _RAND_533;
  reg [63:0] _RAND_534;
  reg [63:0] _RAND_535;
  reg [63:0] _RAND_536;
  reg [63:0] _RAND_537;
  reg [63:0] _RAND_538;
  reg [63:0] _RAND_539;
  reg [63:0] _RAND_540;
  reg [63:0] _RAND_541;
  reg [63:0] _RAND_542;
  reg [63:0] _RAND_543;
  reg [63:0] _RAND_544;
  reg [63:0] _RAND_545;
  reg [63:0] _RAND_546;
  reg [63:0] _RAND_547;
  reg [63:0] _RAND_548;
  reg [63:0] _RAND_549;
  reg [63:0] _RAND_550;
  reg [63:0] _RAND_551;
  reg [63:0] _RAND_552;
  reg [63:0] _RAND_553;
  reg [63:0] _RAND_554;
  reg [63:0] _RAND_555;
  reg [63:0] _RAND_556;
  reg [63:0] _RAND_557;
  reg [63:0] _RAND_558;
  reg [63:0] _RAND_559;
  reg [63:0] _RAND_560;
  reg [63:0] _RAND_561;
  reg [63:0] _RAND_562;
  reg [63:0] _RAND_563;
  reg [63:0] _RAND_564;
  reg [63:0] _RAND_565;
  reg [63:0] _RAND_566;
  reg [63:0] _RAND_567;
  reg [63:0] _RAND_568;
  reg [63:0] _RAND_569;
  reg [63:0] _RAND_570;
  reg [63:0] _RAND_571;
  reg [63:0] _RAND_572;
  reg [63:0] _RAND_573;
  reg [63:0] _RAND_574;
  reg [63:0] _RAND_575;
  reg [63:0] _RAND_576;
  reg [63:0] _RAND_577;
  reg [63:0] _RAND_578;
  reg [63:0] _RAND_579;
  reg [63:0] _RAND_580;
  reg [63:0] _RAND_581;
  reg [63:0] _RAND_582;
  reg [63:0] _RAND_583;
  reg [63:0] _RAND_584;
  reg [63:0] _RAND_585;
  reg [63:0] _RAND_586;
  reg [63:0] _RAND_587;
  reg [63:0] _RAND_588;
  reg [63:0] _RAND_589;
  reg [63:0] _RAND_590;
  reg [63:0] _RAND_591;
  reg [63:0] _RAND_592;
  reg [63:0] _RAND_593;
  reg [63:0] _RAND_594;
  reg [63:0] _RAND_595;
  reg [63:0] _RAND_596;
  reg [63:0] _RAND_597;
  reg [63:0] _RAND_598;
  reg [63:0] _RAND_599;
  reg [63:0] _RAND_600;
  reg [63:0] _RAND_601;
  reg [63:0] _RAND_602;
  reg [63:0] _RAND_603;
  reg [63:0] _RAND_604;
  reg [63:0] _RAND_605;
  reg [63:0] _RAND_606;
  reg [63:0] _RAND_607;
  reg [63:0] _RAND_608;
  reg [63:0] _RAND_609;
  reg [63:0] _RAND_610;
  reg [63:0] _RAND_611;
  reg [63:0] _RAND_612;
  reg [63:0] _RAND_613;
  reg [63:0] _RAND_614;
  reg [63:0] _RAND_615;
  reg [63:0] _RAND_616;
  reg [63:0] _RAND_617;
  reg [63:0] _RAND_618;
  reg [63:0] _RAND_619;
  reg [63:0] _RAND_620;
  reg [63:0] _RAND_621;
  reg [63:0] _RAND_622;
  reg [63:0] _RAND_623;
  reg [63:0] _RAND_624;
  reg [63:0] _RAND_625;
  reg [63:0] _RAND_626;
  reg [63:0] _RAND_627;
  reg [63:0] _RAND_628;
  reg [63:0] _RAND_629;
  reg [63:0] _RAND_630;
  reg [63:0] _RAND_631;
  reg [63:0] _RAND_632;
  reg [63:0] _RAND_633;
  reg [63:0] _RAND_634;
  reg [63:0] _RAND_635;
  reg [63:0] _RAND_636;
  reg [63:0] _RAND_637;
  reg [63:0] _RAND_638;
  reg [63:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [63:0] _RAND_768;
  reg [63:0] _RAND_769;
  reg [63:0] _RAND_770;
  reg [63:0] _RAND_771;
  reg [63:0] _RAND_772;
  reg [63:0] _RAND_773;
  reg [63:0] _RAND_774;
  reg [63:0] _RAND_775;
  reg [63:0] _RAND_776;
  reg [63:0] _RAND_777;
  reg [63:0] _RAND_778;
  reg [63:0] _RAND_779;
  reg [63:0] _RAND_780;
  reg [63:0] _RAND_781;
  reg [63:0] _RAND_782;
  reg [63:0] _RAND_783;
  reg [63:0] _RAND_784;
  reg [63:0] _RAND_785;
  reg [63:0] _RAND_786;
  reg [63:0] _RAND_787;
  reg [63:0] _RAND_788;
  reg [63:0] _RAND_789;
  reg [63:0] _RAND_790;
  reg [63:0] _RAND_791;
  reg [63:0] _RAND_792;
  reg [63:0] _RAND_793;
  reg [63:0] _RAND_794;
  reg [63:0] _RAND_795;
  reg [63:0] _RAND_796;
  reg [63:0] _RAND_797;
  reg [63:0] _RAND_798;
  reg [63:0] _RAND_799;
  reg [63:0] _RAND_800;
  reg [63:0] _RAND_801;
  reg [63:0] _RAND_802;
  reg [63:0] _RAND_803;
  reg [63:0] _RAND_804;
  reg [63:0] _RAND_805;
  reg [63:0] _RAND_806;
  reg [63:0] _RAND_807;
  reg [63:0] _RAND_808;
  reg [63:0] _RAND_809;
  reg [63:0] _RAND_810;
  reg [63:0] _RAND_811;
  reg [63:0] _RAND_812;
  reg [63:0] _RAND_813;
  reg [63:0] _RAND_814;
  reg [63:0] _RAND_815;
  reg [63:0] _RAND_816;
  reg [63:0] _RAND_817;
  reg [63:0] _RAND_818;
  reg [63:0] _RAND_819;
  reg [63:0] _RAND_820;
  reg [63:0] _RAND_821;
  reg [63:0] _RAND_822;
  reg [63:0] _RAND_823;
  reg [63:0] _RAND_824;
  reg [63:0] _RAND_825;
  reg [63:0] _RAND_826;
  reg [63:0] _RAND_827;
  reg [63:0] _RAND_828;
  reg [63:0] _RAND_829;
  reg [63:0] _RAND_830;
  reg [63:0] _RAND_831;
  reg [63:0] _RAND_832;
  reg [63:0] _RAND_833;
  reg [63:0] _RAND_834;
  reg [63:0] _RAND_835;
  reg [63:0] _RAND_836;
  reg [63:0] _RAND_837;
  reg [63:0] _RAND_838;
  reg [63:0] _RAND_839;
  reg [63:0] _RAND_840;
  reg [63:0] _RAND_841;
  reg [63:0] _RAND_842;
  reg [63:0] _RAND_843;
  reg [63:0] _RAND_844;
  reg [63:0] _RAND_845;
  reg [63:0] _RAND_846;
  reg [63:0] _RAND_847;
  reg [63:0] _RAND_848;
  reg [63:0] _RAND_849;
  reg [63:0] _RAND_850;
  reg [63:0] _RAND_851;
  reg [63:0] _RAND_852;
  reg [63:0] _RAND_853;
  reg [63:0] _RAND_854;
  reg [63:0] _RAND_855;
  reg [63:0] _RAND_856;
  reg [63:0] _RAND_857;
  reg [63:0] _RAND_858;
  reg [63:0] _RAND_859;
  reg [63:0] _RAND_860;
  reg [63:0] _RAND_861;
  reg [63:0] _RAND_862;
  reg [63:0] _RAND_863;
  reg [63:0] _RAND_864;
  reg [63:0] _RAND_865;
  reg [63:0] _RAND_866;
  reg [63:0] _RAND_867;
  reg [63:0] _RAND_868;
  reg [63:0] _RAND_869;
  reg [63:0] _RAND_870;
  reg [63:0] _RAND_871;
  reg [63:0] _RAND_872;
  reg [63:0] _RAND_873;
  reg [63:0] _RAND_874;
  reg [63:0] _RAND_875;
  reg [63:0] _RAND_876;
  reg [63:0] _RAND_877;
  reg [63:0] _RAND_878;
  reg [63:0] _RAND_879;
  reg [63:0] _RAND_880;
  reg [63:0] _RAND_881;
  reg [63:0] _RAND_882;
  reg [63:0] _RAND_883;
  reg [63:0] _RAND_884;
  reg [63:0] _RAND_885;
  reg [63:0] _RAND_886;
  reg [63:0] _RAND_887;
  reg [63:0] _RAND_888;
  reg [63:0] _RAND_889;
  reg [63:0] _RAND_890;
  reg [63:0] _RAND_891;
  reg [63:0] _RAND_892;
  reg [63:0] _RAND_893;
  reg [63:0] _RAND_894;
  reg [63:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [63:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [63:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = ~reset; // @[d_cache.scala 16:11]
  reg [63:0] ram_0_0; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_1; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_2; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_3; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_4; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_5; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_6; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_7; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_8; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_9; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_10; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_11; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_12; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_13; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_14; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_15; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_16; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_17; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_18; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_19; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_20; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_21; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_22; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_23; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_24; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_25; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_26; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_27; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_28; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_29; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_30; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_31; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_32; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_33; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_34; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_35; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_36; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_37; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_38; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_39; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_40; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_41; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_42; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_43; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_44; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_45; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_46; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_47; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_48; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_49; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_50; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_51; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_52; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_53; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_54; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_55; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_56; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_57; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_58; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_59; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_60; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_61; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_62; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_63; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_64; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_65; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_66; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_67; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_68; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_69; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_70; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_71; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_72; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_73; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_74; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_75; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_76; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_77; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_78; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_79; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_80; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_81; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_82; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_83; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_84; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_85; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_86; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_87; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_88; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_89; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_90; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_91; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_92; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_93; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_94; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_95; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_96; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_97; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_98; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_99; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_100; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_101; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_102; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_103; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_104; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_105; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_106; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_107; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_108; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_109; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_110; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_111; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_112; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_113; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_114; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_115; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_116; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_117; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_118; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_119; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_120; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_121; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_122; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_123; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_124; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_125; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_126; // @[d_cache.scala 19:24]
  reg [63:0] ram_0_127; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_0; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_1; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_2; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_3; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_4; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_5; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_6; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_7; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_8; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_9; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_10; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_11; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_12; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_13; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_14; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_15; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_16; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_17; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_18; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_19; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_20; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_21; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_22; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_23; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_24; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_25; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_26; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_27; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_28; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_29; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_30; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_31; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_32; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_33; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_34; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_35; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_36; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_37; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_38; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_39; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_40; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_41; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_42; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_43; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_44; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_45; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_46; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_47; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_48; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_49; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_50; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_51; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_52; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_53; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_54; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_55; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_56; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_57; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_58; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_59; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_60; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_61; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_62; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_63; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_64; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_65; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_66; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_67; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_68; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_69; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_70; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_71; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_72; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_73; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_74; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_75; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_76; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_77; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_78; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_79; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_80; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_81; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_82; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_83; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_84; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_85; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_86; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_87; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_88; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_89; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_90; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_91; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_92; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_93; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_94; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_95; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_96; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_97; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_98; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_99; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_100; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_101; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_102; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_103; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_104; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_105; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_106; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_107; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_108; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_109; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_110; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_111; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_112; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_113; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_114; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_115; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_116; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_117; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_118; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_119; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_120; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_121; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_122; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_123; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_124; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_125; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_126; // @[d_cache.scala 20:24]
  reg [63:0] ram_1_127; // @[d_cache.scala 20:24]
  reg [63:0] record_wdata1_0; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_1; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_2; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_3; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_4; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_5; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_6; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_7; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_8; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_9; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_10; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_11; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_12; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_13; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_14; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_15; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_16; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_17; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_18; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_19; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_20; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_21; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_22; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_23; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_24; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_25; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_26; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_27; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_28; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_29; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_30; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_31; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_32; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_33; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_34; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_35; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_36; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_37; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_38; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_39; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_40; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_41; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_42; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_43; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_44; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_45; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_46; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_47; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_48; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_49; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_50; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_51; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_52; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_53; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_54; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_55; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_56; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_57; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_58; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_59; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_60; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_61; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_62; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_63; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_64; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_65; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_66; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_67; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_68; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_69; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_70; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_71; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_72; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_73; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_74; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_75; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_76; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_77; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_78; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_79; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_80; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_81; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_82; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_83; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_84; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_85; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_86; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_87; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_88; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_89; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_90; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_91; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_92; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_93; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_94; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_95; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_96; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_97; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_98; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_99; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_100; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_101; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_102; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_103; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_104; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_105; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_106; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_107; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_108; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_109; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_110; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_111; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_112; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_113; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_114; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_115; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_116; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_117; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_118; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_119; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_120; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_121; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_122; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_123; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_124; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_125; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_126; // @[d_cache.scala 21:32]
  reg [63:0] record_wdata1_127; // @[d_cache.scala 21:32]
  reg [7:0] record_wstrb1_0; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_1; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_2; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_3; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_4; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_5; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_6; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_7; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_8; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_9; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_10; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_11; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_12; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_13; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_14; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_15; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_16; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_17; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_18; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_19; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_20; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_21; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_22; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_23; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_24; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_25; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_26; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_27; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_28; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_29; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_30; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_31; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_32; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_33; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_34; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_35; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_36; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_37; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_38; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_39; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_40; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_41; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_42; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_43; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_44; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_45; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_46; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_47; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_48; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_49; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_50; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_51; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_52; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_53; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_54; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_55; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_56; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_57; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_58; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_59; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_60; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_61; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_62; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_63; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_64; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_65; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_66; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_67; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_68; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_69; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_70; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_71; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_72; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_73; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_74; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_75; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_76; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_77; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_78; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_79; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_80; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_81; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_82; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_83; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_84; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_85; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_86; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_87; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_88; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_89; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_90; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_91; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_92; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_93; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_94; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_95; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_96; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_97; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_98; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_99; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_100; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_101; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_102; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_103; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_104; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_105; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_106; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_107; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_108; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_109; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_110; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_111; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_112; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_113; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_114; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_115; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_116; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_117; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_118; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_119; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_120; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_121; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_122; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_123; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_124; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_125; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_126; // @[d_cache.scala 22:32]
  reg [7:0] record_wstrb1_127; // @[d_cache.scala 22:32]
  reg [63:0] record_pc_0; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_1; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_2; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_3; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_4; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_5; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_6; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_7; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_8; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_9; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_10; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_11; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_12; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_13; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_14; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_15; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_16; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_17; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_18; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_19; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_20; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_21; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_22; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_23; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_24; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_25; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_26; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_27; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_28; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_29; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_30; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_31; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_32; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_33; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_34; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_35; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_36; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_37; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_38; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_39; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_40; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_41; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_42; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_43; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_44; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_45; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_46; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_47; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_48; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_49; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_50; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_51; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_52; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_53; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_54; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_55; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_56; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_57; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_58; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_59; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_60; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_61; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_62; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_63; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_64; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_65; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_66; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_67; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_68; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_69; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_70; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_71; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_72; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_73; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_74; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_75; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_76; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_77; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_78; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_79; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_80; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_81; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_82; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_83; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_84; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_85; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_86; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_87; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_88; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_89; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_90; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_91; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_92; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_93; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_94; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_95; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_96; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_97; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_98; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_99; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_100; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_101; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_102; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_103; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_104; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_105; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_106; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_107; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_108; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_109; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_110; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_111; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_112; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_113; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_114; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_115; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_116; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_117; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_118; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_119; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_120; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_121; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_122; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_123; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_124; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_125; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_126; // @[d_cache.scala 23:28]
  reg [63:0] record_pc_127; // @[d_cache.scala 23:28]
  reg [31:0] record_addr_0; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_1; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_2; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_3; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_4; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_5; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_6; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_7; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_8; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_9; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_10; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_11; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_12; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_13; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_14; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_15; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_16; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_17; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_18; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_19; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_20; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_21; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_22; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_23; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_24; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_25; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_26; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_27; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_28; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_29; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_30; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_31; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_32; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_33; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_34; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_35; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_36; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_37; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_38; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_39; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_40; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_41; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_42; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_43; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_44; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_45; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_46; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_47; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_48; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_49; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_50; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_51; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_52; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_53; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_54; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_55; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_56; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_57; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_58; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_59; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_60; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_61; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_62; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_63; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_64; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_65; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_66; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_67; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_68; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_69; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_70; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_71; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_72; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_73; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_74; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_75; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_76; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_77; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_78; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_79; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_80; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_81; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_82; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_83; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_84; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_85; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_86; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_87; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_88; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_89; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_90; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_91; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_92; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_93; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_94; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_95; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_96; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_97; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_98; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_99; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_100; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_101; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_102; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_103; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_104; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_105; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_106; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_107; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_108; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_109; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_110; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_111; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_112; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_113; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_114; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_115; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_116; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_117; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_118; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_119; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_120; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_121; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_122; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_123; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_124; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_125; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_126; // @[d_cache.scala 24:30]
  reg [31:0] record_addr_127; // @[d_cache.scala 24:30]
  reg [63:0] record_olddata_0; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_1; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_2; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_3; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_4; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_5; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_6; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_7; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_8; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_9; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_10; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_11; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_12; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_13; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_14; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_15; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_16; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_17; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_18; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_19; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_20; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_21; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_22; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_23; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_24; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_25; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_26; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_27; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_28; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_29; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_30; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_31; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_32; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_33; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_34; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_35; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_36; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_37; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_38; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_39; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_40; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_41; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_42; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_43; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_44; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_45; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_46; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_47; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_48; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_49; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_50; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_51; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_52; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_53; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_54; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_55; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_56; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_57; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_58; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_59; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_60; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_61; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_62; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_63; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_64; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_65; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_66; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_67; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_68; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_69; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_70; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_71; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_72; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_73; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_74; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_75; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_76; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_77; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_78; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_79; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_80; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_81; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_82; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_83; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_84; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_85; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_86; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_87; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_88; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_89; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_90; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_91; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_92; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_93; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_94; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_95; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_96; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_97; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_98; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_99; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_100; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_101; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_102; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_103; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_104; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_105; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_106; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_107; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_108; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_109; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_110; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_111; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_112; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_113; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_114; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_115; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_116; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_117; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_118; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_119; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_120; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_121; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_122; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_123; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_124; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_125; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_126; // @[d_cache.scala 25:33]
  reg [63:0] record_olddata_127; // @[d_cache.scala 25:33]
  reg [31:0] tag_0_0; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_1; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_2; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_3; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_4; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_5; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_6; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_7; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_8; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_9; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_10; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_11; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_12; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_13; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_14; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_15; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_16; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_17; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_18; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_19; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_20; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_21; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_22; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_23; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_24; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_25; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_26; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_27; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_28; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_29; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_30; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_31; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_32; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_33; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_34; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_35; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_36; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_37; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_38; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_39; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_40; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_41; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_42; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_43; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_44; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_45; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_46; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_47; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_48; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_49; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_50; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_51; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_52; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_53; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_54; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_55; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_56; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_57; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_58; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_59; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_60; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_61; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_62; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_63; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_64; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_65; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_66; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_67; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_68; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_69; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_70; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_71; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_72; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_73; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_74; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_75; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_76; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_77; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_78; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_79; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_80; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_81; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_82; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_83; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_84; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_85; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_86; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_87; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_88; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_89; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_90; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_91; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_92; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_93; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_94; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_95; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_96; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_97; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_98; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_99; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_100; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_101; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_102; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_103; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_104; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_105; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_106; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_107; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_108; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_109; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_110; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_111; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_112; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_113; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_114; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_115; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_116; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_117; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_118; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_119; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_120; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_121; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_122; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_123; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_124; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_125; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_126; // @[d_cache.scala 28:24]
  reg [31:0] tag_0_127; // @[d_cache.scala 28:24]
  reg [31:0] tag_1_0; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_1; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_2; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_3; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_4; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_5; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_6; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_7; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_8; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_9; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_10; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_11; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_12; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_13; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_14; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_15; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_16; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_17; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_18; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_19; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_20; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_21; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_22; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_23; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_24; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_25; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_26; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_27; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_28; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_29; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_30; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_31; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_32; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_33; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_34; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_35; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_36; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_37; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_38; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_39; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_40; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_41; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_42; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_43; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_44; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_45; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_46; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_47; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_48; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_49; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_50; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_51; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_52; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_53; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_54; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_55; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_56; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_57; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_58; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_59; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_60; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_61; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_62; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_63; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_64; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_65; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_66; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_67; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_68; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_69; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_70; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_71; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_72; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_73; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_74; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_75; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_76; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_77; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_78; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_79; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_80; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_81; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_82; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_83; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_84; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_85; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_86; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_87; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_88; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_89; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_90; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_91; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_92; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_93; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_94; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_95; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_96; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_97; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_98; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_99; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_100; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_101; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_102; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_103; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_104; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_105; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_106; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_107; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_108; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_109; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_110; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_111; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_112; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_113; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_114; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_115; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_116; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_117; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_118; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_119; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_120; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_121; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_122; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_123; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_124; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_125; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_126; // @[d_cache.scala 29:24]
  reg [31:0] tag_1_127; // @[d_cache.scala 29:24]
  reg  valid_0_0; // @[d_cache.scala 30:26]
  reg  valid_0_1; // @[d_cache.scala 30:26]
  reg  valid_0_2; // @[d_cache.scala 30:26]
  reg  valid_0_3; // @[d_cache.scala 30:26]
  reg  valid_0_4; // @[d_cache.scala 30:26]
  reg  valid_0_5; // @[d_cache.scala 30:26]
  reg  valid_0_6; // @[d_cache.scala 30:26]
  reg  valid_0_7; // @[d_cache.scala 30:26]
  reg  valid_0_8; // @[d_cache.scala 30:26]
  reg  valid_0_9; // @[d_cache.scala 30:26]
  reg  valid_0_10; // @[d_cache.scala 30:26]
  reg  valid_0_11; // @[d_cache.scala 30:26]
  reg  valid_0_12; // @[d_cache.scala 30:26]
  reg  valid_0_13; // @[d_cache.scala 30:26]
  reg  valid_0_14; // @[d_cache.scala 30:26]
  reg  valid_0_15; // @[d_cache.scala 30:26]
  reg  valid_0_16; // @[d_cache.scala 30:26]
  reg  valid_0_17; // @[d_cache.scala 30:26]
  reg  valid_0_18; // @[d_cache.scala 30:26]
  reg  valid_0_19; // @[d_cache.scala 30:26]
  reg  valid_0_20; // @[d_cache.scala 30:26]
  reg  valid_0_21; // @[d_cache.scala 30:26]
  reg  valid_0_22; // @[d_cache.scala 30:26]
  reg  valid_0_23; // @[d_cache.scala 30:26]
  reg  valid_0_24; // @[d_cache.scala 30:26]
  reg  valid_0_25; // @[d_cache.scala 30:26]
  reg  valid_0_26; // @[d_cache.scala 30:26]
  reg  valid_0_27; // @[d_cache.scala 30:26]
  reg  valid_0_28; // @[d_cache.scala 30:26]
  reg  valid_0_29; // @[d_cache.scala 30:26]
  reg  valid_0_30; // @[d_cache.scala 30:26]
  reg  valid_0_31; // @[d_cache.scala 30:26]
  reg  valid_0_32; // @[d_cache.scala 30:26]
  reg  valid_0_33; // @[d_cache.scala 30:26]
  reg  valid_0_34; // @[d_cache.scala 30:26]
  reg  valid_0_35; // @[d_cache.scala 30:26]
  reg  valid_0_36; // @[d_cache.scala 30:26]
  reg  valid_0_37; // @[d_cache.scala 30:26]
  reg  valid_0_38; // @[d_cache.scala 30:26]
  reg  valid_0_39; // @[d_cache.scala 30:26]
  reg  valid_0_40; // @[d_cache.scala 30:26]
  reg  valid_0_41; // @[d_cache.scala 30:26]
  reg  valid_0_42; // @[d_cache.scala 30:26]
  reg  valid_0_43; // @[d_cache.scala 30:26]
  reg  valid_0_44; // @[d_cache.scala 30:26]
  reg  valid_0_45; // @[d_cache.scala 30:26]
  reg  valid_0_46; // @[d_cache.scala 30:26]
  reg  valid_0_47; // @[d_cache.scala 30:26]
  reg  valid_0_48; // @[d_cache.scala 30:26]
  reg  valid_0_49; // @[d_cache.scala 30:26]
  reg  valid_0_50; // @[d_cache.scala 30:26]
  reg  valid_0_51; // @[d_cache.scala 30:26]
  reg  valid_0_52; // @[d_cache.scala 30:26]
  reg  valid_0_53; // @[d_cache.scala 30:26]
  reg  valid_0_54; // @[d_cache.scala 30:26]
  reg  valid_0_55; // @[d_cache.scala 30:26]
  reg  valid_0_56; // @[d_cache.scala 30:26]
  reg  valid_0_57; // @[d_cache.scala 30:26]
  reg  valid_0_58; // @[d_cache.scala 30:26]
  reg  valid_0_59; // @[d_cache.scala 30:26]
  reg  valid_0_60; // @[d_cache.scala 30:26]
  reg  valid_0_61; // @[d_cache.scala 30:26]
  reg  valid_0_62; // @[d_cache.scala 30:26]
  reg  valid_0_63; // @[d_cache.scala 30:26]
  reg  valid_0_64; // @[d_cache.scala 30:26]
  reg  valid_0_65; // @[d_cache.scala 30:26]
  reg  valid_0_66; // @[d_cache.scala 30:26]
  reg  valid_0_67; // @[d_cache.scala 30:26]
  reg  valid_0_68; // @[d_cache.scala 30:26]
  reg  valid_0_69; // @[d_cache.scala 30:26]
  reg  valid_0_70; // @[d_cache.scala 30:26]
  reg  valid_0_71; // @[d_cache.scala 30:26]
  reg  valid_0_72; // @[d_cache.scala 30:26]
  reg  valid_0_73; // @[d_cache.scala 30:26]
  reg  valid_0_74; // @[d_cache.scala 30:26]
  reg  valid_0_75; // @[d_cache.scala 30:26]
  reg  valid_0_76; // @[d_cache.scala 30:26]
  reg  valid_0_77; // @[d_cache.scala 30:26]
  reg  valid_0_78; // @[d_cache.scala 30:26]
  reg  valid_0_79; // @[d_cache.scala 30:26]
  reg  valid_0_80; // @[d_cache.scala 30:26]
  reg  valid_0_81; // @[d_cache.scala 30:26]
  reg  valid_0_82; // @[d_cache.scala 30:26]
  reg  valid_0_83; // @[d_cache.scala 30:26]
  reg  valid_0_84; // @[d_cache.scala 30:26]
  reg  valid_0_85; // @[d_cache.scala 30:26]
  reg  valid_0_86; // @[d_cache.scala 30:26]
  reg  valid_0_87; // @[d_cache.scala 30:26]
  reg  valid_0_88; // @[d_cache.scala 30:26]
  reg  valid_0_89; // @[d_cache.scala 30:26]
  reg  valid_0_90; // @[d_cache.scala 30:26]
  reg  valid_0_91; // @[d_cache.scala 30:26]
  reg  valid_0_92; // @[d_cache.scala 30:26]
  reg  valid_0_93; // @[d_cache.scala 30:26]
  reg  valid_0_94; // @[d_cache.scala 30:26]
  reg  valid_0_95; // @[d_cache.scala 30:26]
  reg  valid_0_96; // @[d_cache.scala 30:26]
  reg  valid_0_97; // @[d_cache.scala 30:26]
  reg  valid_0_98; // @[d_cache.scala 30:26]
  reg  valid_0_99; // @[d_cache.scala 30:26]
  reg  valid_0_100; // @[d_cache.scala 30:26]
  reg  valid_0_101; // @[d_cache.scala 30:26]
  reg  valid_0_102; // @[d_cache.scala 30:26]
  reg  valid_0_103; // @[d_cache.scala 30:26]
  reg  valid_0_104; // @[d_cache.scala 30:26]
  reg  valid_0_105; // @[d_cache.scala 30:26]
  reg  valid_0_106; // @[d_cache.scala 30:26]
  reg  valid_0_107; // @[d_cache.scala 30:26]
  reg  valid_0_108; // @[d_cache.scala 30:26]
  reg  valid_0_109; // @[d_cache.scala 30:26]
  reg  valid_0_110; // @[d_cache.scala 30:26]
  reg  valid_0_111; // @[d_cache.scala 30:26]
  reg  valid_0_112; // @[d_cache.scala 30:26]
  reg  valid_0_113; // @[d_cache.scala 30:26]
  reg  valid_0_114; // @[d_cache.scala 30:26]
  reg  valid_0_115; // @[d_cache.scala 30:26]
  reg  valid_0_116; // @[d_cache.scala 30:26]
  reg  valid_0_117; // @[d_cache.scala 30:26]
  reg  valid_0_118; // @[d_cache.scala 30:26]
  reg  valid_0_119; // @[d_cache.scala 30:26]
  reg  valid_0_120; // @[d_cache.scala 30:26]
  reg  valid_0_121; // @[d_cache.scala 30:26]
  reg  valid_0_122; // @[d_cache.scala 30:26]
  reg  valid_0_123; // @[d_cache.scala 30:26]
  reg  valid_0_124; // @[d_cache.scala 30:26]
  reg  valid_0_125; // @[d_cache.scala 30:26]
  reg  valid_0_126; // @[d_cache.scala 30:26]
  reg  valid_0_127; // @[d_cache.scala 30:26]
  reg  valid_1_0; // @[d_cache.scala 31:26]
  reg  valid_1_1; // @[d_cache.scala 31:26]
  reg  valid_1_2; // @[d_cache.scala 31:26]
  reg  valid_1_3; // @[d_cache.scala 31:26]
  reg  valid_1_4; // @[d_cache.scala 31:26]
  reg  valid_1_5; // @[d_cache.scala 31:26]
  reg  valid_1_6; // @[d_cache.scala 31:26]
  reg  valid_1_7; // @[d_cache.scala 31:26]
  reg  valid_1_8; // @[d_cache.scala 31:26]
  reg  valid_1_9; // @[d_cache.scala 31:26]
  reg  valid_1_10; // @[d_cache.scala 31:26]
  reg  valid_1_11; // @[d_cache.scala 31:26]
  reg  valid_1_12; // @[d_cache.scala 31:26]
  reg  valid_1_13; // @[d_cache.scala 31:26]
  reg  valid_1_14; // @[d_cache.scala 31:26]
  reg  valid_1_15; // @[d_cache.scala 31:26]
  reg  valid_1_16; // @[d_cache.scala 31:26]
  reg  valid_1_17; // @[d_cache.scala 31:26]
  reg  valid_1_18; // @[d_cache.scala 31:26]
  reg  valid_1_19; // @[d_cache.scala 31:26]
  reg  valid_1_20; // @[d_cache.scala 31:26]
  reg  valid_1_21; // @[d_cache.scala 31:26]
  reg  valid_1_22; // @[d_cache.scala 31:26]
  reg  valid_1_23; // @[d_cache.scala 31:26]
  reg  valid_1_24; // @[d_cache.scala 31:26]
  reg  valid_1_25; // @[d_cache.scala 31:26]
  reg  valid_1_26; // @[d_cache.scala 31:26]
  reg  valid_1_27; // @[d_cache.scala 31:26]
  reg  valid_1_28; // @[d_cache.scala 31:26]
  reg  valid_1_29; // @[d_cache.scala 31:26]
  reg  valid_1_30; // @[d_cache.scala 31:26]
  reg  valid_1_31; // @[d_cache.scala 31:26]
  reg  valid_1_32; // @[d_cache.scala 31:26]
  reg  valid_1_33; // @[d_cache.scala 31:26]
  reg  valid_1_34; // @[d_cache.scala 31:26]
  reg  valid_1_35; // @[d_cache.scala 31:26]
  reg  valid_1_36; // @[d_cache.scala 31:26]
  reg  valid_1_37; // @[d_cache.scala 31:26]
  reg  valid_1_38; // @[d_cache.scala 31:26]
  reg  valid_1_39; // @[d_cache.scala 31:26]
  reg  valid_1_40; // @[d_cache.scala 31:26]
  reg  valid_1_41; // @[d_cache.scala 31:26]
  reg  valid_1_42; // @[d_cache.scala 31:26]
  reg  valid_1_43; // @[d_cache.scala 31:26]
  reg  valid_1_44; // @[d_cache.scala 31:26]
  reg  valid_1_45; // @[d_cache.scala 31:26]
  reg  valid_1_46; // @[d_cache.scala 31:26]
  reg  valid_1_47; // @[d_cache.scala 31:26]
  reg  valid_1_48; // @[d_cache.scala 31:26]
  reg  valid_1_49; // @[d_cache.scala 31:26]
  reg  valid_1_50; // @[d_cache.scala 31:26]
  reg  valid_1_51; // @[d_cache.scala 31:26]
  reg  valid_1_52; // @[d_cache.scala 31:26]
  reg  valid_1_53; // @[d_cache.scala 31:26]
  reg  valid_1_54; // @[d_cache.scala 31:26]
  reg  valid_1_55; // @[d_cache.scala 31:26]
  reg  valid_1_56; // @[d_cache.scala 31:26]
  reg  valid_1_57; // @[d_cache.scala 31:26]
  reg  valid_1_58; // @[d_cache.scala 31:26]
  reg  valid_1_59; // @[d_cache.scala 31:26]
  reg  valid_1_60; // @[d_cache.scala 31:26]
  reg  valid_1_61; // @[d_cache.scala 31:26]
  reg  valid_1_62; // @[d_cache.scala 31:26]
  reg  valid_1_63; // @[d_cache.scala 31:26]
  reg  valid_1_64; // @[d_cache.scala 31:26]
  reg  valid_1_65; // @[d_cache.scala 31:26]
  reg  valid_1_66; // @[d_cache.scala 31:26]
  reg  valid_1_67; // @[d_cache.scala 31:26]
  reg  valid_1_68; // @[d_cache.scala 31:26]
  reg  valid_1_69; // @[d_cache.scala 31:26]
  reg  valid_1_70; // @[d_cache.scala 31:26]
  reg  valid_1_71; // @[d_cache.scala 31:26]
  reg  valid_1_72; // @[d_cache.scala 31:26]
  reg  valid_1_73; // @[d_cache.scala 31:26]
  reg  valid_1_74; // @[d_cache.scala 31:26]
  reg  valid_1_75; // @[d_cache.scala 31:26]
  reg  valid_1_76; // @[d_cache.scala 31:26]
  reg  valid_1_77; // @[d_cache.scala 31:26]
  reg  valid_1_78; // @[d_cache.scala 31:26]
  reg  valid_1_79; // @[d_cache.scala 31:26]
  reg  valid_1_80; // @[d_cache.scala 31:26]
  reg  valid_1_81; // @[d_cache.scala 31:26]
  reg  valid_1_82; // @[d_cache.scala 31:26]
  reg  valid_1_83; // @[d_cache.scala 31:26]
  reg  valid_1_84; // @[d_cache.scala 31:26]
  reg  valid_1_85; // @[d_cache.scala 31:26]
  reg  valid_1_86; // @[d_cache.scala 31:26]
  reg  valid_1_87; // @[d_cache.scala 31:26]
  reg  valid_1_88; // @[d_cache.scala 31:26]
  reg  valid_1_89; // @[d_cache.scala 31:26]
  reg  valid_1_90; // @[d_cache.scala 31:26]
  reg  valid_1_91; // @[d_cache.scala 31:26]
  reg  valid_1_92; // @[d_cache.scala 31:26]
  reg  valid_1_93; // @[d_cache.scala 31:26]
  reg  valid_1_94; // @[d_cache.scala 31:26]
  reg  valid_1_95; // @[d_cache.scala 31:26]
  reg  valid_1_96; // @[d_cache.scala 31:26]
  reg  valid_1_97; // @[d_cache.scala 31:26]
  reg  valid_1_98; // @[d_cache.scala 31:26]
  reg  valid_1_99; // @[d_cache.scala 31:26]
  reg  valid_1_100; // @[d_cache.scala 31:26]
  reg  valid_1_101; // @[d_cache.scala 31:26]
  reg  valid_1_102; // @[d_cache.scala 31:26]
  reg  valid_1_103; // @[d_cache.scala 31:26]
  reg  valid_1_104; // @[d_cache.scala 31:26]
  reg  valid_1_105; // @[d_cache.scala 31:26]
  reg  valid_1_106; // @[d_cache.scala 31:26]
  reg  valid_1_107; // @[d_cache.scala 31:26]
  reg  valid_1_108; // @[d_cache.scala 31:26]
  reg  valid_1_109; // @[d_cache.scala 31:26]
  reg  valid_1_110; // @[d_cache.scala 31:26]
  reg  valid_1_111; // @[d_cache.scala 31:26]
  reg  valid_1_112; // @[d_cache.scala 31:26]
  reg  valid_1_113; // @[d_cache.scala 31:26]
  reg  valid_1_114; // @[d_cache.scala 31:26]
  reg  valid_1_115; // @[d_cache.scala 31:26]
  reg  valid_1_116; // @[d_cache.scala 31:26]
  reg  valid_1_117; // @[d_cache.scala 31:26]
  reg  valid_1_118; // @[d_cache.scala 31:26]
  reg  valid_1_119; // @[d_cache.scala 31:26]
  reg  valid_1_120; // @[d_cache.scala 31:26]
  reg  valid_1_121; // @[d_cache.scala 31:26]
  reg  valid_1_122; // @[d_cache.scala 31:26]
  reg  valid_1_123; // @[d_cache.scala 31:26]
  reg  valid_1_124; // @[d_cache.scala 31:26]
  reg  valid_1_125; // @[d_cache.scala 31:26]
  reg  valid_1_126; // @[d_cache.scala 31:26]
  reg  valid_1_127; // @[d_cache.scala 31:26]
  reg  dirty_0_0; // @[d_cache.scala 32:26]
  reg  dirty_0_1; // @[d_cache.scala 32:26]
  reg  dirty_0_2; // @[d_cache.scala 32:26]
  reg  dirty_0_3; // @[d_cache.scala 32:26]
  reg  dirty_0_4; // @[d_cache.scala 32:26]
  reg  dirty_0_5; // @[d_cache.scala 32:26]
  reg  dirty_0_6; // @[d_cache.scala 32:26]
  reg  dirty_0_7; // @[d_cache.scala 32:26]
  reg  dirty_0_8; // @[d_cache.scala 32:26]
  reg  dirty_0_9; // @[d_cache.scala 32:26]
  reg  dirty_0_10; // @[d_cache.scala 32:26]
  reg  dirty_0_11; // @[d_cache.scala 32:26]
  reg  dirty_0_12; // @[d_cache.scala 32:26]
  reg  dirty_0_13; // @[d_cache.scala 32:26]
  reg  dirty_0_14; // @[d_cache.scala 32:26]
  reg  dirty_0_15; // @[d_cache.scala 32:26]
  reg  dirty_0_16; // @[d_cache.scala 32:26]
  reg  dirty_0_17; // @[d_cache.scala 32:26]
  reg  dirty_0_18; // @[d_cache.scala 32:26]
  reg  dirty_0_19; // @[d_cache.scala 32:26]
  reg  dirty_0_20; // @[d_cache.scala 32:26]
  reg  dirty_0_21; // @[d_cache.scala 32:26]
  reg  dirty_0_22; // @[d_cache.scala 32:26]
  reg  dirty_0_23; // @[d_cache.scala 32:26]
  reg  dirty_0_24; // @[d_cache.scala 32:26]
  reg  dirty_0_25; // @[d_cache.scala 32:26]
  reg  dirty_0_26; // @[d_cache.scala 32:26]
  reg  dirty_0_27; // @[d_cache.scala 32:26]
  reg  dirty_0_28; // @[d_cache.scala 32:26]
  reg  dirty_0_29; // @[d_cache.scala 32:26]
  reg  dirty_0_30; // @[d_cache.scala 32:26]
  reg  dirty_0_31; // @[d_cache.scala 32:26]
  reg  dirty_0_32; // @[d_cache.scala 32:26]
  reg  dirty_0_33; // @[d_cache.scala 32:26]
  reg  dirty_0_34; // @[d_cache.scala 32:26]
  reg  dirty_0_35; // @[d_cache.scala 32:26]
  reg  dirty_0_36; // @[d_cache.scala 32:26]
  reg  dirty_0_37; // @[d_cache.scala 32:26]
  reg  dirty_0_38; // @[d_cache.scala 32:26]
  reg  dirty_0_39; // @[d_cache.scala 32:26]
  reg  dirty_0_40; // @[d_cache.scala 32:26]
  reg  dirty_0_41; // @[d_cache.scala 32:26]
  reg  dirty_0_42; // @[d_cache.scala 32:26]
  reg  dirty_0_43; // @[d_cache.scala 32:26]
  reg  dirty_0_44; // @[d_cache.scala 32:26]
  reg  dirty_0_45; // @[d_cache.scala 32:26]
  reg  dirty_0_46; // @[d_cache.scala 32:26]
  reg  dirty_0_47; // @[d_cache.scala 32:26]
  reg  dirty_0_48; // @[d_cache.scala 32:26]
  reg  dirty_0_49; // @[d_cache.scala 32:26]
  reg  dirty_0_50; // @[d_cache.scala 32:26]
  reg  dirty_0_51; // @[d_cache.scala 32:26]
  reg  dirty_0_52; // @[d_cache.scala 32:26]
  reg  dirty_0_53; // @[d_cache.scala 32:26]
  reg  dirty_0_54; // @[d_cache.scala 32:26]
  reg  dirty_0_55; // @[d_cache.scala 32:26]
  reg  dirty_0_56; // @[d_cache.scala 32:26]
  reg  dirty_0_57; // @[d_cache.scala 32:26]
  reg  dirty_0_58; // @[d_cache.scala 32:26]
  reg  dirty_0_59; // @[d_cache.scala 32:26]
  reg  dirty_0_60; // @[d_cache.scala 32:26]
  reg  dirty_0_61; // @[d_cache.scala 32:26]
  reg  dirty_0_62; // @[d_cache.scala 32:26]
  reg  dirty_0_63; // @[d_cache.scala 32:26]
  reg  dirty_0_64; // @[d_cache.scala 32:26]
  reg  dirty_0_65; // @[d_cache.scala 32:26]
  reg  dirty_0_66; // @[d_cache.scala 32:26]
  reg  dirty_0_67; // @[d_cache.scala 32:26]
  reg  dirty_0_68; // @[d_cache.scala 32:26]
  reg  dirty_0_69; // @[d_cache.scala 32:26]
  reg  dirty_0_70; // @[d_cache.scala 32:26]
  reg  dirty_0_71; // @[d_cache.scala 32:26]
  reg  dirty_0_72; // @[d_cache.scala 32:26]
  reg  dirty_0_73; // @[d_cache.scala 32:26]
  reg  dirty_0_74; // @[d_cache.scala 32:26]
  reg  dirty_0_75; // @[d_cache.scala 32:26]
  reg  dirty_0_76; // @[d_cache.scala 32:26]
  reg  dirty_0_77; // @[d_cache.scala 32:26]
  reg  dirty_0_78; // @[d_cache.scala 32:26]
  reg  dirty_0_79; // @[d_cache.scala 32:26]
  reg  dirty_0_80; // @[d_cache.scala 32:26]
  reg  dirty_0_81; // @[d_cache.scala 32:26]
  reg  dirty_0_82; // @[d_cache.scala 32:26]
  reg  dirty_0_83; // @[d_cache.scala 32:26]
  reg  dirty_0_84; // @[d_cache.scala 32:26]
  reg  dirty_0_85; // @[d_cache.scala 32:26]
  reg  dirty_0_86; // @[d_cache.scala 32:26]
  reg  dirty_0_87; // @[d_cache.scala 32:26]
  reg  dirty_0_88; // @[d_cache.scala 32:26]
  reg  dirty_0_89; // @[d_cache.scala 32:26]
  reg  dirty_0_90; // @[d_cache.scala 32:26]
  reg  dirty_0_91; // @[d_cache.scala 32:26]
  reg  dirty_0_92; // @[d_cache.scala 32:26]
  reg  dirty_0_93; // @[d_cache.scala 32:26]
  reg  dirty_0_94; // @[d_cache.scala 32:26]
  reg  dirty_0_95; // @[d_cache.scala 32:26]
  reg  dirty_0_96; // @[d_cache.scala 32:26]
  reg  dirty_0_97; // @[d_cache.scala 32:26]
  reg  dirty_0_98; // @[d_cache.scala 32:26]
  reg  dirty_0_99; // @[d_cache.scala 32:26]
  reg  dirty_0_100; // @[d_cache.scala 32:26]
  reg  dirty_0_101; // @[d_cache.scala 32:26]
  reg  dirty_0_102; // @[d_cache.scala 32:26]
  reg  dirty_0_103; // @[d_cache.scala 32:26]
  reg  dirty_0_104; // @[d_cache.scala 32:26]
  reg  dirty_0_105; // @[d_cache.scala 32:26]
  reg  dirty_0_106; // @[d_cache.scala 32:26]
  reg  dirty_0_107; // @[d_cache.scala 32:26]
  reg  dirty_0_108; // @[d_cache.scala 32:26]
  reg  dirty_0_109; // @[d_cache.scala 32:26]
  reg  dirty_0_110; // @[d_cache.scala 32:26]
  reg  dirty_0_111; // @[d_cache.scala 32:26]
  reg  dirty_0_112; // @[d_cache.scala 32:26]
  reg  dirty_0_113; // @[d_cache.scala 32:26]
  reg  dirty_0_114; // @[d_cache.scala 32:26]
  reg  dirty_0_115; // @[d_cache.scala 32:26]
  reg  dirty_0_116; // @[d_cache.scala 32:26]
  reg  dirty_0_117; // @[d_cache.scala 32:26]
  reg  dirty_0_118; // @[d_cache.scala 32:26]
  reg  dirty_0_119; // @[d_cache.scala 32:26]
  reg  dirty_0_120; // @[d_cache.scala 32:26]
  reg  dirty_0_121; // @[d_cache.scala 32:26]
  reg  dirty_0_122; // @[d_cache.scala 32:26]
  reg  dirty_0_123; // @[d_cache.scala 32:26]
  reg  dirty_0_124; // @[d_cache.scala 32:26]
  reg  dirty_0_125; // @[d_cache.scala 32:26]
  reg  dirty_0_126; // @[d_cache.scala 32:26]
  reg  dirty_0_127; // @[d_cache.scala 32:26]
  reg  dirty_1_0; // @[d_cache.scala 33:26]
  reg  dirty_1_1; // @[d_cache.scala 33:26]
  reg  dirty_1_2; // @[d_cache.scala 33:26]
  reg  dirty_1_3; // @[d_cache.scala 33:26]
  reg  dirty_1_4; // @[d_cache.scala 33:26]
  reg  dirty_1_5; // @[d_cache.scala 33:26]
  reg  dirty_1_6; // @[d_cache.scala 33:26]
  reg  dirty_1_7; // @[d_cache.scala 33:26]
  reg  dirty_1_8; // @[d_cache.scala 33:26]
  reg  dirty_1_9; // @[d_cache.scala 33:26]
  reg  dirty_1_10; // @[d_cache.scala 33:26]
  reg  dirty_1_11; // @[d_cache.scala 33:26]
  reg  dirty_1_12; // @[d_cache.scala 33:26]
  reg  dirty_1_13; // @[d_cache.scala 33:26]
  reg  dirty_1_14; // @[d_cache.scala 33:26]
  reg  dirty_1_15; // @[d_cache.scala 33:26]
  reg  dirty_1_16; // @[d_cache.scala 33:26]
  reg  dirty_1_17; // @[d_cache.scala 33:26]
  reg  dirty_1_18; // @[d_cache.scala 33:26]
  reg  dirty_1_19; // @[d_cache.scala 33:26]
  reg  dirty_1_20; // @[d_cache.scala 33:26]
  reg  dirty_1_21; // @[d_cache.scala 33:26]
  reg  dirty_1_22; // @[d_cache.scala 33:26]
  reg  dirty_1_23; // @[d_cache.scala 33:26]
  reg  dirty_1_24; // @[d_cache.scala 33:26]
  reg  dirty_1_25; // @[d_cache.scala 33:26]
  reg  dirty_1_26; // @[d_cache.scala 33:26]
  reg  dirty_1_27; // @[d_cache.scala 33:26]
  reg  dirty_1_28; // @[d_cache.scala 33:26]
  reg  dirty_1_29; // @[d_cache.scala 33:26]
  reg  dirty_1_30; // @[d_cache.scala 33:26]
  reg  dirty_1_31; // @[d_cache.scala 33:26]
  reg  dirty_1_32; // @[d_cache.scala 33:26]
  reg  dirty_1_33; // @[d_cache.scala 33:26]
  reg  dirty_1_34; // @[d_cache.scala 33:26]
  reg  dirty_1_35; // @[d_cache.scala 33:26]
  reg  dirty_1_36; // @[d_cache.scala 33:26]
  reg  dirty_1_37; // @[d_cache.scala 33:26]
  reg  dirty_1_38; // @[d_cache.scala 33:26]
  reg  dirty_1_39; // @[d_cache.scala 33:26]
  reg  dirty_1_40; // @[d_cache.scala 33:26]
  reg  dirty_1_41; // @[d_cache.scala 33:26]
  reg  dirty_1_42; // @[d_cache.scala 33:26]
  reg  dirty_1_43; // @[d_cache.scala 33:26]
  reg  dirty_1_44; // @[d_cache.scala 33:26]
  reg  dirty_1_45; // @[d_cache.scala 33:26]
  reg  dirty_1_46; // @[d_cache.scala 33:26]
  reg  dirty_1_47; // @[d_cache.scala 33:26]
  reg  dirty_1_48; // @[d_cache.scala 33:26]
  reg  dirty_1_49; // @[d_cache.scala 33:26]
  reg  dirty_1_50; // @[d_cache.scala 33:26]
  reg  dirty_1_51; // @[d_cache.scala 33:26]
  reg  dirty_1_52; // @[d_cache.scala 33:26]
  reg  dirty_1_53; // @[d_cache.scala 33:26]
  reg  dirty_1_54; // @[d_cache.scala 33:26]
  reg  dirty_1_55; // @[d_cache.scala 33:26]
  reg  dirty_1_56; // @[d_cache.scala 33:26]
  reg  dirty_1_57; // @[d_cache.scala 33:26]
  reg  dirty_1_58; // @[d_cache.scala 33:26]
  reg  dirty_1_59; // @[d_cache.scala 33:26]
  reg  dirty_1_60; // @[d_cache.scala 33:26]
  reg  dirty_1_61; // @[d_cache.scala 33:26]
  reg  dirty_1_62; // @[d_cache.scala 33:26]
  reg  dirty_1_63; // @[d_cache.scala 33:26]
  reg  dirty_1_64; // @[d_cache.scala 33:26]
  reg  dirty_1_65; // @[d_cache.scala 33:26]
  reg  dirty_1_66; // @[d_cache.scala 33:26]
  reg  dirty_1_67; // @[d_cache.scala 33:26]
  reg  dirty_1_68; // @[d_cache.scala 33:26]
  reg  dirty_1_69; // @[d_cache.scala 33:26]
  reg  dirty_1_70; // @[d_cache.scala 33:26]
  reg  dirty_1_71; // @[d_cache.scala 33:26]
  reg  dirty_1_72; // @[d_cache.scala 33:26]
  reg  dirty_1_73; // @[d_cache.scala 33:26]
  reg  dirty_1_74; // @[d_cache.scala 33:26]
  reg  dirty_1_75; // @[d_cache.scala 33:26]
  reg  dirty_1_76; // @[d_cache.scala 33:26]
  reg  dirty_1_77; // @[d_cache.scala 33:26]
  reg  dirty_1_78; // @[d_cache.scala 33:26]
  reg  dirty_1_79; // @[d_cache.scala 33:26]
  reg  dirty_1_80; // @[d_cache.scala 33:26]
  reg  dirty_1_81; // @[d_cache.scala 33:26]
  reg  dirty_1_82; // @[d_cache.scala 33:26]
  reg  dirty_1_83; // @[d_cache.scala 33:26]
  reg  dirty_1_84; // @[d_cache.scala 33:26]
  reg  dirty_1_85; // @[d_cache.scala 33:26]
  reg  dirty_1_86; // @[d_cache.scala 33:26]
  reg  dirty_1_87; // @[d_cache.scala 33:26]
  reg  dirty_1_88; // @[d_cache.scala 33:26]
  reg  dirty_1_89; // @[d_cache.scala 33:26]
  reg  dirty_1_90; // @[d_cache.scala 33:26]
  reg  dirty_1_91; // @[d_cache.scala 33:26]
  reg  dirty_1_92; // @[d_cache.scala 33:26]
  reg  dirty_1_93; // @[d_cache.scala 33:26]
  reg  dirty_1_94; // @[d_cache.scala 33:26]
  reg  dirty_1_95; // @[d_cache.scala 33:26]
  reg  dirty_1_96; // @[d_cache.scala 33:26]
  reg  dirty_1_97; // @[d_cache.scala 33:26]
  reg  dirty_1_98; // @[d_cache.scala 33:26]
  reg  dirty_1_99; // @[d_cache.scala 33:26]
  reg  dirty_1_100; // @[d_cache.scala 33:26]
  reg  dirty_1_101; // @[d_cache.scala 33:26]
  reg  dirty_1_102; // @[d_cache.scala 33:26]
  reg  dirty_1_103; // @[d_cache.scala 33:26]
  reg  dirty_1_104; // @[d_cache.scala 33:26]
  reg  dirty_1_105; // @[d_cache.scala 33:26]
  reg  dirty_1_106; // @[d_cache.scala 33:26]
  reg  dirty_1_107; // @[d_cache.scala 33:26]
  reg  dirty_1_108; // @[d_cache.scala 33:26]
  reg  dirty_1_109; // @[d_cache.scala 33:26]
  reg  dirty_1_110; // @[d_cache.scala 33:26]
  reg  dirty_1_111; // @[d_cache.scala 33:26]
  reg  dirty_1_112; // @[d_cache.scala 33:26]
  reg  dirty_1_113; // @[d_cache.scala 33:26]
  reg  dirty_1_114; // @[d_cache.scala 33:26]
  reg  dirty_1_115; // @[d_cache.scala 33:26]
  reg  dirty_1_116; // @[d_cache.scala 33:26]
  reg  dirty_1_117; // @[d_cache.scala 33:26]
  reg  dirty_1_118; // @[d_cache.scala 33:26]
  reg  dirty_1_119; // @[d_cache.scala 33:26]
  reg  dirty_1_120; // @[d_cache.scala 33:26]
  reg  dirty_1_121; // @[d_cache.scala 33:26]
  reg  dirty_1_122; // @[d_cache.scala 33:26]
  reg  dirty_1_123; // @[d_cache.scala 33:26]
  reg  dirty_1_124; // @[d_cache.scala 33:26]
  reg  dirty_1_125; // @[d_cache.scala 33:26]
  reg  dirty_1_126; // @[d_cache.scala 33:26]
  reg  dirty_1_127; // @[d_cache.scala 33:26]
  reg  way0_hit; // @[d_cache.scala 34:27]
  reg  way1_hit; // @[d_cache.scala 35:27]
  reg [63:0] write_back_data; // @[d_cache.scala 37:34]
  reg [31:0] write_back_addr; // @[d_cache.scala 38:34]
  reg [1:0] unuse_way; // @[d_cache.scala 41:28]
  reg [63:0] receive_data; // @[d_cache.scala 42:31]
  reg  quene; // @[d_cache.scala 43:24]
  wire [2:0] offset = io_from_lsu_araddr[2:0]; // @[d_cache.scala 45:36]
  wire [6:0] index = io_from_lsu_araddr[9:3]; // @[d_cache.scala 46:35]
  wire [21:0] tag = io_from_lsu_araddr[31:10]; // @[d_cache.scala 47:33]
  wire [5:0] _shift_bit_T_8 = offset == 3'h7 ? 6'h38 : 6'h0; // @[d_cache.scala 56:24]
  wire [5:0] _shift_bit_T_9 = offset == 3'h6 ? 6'h30 : _shift_bit_T_8; // @[d_cache.scala 55:24]
  wire [5:0] _shift_bit_T_10 = offset == 3'h5 ? 6'h28 : _shift_bit_T_9; // @[d_cache.scala 54:24]
  wire [5:0] _shift_bit_T_11 = offset == 3'h4 ? 6'h20 : _shift_bit_T_10; // @[d_cache.scala 53:24]
  wire [5:0] _shift_bit_T_12 = offset == 3'h3 ? 6'h18 : _shift_bit_T_11; // @[d_cache.scala 52:24]
  wire [5:0] _shift_bit_T_13 = offset == 3'h2 ? 6'h10 : _shift_bit_T_12; // @[d_cache.scala 51:24]
  wire [5:0] _shift_bit_T_14 = offset == 3'h1 ? 6'h8 : _shift_bit_T_13; // @[d_cache.scala 50:24]
  wire [5:0] shift_bit = offset == 3'h0 ? 6'h0 : _shift_bit_T_14; // @[d_cache.scala 49:24]
  wire [63:0] _wmask_T_4 = io_from_lsu_wstrb == 8'hff ? 64'hffffffffffffffff : 64'h0; // @[d_cache.scala 61:20]
  wire [63:0] _wmask_T_5 = io_from_lsu_wstrb == 8'hf ? 64'hffffffff : _wmask_T_4; // @[d_cache.scala 60:20]
  wire [63:0] _wmask_T_6 = io_from_lsu_wstrb == 8'h3 ? 64'hffff : _wmask_T_5; // @[d_cache.scala 59:20]
  wire [63:0] wmask = io_from_lsu_wstrb == 8'h1 ? 64'hff : _wmask_T_6; // @[d_cache.scala 58:20]
  wire [31:0] _GEN_1 = 7'h1 == index ? tag_0_1 : tag_0_0; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_2 = 7'h2 == index ? tag_0_2 : _GEN_1; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_3 = 7'h3 == index ? tag_0_3 : _GEN_2; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_4 = 7'h4 == index ? tag_0_4 : _GEN_3; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_5 = 7'h5 == index ? tag_0_5 : _GEN_4; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_6 = 7'h6 == index ? tag_0_6 : _GEN_5; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_7 = 7'h7 == index ? tag_0_7 : _GEN_6; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_8 = 7'h8 == index ? tag_0_8 : _GEN_7; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_9 = 7'h9 == index ? tag_0_9 : _GEN_8; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_10 = 7'ha == index ? tag_0_10 : _GEN_9; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_11 = 7'hb == index ? tag_0_11 : _GEN_10; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_12 = 7'hc == index ? tag_0_12 : _GEN_11; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_13 = 7'hd == index ? tag_0_13 : _GEN_12; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_14 = 7'he == index ? tag_0_14 : _GEN_13; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_15 = 7'hf == index ? tag_0_15 : _GEN_14; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_16 = 7'h10 == index ? tag_0_16 : _GEN_15; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_17 = 7'h11 == index ? tag_0_17 : _GEN_16; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_18 = 7'h12 == index ? tag_0_18 : _GEN_17; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_19 = 7'h13 == index ? tag_0_19 : _GEN_18; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_20 = 7'h14 == index ? tag_0_20 : _GEN_19; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_21 = 7'h15 == index ? tag_0_21 : _GEN_20; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_22 = 7'h16 == index ? tag_0_22 : _GEN_21; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_23 = 7'h17 == index ? tag_0_23 : _GEN_22; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_24 = 7'h18 == index ? tag_0_24 : _GEN_23; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_25 = 7'h19 == index ? tag_0_25 : _GEN_24; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_26 = 7'h1a == index ? tag_0_26 : _GEN_25; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_27 = 7'h1b == index ? tag_0_27 : _GEN_26; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_28 = 7'h1c == index ? tag_0_28 : _GEN_27; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_29 = 7'h1d == index ? tag_0_29 : _GEN_28; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_30 = 7'h1e == index ? tag_0_30 : _GEN_29; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_31 = 7'h1f == index ? tag_0_31 : _GEN_30; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_32 = 7'h20 == index ? tag_0_32 : _GEN_31; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_33 = 7'h21 == index ? tag_0_33 : _GEN_32; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_34 = 7'h22 == index ? tag_0_34 : _GEN_33; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_35 = 7'h23 == index ? tag_0_35 : _GEN_34; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_36 = 7'h24 == index ? tag_0_36 : _GEN_35; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_37 = 7'h25 == index ? tag_0_37 : _GEN_36; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_38 = 7'h26 == index ? tag_0_38 : _GEN_37; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_39 = 7'h27 == index ? tag_0_39 : _GEN_38; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_40 = 7'h28 == index ? tag_0_40 : _GEN_39; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_41 = 7'h29 == index ? tag_0_41 : _GEN_40; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_42 = 7'h2a == index ? tag_0_42 : _GEN_41; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_43 = 7'h2b == index ? tag_0_43 : _GEN_42; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_44 = 7'h2c == index ? tag_0_44 : _GEN_43; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_45 = 7'h2d == index ? tag_0_45 : _GEN_44; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_46 = 7'h2e == index ? tag_0_46 : _GEN_45; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_47 = 7'h2f == index ? tag_0_47 : _GEN_46; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_48 = 7'h30 == index ? tag_0_48 : _GEN_47; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_49 = 7'h31 == index ? tag_0_49 : _GEN_48; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_50 = 7'h32 == index ? tag_0_50 : _GEN_49; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_51 = 7'h33 == index ? tag_0_51 : _GEN_50; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_52 = 7'h34 == index ? tag_0_52 : _GEN_51; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_53 = 7'h35 == index ? tag_0_53 : _GEN_52; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_54 = 7'h36 == index ? tag_0_54 : _GEN_53; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_55 = 7'h37 == index ? tag_0_55 : _GEN_54; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_56 = 7'h38 == index ? tag_0_56 : _GEN_55; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_57 = 7'h39 == index ? tag_0_57 : _GEN_56; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_58 = 7'h3a == index ? tag_0_58 : _GEN_57; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_59 = 7'h3b == index ? tag_0_59 : _GEN_58; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_60 = 7'h3c == index ? tag_0_60 : _GEN_59; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_61 = 7'h3d == index ? tag_0_61 : _GEN_60; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_62 = 7'h3e == index ? tag_0_62 : _GEN_61; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_63 = 7'h3f == index ? tag_0_63 : _GEN_62; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_64 = 7'h40 == index ? tag_0_64 : _GEN_63; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_65 = 7'h41 == index ? tag_0_65 : _GEN_64; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_66 = 7'h42 == index ? tag_0_66 : _GEN_65; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_67 = 7'h43 == index ? tag_0_67 : _GEN_66; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_68 = 7'h44 == index ? tag_0_68 : _GEN_67; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_69 = 7'h45 == index ? tag_0_69 : _GEN_68; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_70 = 7'h46 == index ? tag_0_70 : _GEN_69; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_71 = 7'h47 == index ? tag_0_71 : _GEN_70; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_72 = 7'h48 == index ? tag_0_72 : _GEN_71; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_73 = 7'h49 == index ? tag_0_73 : _GEN_72; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_74 = 7'h4a == index ? tag_0_74 : _GEN_73; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_75 = 7'h4b == index ? tag_0_75 : _GEN_74; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_76 = 7'h4c == index ? tag_0_76 : _GEN_75; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_77 = 7'h4d == index ? tag_0_77 : _GEN_76; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_78 = 7'h4e == index ? tag_0_78 : _GEN_77; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_79 = 7'h4f == index ? tag_0_79 : _GEN_78; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_80 = 7'h50 == index ? tag_0_80 : _GEN_79; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_81 = 7'h51 == index ? tag_0_81 : _GEN_80; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_82 = 7'h52 == index ? tag_0_82 : _GEN_81; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_83 = 7'h53 == index ? tag_0_83 : _GEN_82; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_84 = 7'h54 == index ? tag_0_84 : _GEN_83; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_85 = 7'h55 == index ? tag_0_85 : _GEN_84; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_86 = 7'h56 == index ? tag_0_86 : _GEN_85; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_87 = 7'h57 == index ? tag_0_87 : _GEN_86; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_88 = 7'h58 == index ? tag_0_88 : _GEN_87; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_89 = 7'h59 == index ? tag_0_89 : _GEN_88; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_90 = 7'h5a == index ? tag_0_90 : _GEN_89; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_91 = 7'h5b == index ? tag_0_91 : _GEN_90; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_92 = 7'h5c == index ? tag_0_92 : _GEN_91; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_93 = 7'h5d == index ? tag_0_93 : _GEN_92; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_94 = 7'h5e == index ? tag_0_94 : _GEN_93; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_95 = 7'h5f == index ? tag_0_95 : _GEN_94; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_96 = 7'h60 == index ? tag_0_96 : _GEN_95; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_97 = 7'h61 == index ? tag_0_97 : _GEN_96; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_98 = 7'h62 == index ? tag_0_98 : _GEN_97; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_99 = 7'h63 == index ? tag_0_99 : _GEN_98; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_100 = 7'h64 == index ? tag_0_100 : _GEN_99; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_101 = 7'h65 == index ? tag_0_101 : _GEN_100; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_102 = 7'h66 == index ? tag_0_102 : _GEN_101; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_103 = 7'h67 == index ? tag_0_103 : _GEN_102; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_104 = 7'h68 == index ? tag_0_104 : _GEN_103; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_105 = 7'h69 == index ? tag_0_105 : _GEN_104; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_106 = 7'h6a == index ? tag_0_106 : _GEN_105; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_107 = 7'h6b == index ? tag_0_107 : _GEN_106; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_108 = 7'h6c == index ? tag_0_108 : _GEN_107; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_109 = 7'h6d == index ? tag_0_109 : _GEN_108; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_110 = 7'h6e == index ? tag_0_110 : _GEN_109; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_111 = 7'h6f == index ? tag_0_111 : _GEN_110; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_112 = 7'h70 == index ? tag_0_112 : _GEN_111; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_113 = 7'h71 == index ? tag_0_113 : _GEN_112; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_114 = 7'h72 == index ? tag_0_114 : _GEN_113; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_115 = 7'h73 == index ? tag_0_115 : _GEN_114; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_116 = 7'h74 == index ? tag_0_116 : _GEN_115; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_117 = 7'h75 == index ? tag_0_117 : _GEN_116; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_118 = 7'h76 == index ? tag_0_118 : _GEN_117; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_119 = 7'h77 == index ? tag_0_119 : _GEN_118; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_120 = 7'h78 == index ? tag_0_120 : _GEN_119; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_121 = 7'h79 == index ? tag_0_121 : _GEN_120; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_122 = 7'h7a == index ? tag_0_122 : _GEN_121; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_123 = 7'h7b == index ? tag_0_123 : _GEN_122; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_124 = 7'h7c == index ? tag_0_124 : _GEN_123; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_125 = 7'h7d == index ? tag_0_125 : _GEN_124; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_126 = 7'h7e == index ? tag_0_126 : _GEN_125; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_127 = 7'h7f == index ? tag_0_127 : _GEN_126; // @[d_cache.scala 63:{24,24}]
  wire [31:0] _GEN_19745 = {{10'd0}, tag}; // @[d_cache.scala 63:24]
  wire  _GEN_129 = 7'h1 == index ? valid_0_1 : valid_0_0; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_130 = 7'h2 == index ? valid_0_2 : _GEN_129; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_131 = 7'h3 == index ? valid_0_3 : _GEN_130; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_132 = 7'h4 == index ? valid_0_4 : _GEN_131; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_133 = 7'h5 == index ? valid_0_5 : _GEN_132; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_134 = 7'h6 == index ? valid_0_6 : _GEN_133; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_135 = 7'h7 == index ? valid_0_7 : _GEN_134; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_136 = 7'h8 == index ? valid_0_8 : _GEN_135; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_137 = 7'h9 == index ? valid_0_9 : _GEN_136; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_138 = 7'ha == index ? valid_0_10 : _GEN_137; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_139 = 7'hb == index ? valid_0_11 : _GEN_138; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_140 = 7'hc == index ? valid_0_12 : _GEN_139; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_141 = 7'hd == index ? valid_0_13 : _GEN_140; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_142 = 7'he == index ? valid_0_14 : _GEN_141; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_143 = 7'hf == index ? valid_0_15 : _GEN_142; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_144 = 7'h10 == index ? valid_0_16 : _GEN_143; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_145 = 7'h11 == index ? valid_0_17 : _GEN_144; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_146 = 7'h12 == index ? valid_0_18 : _GEN_145; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_147 = 7'h13 == index ? valid_0_19 : _GEN_146; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_148 = 7'h14 == index ? valid_0_20 : _GEN_147; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_149 = 7'h15 == index ? valid_0_21 : _GEN_148; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_150 = 7'h16 == index ? valid_0_22 : _GEN_149; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_151 = 7'h17 == index ? valid_0_23 : _GEN_150; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_152 = 7'h18 == index ? valid_0_24 : _GEN_151; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_153 = 7'h19 == index ? valid_0_25 : _GEN_152; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_154 = 7'h1a == index ? valid_0_26 : _GEN_153; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_155 = 7'h1b == index ? valid_0_27 : _GEN_154; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_156 = 7'h1c == index ? valid_0_28 : _GEN_155; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_157 = 7'h1d == index ? valid_0_29 : _GEN_156; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_158 = 7'h1e == index ? valid_0_30 : _GEN_157; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_159 = 7'h1f == index ? valid_0_31 : _GEN_158; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_160 = 7'h20 == index ? valid_0_32 : _GEN_159; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_161 = 7'h21 == index ? valid_0_33 : _GEN_160; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_162 = 7'h22 == index ? valid_0_34 : _GEN_161; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_163 = 7'h23 == index ? valid_0_35 : _GEN_162; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_164 = 7'h24 == index ? valid_0_36 : _GEN_163; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_165 = 7'h25 == index ? valid_0_37 : _GEN_164; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_166 = 7'h26 == index ? valid_0_38 : _GEN_165; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_167 = 7'h27 == index ? valid_0_39 : _GEN_166; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_168 = 7'h28 == index ? valid_0_40 : _GEN_167; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_169 = 7'h29 == index ? valid_0_41 : _GEN_168; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_170 = 7'h2a == index ? valid_0_42 : _GEN_169; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_171 = 7'h2b == index ? valid_0_43 : _GEN_170; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_172 = 7'h2c == index ? valid_0_44 : _GEN_171; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_173 = 7'h2d == index ? valid_0_45 : _GEN_172; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_174 = 7'h2e == index ? valid_0_46 : _GEN_173; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_175 = 7'h2f == index ? valid_0_47 : _GEN_174; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_176 = 7'h30 == index ? valid_0_48 : _GEN_175; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_177 = 7'h31 == index ? valid_0_49 : _GEN_176; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_178 = 7'h32 == index ? valid_0_50 : _GEN_177; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_179 = 7'h33 == index ? valid_0_51 : _GEN_178; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_180 = 7'h34 == index ? valid_0_52 : _GEN_179; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_181 = 7'h35 == index ? valid_0_53 : _GEN_180; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_182 = 7'h36 == index ? valid_0_54 : _GEN_181; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_183 = 7'h37 == index ? valid_0_55 : _GEN_182; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_184 = 7'h38 == index ? valid_0_56 : _GEN_183; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_185 = 7'h39 == index ? valid_0_57 : _GEN_184; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_186 = 7'h3a == index ? valid_0_58 : _GEN_185; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_187 = 7'h3b == index ? valid_0_59 : _GEN_186; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_188 = 7'h3c == index ? valid_0_60 : _GEN_187; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_189 = 7'h3d == index ? valid_0_61 : _GEN_188; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_190 = 7'h3e == index ? valid_0_62 : _GEN_189; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_191 = 7'h3f == index ? valid_0_63 : _GEN_190; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_192 = 7'h40 == index ? valid_0_64 : _GEN_191; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_193 = 7'h41 == index ? valid_0_65 : _GEN_192; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_194 = 7'h42 == index ? valid_0_66 : _GEN_193; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_195 = 7'h43 == index ? valid_0_67 : _GEN_194; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_196 = 7'h44 == index ? valid_0_68 : _GEN_195; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_197 = 7'h45 == index ? valid_0_69 : _GEN_196; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_198 = 7'h46 == index ? valid_0_70 : _GEN_197; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_199 = 7'h47 == index ? valid_0_71 : _GEN_198; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_200 = 7'h48 == index ? valid_0_72 : _GEN_199; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_201 = 7'h49 == index ? valid_0_73 : _GEN_200; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_202 = 7'h4a == index ? valid_0_74 : _GEN_201; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_203 = 7'h4b == index ? valid_0_75 : _GEN_202; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_204 = 7'h4c == index ? valid_0_76 : _GEN_203; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_205 = 7'h4d == index ? valid_0_77 : _GEN_204; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_206 = 7'h4e == index ? valid_0_78 : _GEN_205; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_207 = 7'h4f == index ? valid_0_79 : _GEN_206; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_208 = 7'h50 == index ? valid_0_80 : _GEN_207; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_209 = 7'h51 == index ? valid_0_81 : _GEN_208; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_210 = 7'h52 == index ? valid_0_82 : _GEN_209; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_211 = 7'h53 == index ? valid_0_83 : _GEN_210; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_212 = 7'h54 == index ? valid_0_84 : _GEN_211; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_213 = 7'h55 == index ? valid_0_85 : _GEN_212; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_214 = 7'h56 == index ? valid_0_86 : _GEN_213; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_215 = 7'h57 == index ? valid_0_87 : _GEN_214; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_216 = 7'h58 == index ? valid_0_88 : _GEN_215; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_217 = 7'h59 == index ? valid_0_89 : _GEN_216; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_218 = 7'h5a == index ? valid_0_90 : _GEN_217; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_219 = 7'h5b == index ? valid_0_91 : _GEN_218; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_220 = 7'h5c == index ? valid_0_92 : _GEN_219; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_221 = 7'h5d == index ? valid_0_93 : _GEN_220; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_222 = 7'h5e == index ? valid_0_94 : _GEN_221; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_223 = 7'h5f == index ? valid_0_95 : _GEN_222; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_224 = 7'h60 == index ? valid_0_96 : _GEN_223; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_225 = 7'h61 == index ? valid_0_97 : _GEN_224; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_226 = 7'h62 == index ? valid_0_98 : _GEN_225; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_227 = 7'h63 == index ? valid_0_99 : _GEN_226; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_228 = 7'h64 == index ? valid_0_100 : _GEN_227; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_229 = 7'h65 == index ? valid_0_101 : _GEN_228; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_230 = 7'h66 == index ? valid_0_102 : _GEN_229; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_231 = 7'h67 == index ? valid_0_103 : _GEN_230; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_232 = 7'h68 == index ? valid_0_104 : _GEN_231; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_233 = 7'h69 == index ? valid_0_105 : _GEN_232; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_234 = 7'h6a == index ? valid_0_106 : _GEN_233; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_235 = 7'h6b == index ? valid_0_107 : _GEN_234; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_236 = 7'h6c == index ? valid_0_108 : _GEN_235; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_237 = 7'h6d == index ? valid_0_109 : _GEN_236; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_238 = 7'h6e == index ? valid_0_110 : _GEN_237; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_239 = 7'h6f == index ? valid_0_111 : _GEN_238; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_240 = 7'h70 == index ? valid_0_112 : _GEN_239; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_241 = 7'h71 == index ? valid_0_113 : _GEN_240; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_242 = 7'h72 == index ? valid_0_114 : _GEN_241; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_243 = 7'h73 == index ? valid_0_115 : _GEN_242; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_244 = 7'h74 == index ? valid_0_116 : _GEN_243; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_245 = 7'h75 == index ? valid_0_117 : _GEN_244; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_246 = 7'h76 == index ? valid_0_118 : _GEN_245; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_247 = 7'h77 == index ? valid_0_119 : _GEN_246; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_248 = 7'h78 == index ? valid_0_120 : _GEN_247; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_249 = 7'h79 == index ? valid_0_121 : _GEN_248; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_250 = 7'h7a == index ? valid_0_122 : _GEN_249; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_251 = 7'h7b == index ? valid_0_123 : _GEN_250; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_252 = 7'h7c == index ? valid_0_124 : _GEN_251; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_253 = 7'h7d == index ? valid_0_125 : _GEN_252; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_254 = 7'h7e == index ? valid_0_126 : _GEN_253; // @[d_cache.scala 63:{50,50}]
  wire  _GEN_255 = 7'h7f == index ? valid_0_127 : _GEN_254; // @[d_cache.scala 63:{50,50}]
  wire  _T_4 = _GEN_127 == _GEN_19745 & _GEN_255; // @[d_cache.scala 63:33]
  wire [31:0] _GEN_258 = 7'h1 == index ? tag_1_1 : tag_1_0; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_259 = 7'h2 == index ? tag_1_2 : _GEN_258; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_260 = 7'h3 == index ? tag_1_3 : _GEN_259; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_261 = 7'h4 == index ? tag_1_4 : _GEN_260; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_262 = 7'h5 == index ? tag_1_5 : _GEN_261; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_263 = 7'h6 == index ? tag_1_6 : _GEN_262; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_264 = 7'h7 == index ? tag_1_7 : _GEN_263; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_265 = 7'h8 == index ? tag_1_8 : _GEN_264; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_266 = 7'h9 == index ? tag_1_9 : _GEN_265; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_267 = 7'ha == index ? tag_1_10 : _GEN_266; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_268 = 7'hb == index ? tag_1_11 : _GEN_267; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_269 = 7'hc == index ? tag_1_12 : _GEN_268; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_270 = 7'hd == index ? tag_1_13 : _GEN_269; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_271 = 7'he == index ? tag_1_14 : _GEN_270; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_272 = 7'hf == index ? tag_1_15 : _GEN_271; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_273 = 7'h10 == index ? tag_1_16 : _GEN_272; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_274 = 7'h11 == index ? tag_1_17 : _GEN_273; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_275 = 7'h12 == index ? tag_1_18 : _GEN_274; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_276 = 7'h13 == index ? tag_1_19 : _GEN_275; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_277 = 7'h14 == index ? tag_1_20 : _GEN_276; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_278 = 7'h15 == index ? tag_1_21 : _GEN_277; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_279 = 7'h16 == index ? tag_1_22 : _GEN_278; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_280 = 7'h17 == index ? tag_1_23 : _GEN_279; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_281 = 7'h18 == index ? tag_1_24 : _GEN_280; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_282 = 7'h19 == index ? tag_1_25 : _GEN_281; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_283 = 7'h1a == index ? tag_1_26 : _GEN_282; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_284 = 7'h1b == index ? tag_1_27 : _GEN_283; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_285 = 7'h1c == index ? tag_1_28 : _GEN_284; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_286 = 7'h1d == index ? tag_1_29 : _GEN_285; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_287 = 7'h1e == index ? tag_1_30 : _GEN_286; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_288 = 7'h1f == index ? tag_1_31 : _GEN_287; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_289 = 7'h20 == index ? tag_1_32 : _GEN_288; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_290 = 7'h21 == index ? tag_1_33 : _GEN_289; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_291 = 7'h22 == index ? tag_1_34 : _GEN_290; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_292 = 7'h23 == index ? tag_1_35 : _GEN_291; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_293 = 7'h24 == index ? tag_1_36 : _GEN_292; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_294 = 7'h25 == index ? tag_1_37 : _GEN_293; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_295 = 7'h26 == index ? tag_1_38 : _GEN_294; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_296 = 7'h27 == index ? tag_1_39 : _GEN_295; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_297 = 7'h28 == index ? tag_1_40 : _GEN_296; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_298 = 7'h29 == index ? tag_1_41 : _GEN_297; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_299 = 7'h2a == index ? tag_1_42 : _GEN_298; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_300 = 7'h2b == index ? tag_1_43 : _GEN_299; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_301 = 7'h2c == index ? tag_1_44 : _GEN_300; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_302 = 7'h2d == index ? tag_1_45 : _GEN_301; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_303 = 7'h2e == index ? tag_1_46 : _GEN_302; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_304 = 7'h2f == index ? tag_1_47 : _GEN_303; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_305 = 7'h30 == index ? tag_1_48 : _GEN_304; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_306 = 7'h31 == index ? tag_1_49 : _GEN_305; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_307 = 7'h32 == index ? tag_1_50 : _GEN_306; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_308 = 7'h33 == index ? tag_1_51 : _GEN_307; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_309 = 7'h34 == index ? tag_1_52 : _GEN_308; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_310 = 7'h35 == index ? tag_1_53 : _GEN_309; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_311 = 7'h36 == index ? tag_1_54 : _GEN_310; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_312 = 7'h37 == index ? tag_1_55 : _GEN_311; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_313 = 7'h38 == index ? tag_1_56 : _GEN_312; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_314 = 7'h39 == index ? tag_1_57 : _GEN_313; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_315 = 7'h3a == index ? tag_1_58 : _GEN_314; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_316 = 7'h3b == index ? tag_1_59 : _GEN_315; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_317 = 7'h3c == index ? tag_1_60 : _GEN_316; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_318 = 7'h3d == index ? tag_1_61 : _GEN_317; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_319 = 7'h3e == index ? tag_1_62 : _GEN_318; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_320 = 7'h3f == index ? tag_1_63 : _GEN_319; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_321 = 7'h40 == index ? tag_1_64 : _GEN_320; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_322 = 7'h41 == index ? tag_1_65 : _GEN_321; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_323 = 7'h42 == index ? tag_1_66 : _GEN_322; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_324 = 7'h43 == index ? tag_1_67 : _GEN_323; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_325 = 7'h44 == index ? tag_1_68 : _GEN_324; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_326 = 7'h45 == index ? tag_1_69 : _GEN_325; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_327 = 7'h46 == index ? tag_1_70 : _GEN_326; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_328 = 7'h47 == index ? tag_1_71 : _GEN_327; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_329 = 7'h48 == index ? tag_1_72 : _GEN_328; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_330 = 7'h49 == index ? tag_1_73 : _GEN_329; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_331 = 7'h4a == index ? tag_1_74 : _GEN_330; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_332 = 7'h4b == index ? tag_1_75 : _GEN_331; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_333 = 7'h4c == index ? tag_1_76 : _GEN_332; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_334 = 7'h4d == index ? tag_1_77 : _GEN_333; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_335 = 7'h4e == index ? tag_1_78 : _GEN_334; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_336 = 7'h4f == index ? tag_1_79 : _GEN_335; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_337 = 7'h50 == index ? tag_1_80 : _GEN_336; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_338 = 7'h51 == index ? tag_1_81 : _GEN_337; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_339 = 7'h52 == index ? tag_1_82 : _GEN_338; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_340 = 7'h53 == index ? tag_1_83 : _GEN_339; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_341 = 7'h54 == index ? tag_1_84 : _GEN_340; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_342 = 7'h55 == index ? tag_1_85 : _GEN_341; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_343 = 7'h56 == index ? tag_1_86 : _GEN_342; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_344 = 7'h57 == index ? tag_1_87 : _GEN_343; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_345 = 7'h58 == index ? tag_1_88 : _GEN_344; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_346 = 7'h59 == index ? tag_1_89 : _GEN_345; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_347 = 7'h5a == index ? tag_1_90 : _GEN_346; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_348 = 7'h5b == index ? tag_1_91 : _GEN_347; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_349 = 7'h5c == index ? tag_1_92 : _GEN_348; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_350 = 7'h5d == index ? tag_1_93 : _GEN_349; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_351 = 7'h5e == index ? tag_1_94 : _GEN_350; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_352 = 7'h5f == index ? tag_1_95 : _GEN_351; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_353 = 7'h60 == index ? tag_1_96 : _GEN_352; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_354 = 7'h61 == index ? tag_1_97 : _GEN_353; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_355 = 7'h62 == index ? tag_1_98 : _GEN_354; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_356 = 7'h63 == index ? tag_1_99 : _GEN_355; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_357 = 7'h64 == index ? tag_1_100 : _GEN_356; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_358 = 7'h65 == index ? tag_1_101 : _GEN_357; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_359 = 7'h66 == index ? tag_1_102 : _GEN_358; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_360 = 7'h67 == index ? tag_1_103 : _GEN_359; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_361 = 7'h68 == index ? tag_1_104 : _GEN_360; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_362 = 7'h69 == index ? tag_1_105 : _GEN_361; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_363 = 7'h6a == index ? tag_1_106 : _GEN_362; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_364 = 7'h6b == index ? tag_1_107 : _GEN_363; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_365 = 7'h6c == index ? tag_1_108 : _GEN_364; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_366 = 7'h6d == index ? tag_1_109 : _GEN_365; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_367 = 7'h6e == index ? tag_1_110 : _GEN_366; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_368 = 7'h6f == index ? tag_1_111 : _GEN_367; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_369 = 7'h70 == index ? tag_1_112 : _GEN_368; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_370 = 7'h71 == index ? tag_1_113 : _GEN_369; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_371 = 7'h72 == index ? tag_1_114 : _GEN_370; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_372 = 7'h73 == index ? tag_1_115 : _GEN_371; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_373 = 7'h74 == index ? tag_1_116 : _GEN_372; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_374 = 7'h75 == index ? tag_1_117 : _GEN_373; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_375 = 7'h76 == index ? tag_1_118 : _GEN_374; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_376 = 7'h77 == index ? tag_1_119 : _GEN_375; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_377 = 7'h78 == index ? tag_1_120 : _GEN_376; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_378 = 7'h79 == index ? tag_1_121 : _GEN_377; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_379 = 7'h7a == index ? tag_1_122 : _GEN_378; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_380 = 7'h7b == index ? tag_1_123 : _GEN_379; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_381 = 7'h7c == index ? tag_1_124 : _GEN_380; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_382 = 7'h7d == index ? tag_1_125 : _GEN_381; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_383 = 7'h7e == index ? tag_1_126 : _GEN_382; // @[d_cache.scala 68:{24,24}]
  wire [31:0] _GEN_384 = 7'h7f == index ? tag_1_127 : _GEN_383; // @[d_cache.scala 68:{24,24}]
  wire  _GEN_386 = 7'h1 == index ? valid_1_1 : valid_1_0; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_387 = 7'h2 == index ? valid_1_2 : _GEN_386; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_388 = 7'h3 == index ? valid_1_3 : _GEN_387; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_389 = 7'h4 == index ? valid_1_4 : _GEN_388; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_390 = 7'h5 == index ? valid_1_5 : _GEN_389; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_391 = 7'h6 == index ? valid_1_6 : _GEN_390; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_392 = 7'h7 == index ? valid_1_7 : _GEN_391; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_393 = 7'h8 == index ? valid_1_8 : _GEN_392; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_394 = 7'h9 == index ? valid_1_9 : _GEN_393; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_395 = 7'ha == index ? valid_1_10 : _GEN_394; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_396 = 7'hb == index ? valid_1_11 : _GEN_395; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_397 = 7'hc == index ? valid_1_12 : _GEN_396; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_398 = 7'hd == index ? valid_1_13 : _GEN_397; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_399 = 7'he == index ? valid_1_14 : _GEN_398; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_400 = 7'hf == index ? valid_1_15 : _GEN_399; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_401 = 7'h10 == index ? valid_1_16 : _GEN_400; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_402 = 7'h11 == index ? valid_1_17 : _GEN_401; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_403 = 7'h12 == index ? valid_1_18 : _GEN_402; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_404 = 7'h13 == index ? valid_1_19 : _GEN_403; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_405 = 7'h14 == index ? valid_1_20 : _GEN_404; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_406 = 7'h15 == index ? valid_1_21 : _GEN_405; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_407 = 7'h16 == index ? valid_1_22 : _GEN_406; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_408 = 7'h17 == index ? valid_1_23 : _GEN_407; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_409 = 7'h18 == index ? valid_1_24 : _GEN_408; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_410 = 7'h19 == index ? valid_1_25 : _GEN_409; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_411 = 7'h1a == index ? valid_1_26 : _GEN_410; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_412 = 7'h1b == index ? valid_1_27 : _GEN_411; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_413 = 7'h1c == index ? valid_1_28 : _GEN_412; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_414 = 7'h1d == index ? valid_1_29 : _GEN_413; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_415 = 7'h1e == index ? valid_1_30 : _GEN_414; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_416 = 7'h1f == index ? valid_1_31 : _GEN_415; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_417 = 7'h20 == index ? valid_1_32 : _GEN_416; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_418 = 7'h21 == index ? valid_1_33 : _GEN_417; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_419 = 7'h22 == index ? valid_1_34 : _GEN_418; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_420 = 7'h23 == index ? valid_1_35 : _GEN_419; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_421 = 7'h24 == index ? valid_1_36 : _GEN_420; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_422 = 7'h25 == index ? valid_1_37 : _GEN_421; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_423 = 7'h26 == index ? valid_1_38 : _GEN_422; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_424 = 7'h27 == index ? valid_1_39 : _GEN_423; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_425 = 7'h28 == index ? valid_1_40 : _GEN_424; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_426 = 7'h29 == index ? valid_1_41 : _GEN_425; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_427 = 7'h2a == index ? valid_1_42 : _GEN_426; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_428 = 7'h2b == index ? valid_1_43 : _GEN_427; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_429 = 7'h2c == index ? valid_1_44 : _GEN_428; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_430 = 7'h2d == index ? valid_1_45 : _GEN_429; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_431 = 7'h2e == index ? valid_1_46 : _GEN_430; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_432 = 7'h2f == index ? valid_1_47 : _GEN_431; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_433 = 7'h30 == index ? valid_1_48 : _GEN_432; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_434 = 7'h31 == index ? valid_1_49 : _GEN_433; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_435 = 7'h32 == index ? valid_1_50 : _GEN_434; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_436 = 7'h33 == index ? valid_1_51 : _GEN_435; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_437 = 7'h34 == index ? valid_1_52 : _GEN_436; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_438 = 7'h35 == index ? valid_1_53 : _GEN_437; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_439 = 7'h36 == index ? valid_1_54 : _GEN_438; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_440 = 7'h37 == index ? valid_1_55 : _GEN_439; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_441 = 7'h38 == index ? valid_1_56 : _GEN_440; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_442 = 7'h39 == index ? valid_1_57 : _GEN_441; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_443 = 7'h3a == index ? valid_1_58 : _GEN_442; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_444 = 7'h3b == index ? valid_1_59 : _GEN_443; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_445 = 7'h3c == index ? valid_1_60 : _GEN_444; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_446 = 7'h3d == index ? valid_1_61 : _GEN_445; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_447 = 7'h3e == index ? valid_1_62 : _GEN_446; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_448 = 7'h3f == index ? valid_1_63 : _GEN_447; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_449 = 7'h40 == index ? valid_1_64 : _GEN_448; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_450 = 7'h41 == index ? valid_1_65 : _GEN_449; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_451 = 7'h42 == index ? valid_1_66 : _GEN_450; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_452 = 7'h43 == index ? valid_1_67 : _GEN_451; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_453 = 7'h44 == index ? valid_1_68 : _GEN_452; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_454 = 7'h45 == index ? valid_1_69 : _GEN_453; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_455 = 7'h46 == index ? valid_1_70 : _GEN_454; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_456 = 7'h47 == index ? valid_1_71 : _GEN_455; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_457 = 7'h48 == index ? valid_1_72 : _GEN_456; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_458 = 7'h49 == index ? valid_1_73 : _GEN_457; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_459 = 7'h4a == index ? valid_1_74 : _GEN_458; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_460 = 7'h4b == index ? valid_1_75 : _GEN_459; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_461 = 7'h4c == index ? valid_1_76 : _GEN_460; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_462 = 7'h4d == index ? valid_1_77 : _GEN_461; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_463 = 7'h4e == index ? valid_1_78 : _GEN_462; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_464 = 7'h4f == index ? valid_1_79 : _GEN_463; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_465 = 7'h50 == index ? valid_1_80 : _GEN_464; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_466 = 7'h51 == index ? valid_1_81 : _GEN_465; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_467 = 7'h52 == index ? valid_1_82 : _GEN_466; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_468 = 7'h53 == index ? valid_1_83 : _GEN_467; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_469 = 7'h54 == index ? valid_1_84 : _GEN_468; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_470 = 7'h55 == index ? valid_1_85 : _GEN_469; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_471 = 7'h56 == index ? valid_1_86 : _GEN_470; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_472 = 7'h57 == index ? valid_1_87 : _GEN_471; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_473 = 7'h58 == index ? valid_1_88 : _GEN_472; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_474 = 7'h59 == index ? valid_1_89 : _GEN_473; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_475 = 7'h5a == index ? valid_1_90 : _GEN_474; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_476 = 7'h5b == index ? valid_1_91 : _GEN_475; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_477 = 7'h5c == index ? valid_1_92 : _GEN_476; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_478 = 7'h5d == index ? valid_1_93 : _GEN_477; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_479 = 7'h5e == index ? valid_1_94 : _GEN_478; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_480 = 7'h5f == index ? valid_1_95 : _GEN_479; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_481 = 7'h60 == index ? valid_1_96 : _GEN_480; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_482 = 7'h61 == index ? valid_1_97 : _GEN_481; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_483 = 7'h62 == index ? valid_1_98 : _GEN_482; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_484 = 7'h63 == index ? valid_1_99 : _GEN_483; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_485 = 7'h64 == index ? valid_1_100 : _GEN_484; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_486 = 7'h65 == index ? valid_1_101 : _GEN_485; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_487 = 7'h66 == index ? valid_1_102 : _GEN_486; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_488 = 7'h67 == index ? valid_1_103 : _GEN_487; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_489 = 7'h68 == index ? valid_1_104 : _GEN_488; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_490 = 7'h69 == index ? valid_1_105 : _GEN_489; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_491 = 7'h6a == index ? valid_1_106 : _GEN_490; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_492 = 7'h6b == index ? valid_1_107 : _GEN_491; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_493 = 7'h6c == index ? valid_1_108 : _GEN_492; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_494 = 7'h6d == index ? valid_1_109 : _GEN_493; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_495 = 7'h6e == index ? valid_1_110 : _GEN_494; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_496 = 7'h6f == index ? valid_1_111 : _GEN_495; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_497 = 7'h70 == index ? valid_1_112 : _GEN_496; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_498 = 7'h71 == index ? valid_1_113 : _GEN_497; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_499 = 7'h72 == index ? valid_1_114 : _GEN_498; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_500 = 7'h73 == index ? valid_1_115 : _GEN_499; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_501 = 7'h74 == index ? valid_1_116 : _GEN_500; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_502 = 7'h75 == index ? valid_1_117 : _GEN_501; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_503 = 7'h76 == index ? valid_1_118 : _GEN_502; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_504 = 7'h77 == index ? valid_1_119 : _GEN_503; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_505 = 7'h78 == index ? valid_1_120 : _GEN_504; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_506 = 7'h79 == index ? valid_1_121 : _GEN_505; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_507 = 7'h7a == index ? valid_1_122 : _GEN_506; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_508 = 7'h7b == index ? valid_1_123 : _GEN_507; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_509 = 7'h7c == index ? valid_1_124 : _GEN_508; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_510 = 7'h7d == index ? valid_1_125 : _GEN_509; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_511 = 7'h7e == index ? valid_1_126 : _GEN_510; // @[d_cache.scala 68:{50,50}]
  wire  _GEN_512 = 7'h7f == index ? valid_1_127 : _GEN_511; // @[d_cache.scala 68:{50,50}]
  wire  _T_7 = _GEN_384 == _GEN_19745 & _GEN_512; // @[d_cache.scala 68:33]
  reg [2:0] state; // @[d_cache.scala 82:24]
  wire  _T_14 = 3'h0 == state; // @[d_cache.scala 87:18]
  wire  _T_15 = 3'h1 == state; // @[d_cache.scala 87:18]
  wire  _GEN_519 = 7'h1 == index ? dirty_0_1 : dirty_0_0; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_520 = 7'h2 == index ? dirty_0_2 : _GEN_519; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_521 = 7'h3 == index ? dirty_0_3 : _GEN_520; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_522 = 7'h4 == index ? dirty_0_4 : _GEN_521; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_523 = 7'h5 == index ? dirty_0_5 : _GEN_522; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_524 = 7'h6 == index ? dirty_0_6 : _GEN_523; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_525 = 7'h7 == index ? dirty_0_7 : _GEN_524; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_526 = 7'h8 == index ? dirty_0_8 : _GEN_525; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_527 = 7'h9 == index ? dirty_0_9 : _GEN_526; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_528 = 7'ha == index ? dirty_0_10 : _GEN_527; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_529 = 7'hb == index ? dirty_0_11 : _GEN_528; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_530 = 7'hc == index ? dirty_0_12 : _GEN_529; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_531 = 7'hd == index ? dirty_0_13 : _GEN_530; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_532 = 7'he == index ? dirty_0_14 : _GEN_531; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_533 = 7'hf == index ? dirty_0_15 : _GEN_532; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_534 = 7'h10 == index ? dirty_0_16 : _GEN_533; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_535 = 7'h11 == index ? dirty_0_17 : _GEN_534; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_536 = 7'h12 == index ? dirty_0_18 : _GEN_535; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_537 = 7'h13 == index ? dirty_0_19 : _GEN_536; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_538 = 7'h14 == index ? dirty_0_20 : _GEN_537; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_539 = 7'h15 == index ? dirty_0_21 : _GEN_538; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_540 = 7'h16 == index ? dirty_0_22 : _GEN_539; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_541 = 7'h17 == index ? dirty_0_23 : _GEN_540; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_542 = 7'h18 == index ? dirty_0_24 : _GEN_541; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_543 = 7'h19 == index ? dirty_0_25 : _GEN_542; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_544 = 7'h1a == index ? dirty_0_26 : _GEN_543; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_545 = 7'h1b == index ? dirty_0_27 : _GEN_544; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_546 = 7'h1c == index ? dirty_0_28 : _GEN_545; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_547 = 7'h1d == index ? dirty_0_29 : _GEN_546; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_548 = 7'h1e == index ? dirty_0_30 : _GEN_547; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_549 = 7'h1f == index ? dirty_0_31 : _GEN_548; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_550 = 7'h20 == index ? dirty_0_32 : _GEN_549; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_551 = 7'h21 == index ? dirty_0_33 : _GEN_550; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_552 = 7'h22 == index ? dirty_0_34 : _GEN_551; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_553 = 7'h23 == index ? dirty_0_35 : _GEN_552; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_554 = 7'h24 == index ? dirty_0_36 : _GEN_553; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_555 = 7'h25 == index ? dirty_0_37 : _GEN_554; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_556 = 7'h26 == index ? dirty_0_38 : _GEN_555; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_557 = 7'h27 == index ? dirty_0_39 : _GEN_556; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_558 = 7'h28 == index ? dirty_0_40 : _GEN_557; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_559 = 7'h29 == index ? dirty_0_41 : _GEN_558; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_560 = 7'h2a == index ? dirty_0_42 : _GEN_559; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_561 = 7'h2b == index ? dirty_0_43 : _GEN_560; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_562 = 7'h2c == index ? dirty_0_44 : _GEN_561; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_563 = 7'h2d == index ? dirty_0_45 : _GEN_562; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_564 = 7'h2e == index ? dirty_0_46 : _GEN_563; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_565 = 7'h2f == index ? dirty_0_47 : _GEN_564; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_566 = 7'h30 == index ? dirty_0_48 : _GEN_565; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_567 = 7'h31 == index ? dirty_0_49 : _GEN_566; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_568 = 7'h32 == index ? dirty_0_50 : _GEN_567; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_569 = 7'h33 == index ? dirty_0_51 : _GEN_568; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_570 = 7'h34 == index ? dirty_0_52 : _GEN_569; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_571 = 7'h35 == index ? dirty_0_53 : _GEN_570; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_572 = 7'h36 == index ? dirty_0_54 : _GEN_571; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_573 = 7'h37 == index ? dirty_0_55 : _GEN_572; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_574 = 7'h38 == index ? dirty_0_56 : _GEN_573; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_575 = 7'h39 == index ? dirty_0_57 : _GEN_574; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_576 = 7'h3a == index ? dirty_0_58 : _GEN_575; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_577 = 7'h3b == index ? dirty_0_59 : _GEN_576; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_578 = 7'h3c == index ? dirty_0_60 : _GEN_577; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_579 = 7'h3d == index ? dirty_0_61 : _GEN_578; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_580 = 7'h3e == index ? dirty_0_62 : _GEN_579; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_581 = 7'h3f == index ? dirty_0_63 : _GEN_580; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_582 = 7'h40 == index ? dirty_0_64 : _GEN_581; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_583 = 7'h41 == index ? dirty_0_65 : _GEN_582; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_584 = 7'h42 == index ? dirty_0_66 : _GEN_583; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_585 = 7'h43 == index ? dirty_0_67 : _GEN_584; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_586 = 7'h44 == index ? dirty_0_68 : _GEN_585; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_587 = 7'h45 == index ? dirty_0_69 : _GEN_586; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_588 = 7'h46 == index ? dirty_0_70 : _GEN_587; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_589 = 7'h47 == index ? dirty_0_71 : _GEN_588; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_590 = 7'h48 == index ? dirty_0_72 : _GEN_589; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_591 = 7'h49 == index ? dirty_0_73 : _GEN_590; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_592 = 7'h4a == index ? dirty_0_74 : _GEN_591; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_593 = 7'h4b == index ? dirty_0_75 : _GEN_592; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_594 = 7'h4c == index ? dirty_0_76 : _GEN_593; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_595 = 7'h4d == index ? dirty_0_77 : _GEN_594; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_596 = 7'h4e == index ? dirty_0_78 : _GEN_595; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_597 = 7'h4f == index ? dirty_0_79 : _GEN_596; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_598 = 7'h50 == index ? dirty_0_80 : _GEN_597; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_599 = 7'h51 == index ? dirty_0_81 : _GEN_598; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_600 = 7'h52 == index ? dirty_0_82 : _GEN_599; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_601 = 7'h53 == index ? dirty_0_83 : _GEN_600; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_602 = 7'h54 == index ? dirty_0_84 : _GEN_601; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_603 = 7'h55 == index ? dirty_0_85 : _GEN_602; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_604 = 7'h56 == index ? dirty_0_86 : _GEN_603; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_605 = 7'h57 == index ? dirty_0_87 : _GEN_604; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_606 = 7'h58 == index ? dirty_0_88 : _GEN_605; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_607 = 7'h59 == index ? dirty_0_89 : _GEN_606; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_608 = 7'h5a == index ? dirty_0_90 : _GEN_607; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_609 = 7'h5b == index ? dirty_0_91 : _GEN_608; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_610 = 7'h5c == index ? dirty_0_92 : _GEN_609; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_611 = 7'h5d == index ? dirty_0_93 : _GEN_610; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_612 = 7'h5e == index ? dirty_0_94 : _GEN_611; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_613 = 7'h5f == index ? dirty_0_95 : _GEN_612; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_614 = 7'h60 == index ? dirty_0_96 : _GEN_613; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_615 = 7'h61 == index ? dirty_0_97 : _GEN_614; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_616 = 7'h62 == index ? dirty_0_98 : _GEN_615; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_617 = 7'h63 == index ? dirty_0_99 : _GEN_616; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_618 = 7'h64 == index ? dirty_0_100 : _GEN_617; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_619 = 7'h65 == index ? dirty_0_101 : _GEN_618; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_620 = 7'h66 == index ? dirty_0_102 : _GEN_619; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_621 = 7'h67 == index ? dirty_0_103 : _GEN_620; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_622 = 7'h68 == index ? dirty_0_104 : _GEN_621; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_623 = 7'h69 == index ? dirty_0_105 : _GEN_622; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_624 = 7'h6a == index ? dirty_0_106 : _GEN_623; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_625 = 7'h6b == index ? dirty_0_107 : _GEN_624; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_626 = 7'h6c == index ? dirty_0_108 : _GEN_625; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_627 = 7'h6d == index ? dirty_0_109 : _GEN_626; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_628 = 7'h6e == index ? dirty_0_110 : _GEN_627; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_629 = 7'h6f == index ? dirty_0_111 : _GEN_628; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_630 = 7'h70 == index ? dirty_0_112 : _GEN_629; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_631 = 7'h71 == index ? dirty_0_113 : _GEN_630; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_632 = 7'h72 == index ? dirty_0_114 : _GEN_631; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_633 = 7'h73 == index ? dirty_0_115 : _GEN_632; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_634 = 7'h74 == index ? dirty_0_116 : _GEN_633; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_635 = 7'h75 == index ? dirty_0_117 : _GEN_634; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_636 = 7'h76 == index ? dirty_0_118 : _GEN_635; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_637 = 7'h77 == index ? dirty_0_119 : _GEN_636; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_638 = 7'h78 == index ? dirty_0_120 : _GEN_637; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_639 = 7'h79 == index ? dirty_0_121 : _GEN_638; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_640 = 7'h7a == index ? dirty_0_122 : _GEN_639; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_641 = 7'h7b == index ? dirty_0_123 : _GEN_640; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_642 = 7'h7c == index ? dirty_0_124 : _GEN_641; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_643 = 7'h7d == index ? dirty_0_125 : _GEN_642; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_644 = 7'h7e == index ? dirty_0_126 : _GEN_643; // @[d_cache.scala 99:{27,27}]
  wire  _GEN_645 = 7'h7f == index ? dirty_0_127 : _GEN_644; // @[d_cache.scala 99:{27,27}]
  wire [2:0] _GEN_646 = io_from_lsu_rready ? 3'h0 : state; // @[d_cache.scala 100:27 82:24 98:41]
  wire  _GEN_648 = 7'h1 == index ? dirty_1_1 : dirty_1_0; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_649 = 7'h2 == index ? dirty_1_2 : _GEN_648; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_650 = 7'h3 == index ? dirty_1_3 : _GEN_649; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_651 = 7'h4 == index ? dirty_1_4 : _GEN_650; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_652 = 7'h5 == index ? dirty_1_5 : _GEN_651; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_653 = 7'h6 == index ? dirty_1_6 : _GEN_652; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_654 = 7'h7 == index ? dirty_1_7 : _GEN_653; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_655 = 7'h8 == index ? dirty_1_8 : _GEN_654; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_656 = 7'h9 == index ? dirty_1_9 : _GEN_655; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_657 = 7'ha == index ? dirty_1_10 : _GEN_656; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_658 = 7'hb == index ? dirty_1_11 : _GEN_657; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_659 = 7'hc == index ? dirty_1_12 : _GEN_658; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_660 = 7'hd == index ? dirty_1_13 : _GEN_659; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_661 = 7'he == index ? dirty_1_14 : _GEN_660; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_662 = 7'hf == index ? dirty_1_15 : _GEN_661; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_663 = 7'h10 == index ? dirty_1_16 : _GEN_662; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_664 = 7'h11 == index ? dirty_1_17 : _GEN_663; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_665 = 7'h12 == index ? dirty_1_18 : _GEN_664; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_666 = 7'h13 == index ? dirty_1_19 : _GEN_665; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_667 = 7'h14 == index ? dirty_1_20 : _GEN_666; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_668 = 7'h15 == index ? dirty_1_21 : _GEN_667; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_669 = 7'h16 == index ? dirty_1_22 : _GEN_668; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_670 = 7'h17 == index ? dirty_1_23 : _GEN_669; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_671 = 7'h18 == index ? dirty_1_24 : _GEN_670; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_672 = 7'h19 == index ? dirty_1_25 : _GEN_671; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_673 = 7'h1a == index ? dirty_1_26 : _GEN_672; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_674 = 7'h1b == index ? dirty_1_27 : _GEN_673; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_675 = 7'h1c == index ? dirty_1_28 : _GEN_674; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_676 = 7'h1d == index ? dirty_1_29 : _GEN_675; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_677 = 7'h1e == index ? dirty_1_30 : _GEN_676; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_678 = 7'h1f == index ? dirty_1_31 : _GEN_677; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_679 = 7'h20 == index ? dirty_1_32 : _GEN_678; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_680 = 7'h21 == index ? dirty_1_33 : _GEN_679; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_681 = 7'h22 == index ? dirty_1_34 : _GEN_680; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_682 = 7'h23 == index ? dirty_1_35 : _GEN_681; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_683 = 7'h24 == index ? dirty_1_36 : _GEN_682; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_684 = 7'h25 == index ? dirty_1_37 : _GEN_683; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_685 = 7'h26 == index ? dirty_1_38 : _GEN_684; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_686 = 7'h27 == index ? dirty_1_39 : _GEN_685; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_687 = 7'h28 == index ? dirty_1_40 : _GEN_686; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_688 = 7'h29 == index ? dirty_1_41 : _GEN_687; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_689 = 7'h2a == index ? dirty_1_42 : _GEN_688; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_690 = 7'h2b == index ? dirty_1_43 : _GEN_689; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_691 = 7'h2c == index ? dirty_1_44 : _GEN_690; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_692 = 7'h2d == index ? dirty_1_45 : _GEN_691; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_693 = 7'h2e == index ? dirty_1_46 : _GEN_692; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_694 = 7'h2f == index ? dirty_1_47 : _GEN_693; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_695 = 7'h30 == index ? dirty_1_48 : _GEN_694; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_696 = 7'h31 == index ? dirty_1_49 : _GEN_695; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_697 = 7'h32 == index ? dirty_1_50 : _GEN_696; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_698 = 7'h33 == index ? dirty_1_51 : _GEN_697; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_699 = 7'h34 == index ? dirty_1_52 : _GEN_698; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_700 = 7'h35 == index ? dirty_1_53 : _GEN_699; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_701 = 7'h36 == index ? dirty_1_54 : _GEN_700; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_702 = 7'h37 == index ? dirty_1_55 : _GEN_701; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_703 = 7'h38 == index ? dirty_1_56 : _GEN_702; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_704 = 7'h39 == index ? dirty_1_57 : _GEN_703; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_705 = 7'h3a == index ? dirty_1_58 : _GEN_704; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_706 = 7'h3b == index ? dirty_1_59 : _GEN_705; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_707 = 7'h3c == index ? dirty_1_60 : _GEN_706; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_708 = 7'h3d == index ? dirty_1_61 : _GEN_707; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_709 = 7'h3e == index ? dirty_1_62 : _GEN_708; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_710 = 7'h3f == index ? dirty_1_63 : _GEN_709; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_711 = 7'h40 == index ? dirty_1_64 : _GEN_710; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_712 = 7'h41 == index ? dirty_1_65 : _GEN_711; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_713 = 7'h42 == index ? dirty_1_66 : _GEN_712; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_714 = 7'h43 == index ? dirty_1_67 : _GEN_713; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_715 = 7'h44 == index ? dirty_1_68 : _GEN_714; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_716 = 7'h45 == index ? dirty_1_69 : _GEN_715; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_717 = 7'h46 == index ? dirty_1_70 : _GEN_716; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_718 = 7'h47 == index ? dirty_1_71 : _GEN_717; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_719 = 7'h48 == index ? dirty_1_72 : _GEN_718; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_720 = 7'h49 == index ? dirty_1_73 : _GEN_719; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_721 = 7'h4a == index ? dirty_1_74 : _GEN_720; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_722 = 7'h4b == index ? dirty_1_75 : _GEN_721; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_723 = 7'h4c == index ? dirty_1_76 : _GEN_722; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_724 = 7'h4d == index ? dirty_1_77 : _GEN_723; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_725 = 7'h4e == index ? dirty_1_78 : _GEN_724; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_726 = 7'h4f == index ? dirty_1_79 : _GEN_725; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_727 = 7'h50 == index ? dirty_1_80 : _GEN_726; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_728 = 7'h51 == index ? dirty_1_81 : _GEN_727; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_729 = 7'h52 == index ? dirty_1_82 : _GEN_728; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_730 = 7'h53 == index ? dirty_1_83 : _GEN_729; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_731 = 7'h54 == index ? dirty_1_84 : _GEN_730; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_732 = 7'h55 == index ? dirty_1_85 : _GEN_731; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_733 = 7'h56 == index ? dirty_1_86 : _GEN_732; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_734 = 7'h57 == index ? dirty_1_87 : _GEN_733; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_735 = 7'h58 == index ? dirty_1_88 : _GEN_734; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_736 = 7'h59 == index ? dirty_1_89 : _GEN_735; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_737 = 7'h5a == index ? dirty_1_90 : _GEN_736; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_738 = 7'h5b == index ? dirty_1_91 : _GEN_737; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_739 = 7'h5c == index ? dirty_1_92 : _GEN_738; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_740 = 7'h5d == index ? dirty_1_93 : _GEN_739; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_741 = 7'h5e == index ? dirty_1_94 : _GEN_740; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_742 = 7'h5f == index ? dirty_1_95 : _GEN_741; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_743 = 7'h60 == index ? dirty_1_96 : _GEN_742; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_744 = 7'h61 == index ? dirty_1_97 : _GEN_743; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_745 = 7'h62 == index ? dirty_1_98 : _GEN_744; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_746 = 7'h63 == index ? dirty_1_99 : _GEN_745; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_747 = 7'h64 == index ? dirty_1_100 : _GEN_746; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_748 = 7'h65 == index ? dirty_1_101 : _GEN_747; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_749 = 7'h66 == index ? dirty_1_102 : _GEN_748; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_750 = 7'h67 == index ? dirty_1_103 : _GEN_749; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_751 = 7'h68 == index ? dirty_1_104 : _GEN_750; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_752 = 7'h69 == index ? dirty_1_105 : _GEN_751; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_753 = 7'h6a == index ? dirty_1_106 : _GEN_752; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_754 = 7'h6b == index ? dirty_1_107 : _GEN_753; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_755 = 7'h6c == index ? dirty_1_108 : _GEN_754; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_756 = 7'h6d == index ? dirty_1_109 : _GEN_755; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_757 = 7'h6e == index ? dirty_1_110 : _GEN_756; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_758 = 7'h6f == index ? dirty_1_111 : _GEN_757; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_759 = 7'h70 == index ? dirty_1_112 : _GEN_758; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_760 = 7'h71 == index ? dirty_1_113 : _GEN_759; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_761 = 7'h72 == index ? dirty_1_114 : _GEN_760; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_762 = 7'h73 == index ? dirty_1_115 : _GEN_761; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_763 = 7'h74 == index ? dirty_1_116 : _GEN_762; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_764 = 7'h75 == index ? dirty_1_117 : _GEN_763; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_765 = 7'h76 == index ? dirty_1_118 : _GEN_764; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_766 = 7'h77 == index ? dirty_1_119 : _GEN_765; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_767 = 7'h78 == index ? dirty_1_120 : _GEN_766; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_768 = 7'h79 == index ? dirty_1_121 : _GEN_767; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_769 = 7'h7a == index ? dirty_1_122 : _GEN_768; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_770 = 7'h7b == index ? dirty_1_123 : _GEN_769; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_771 = 7'h7c == index ? dirty_1_124 : _GEN_770; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_772 = 7'h7d == index ? dirty_1_125 : _GEN_771; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_773 = 7'h7e == index ? dirty_1_126 : _GEN_772; // @[d_cache.scala 105:{27,27}]
  wire  _GEN_774 = 7'h7f == index ? dirty_1_127 : _GEN_773; // @[d_cache.scala 105:{27,27}]
  wire [2:0] _GEN_775 = way1_hit ? _GEN_646 : 3'h3; // @[d_cache.scala 103:33 109:23]
  wire [63:0] _ram_0_T = io_from_lsu_wdata & wmask; // @[d_cache.scala 115:53]
  wire [126:0] _GEN_20785 = {{63'd0}, _ram_0_T}; // @[d_cache.scala 115:62]
  wire [126:0] _ram_0_T_1 = _GEN_20785 << shift_bit; // @[d_cache.scala 115:62]
  wire [126:0] _GEN_20786 = {{63'd0}, wmask}; // @[d_cache.scala 115:102]
  wire [126:0] _ram_0_T_2 = _GEN_20786 << shift_bit; // @[d_cache.scala 115:102]
  wire [126:0] _ram_0_T_3 = ~_ram_0_T_2; // @[d_cache.scala 115:94]
  wire [63:0] _GEN_778 = 7'h1 == index ? ram_0_1 : ram_0_0; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_779 = 7'h2 == index ? ram_0_2 : _GEN_778; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_780 = 7'h3 == index ? ram_0_3 : _GEN_779; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_781 = 7'h4 == index ? ram_0_4 : _GEN_780; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_782 = 7'h5 == index ? ram_0_5 : _GEN_781; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_783 = 7'h6 == index ? ram_0_6 : _GEN_782; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_784 = 7'h7 == index ? ram_0_7 : _GEN_783; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_785 = 7'h8 == index ? ram_0_8 : _GEN_784; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_786 = 7'h9 == index ? ram_0_9 : _GEN_785; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_787 = 7'ha == index ? ram_0_10 : _GEN_786; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_788 = 7'hb == index ? ram_0_11 : _GEN_787; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_789 = 7'hc == index ? ram_0_12 : _GEN_788; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_790 = 7'hd == index ? ram_0_13 : _GEN_789; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_791 = 7'he == index ? ram_0_14 : _GEN_790; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_792 = 7'hf == index ? ram_0_15 : _GEN_791; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_793 = 7'h10 == index ? ram_0_16 : _GEN_792; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_794 = 7'h11 == index ? ram_0_17 : _GEN_793; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_795 = 7'h12 == index ? ram_0_18 : _GEN_794; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_796 = 7'h13 == index ? ram_0_19 : _GEN_795; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_797 = 7'h14 == index ? ram_0_20 : _GEN_796; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_798 = 7'h15 == index ? ram_0_21 : _GEN_797; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_799 = 7'h16 == index ? ram_0_22 : _GEN_798; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_800 = 7'h17 == index ? ram_0_23 : _GEN_799; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_801 = 7'h18 == index ? ram_0_24 : _GEN_800; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_802 = 7'h19 == index ? ram_0_25 : _GEN_801; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_803 = 7'h1a == index ? ram_0_26 : _GEN_802; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_804 = 7'h1b == index ? ram_0_27 : _GEN_803; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_805 = 7'h1c == index ? ram_0_28 : _GEN_804; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_806 = 7'h1d == index ? ram_0_29 : _GEN_805; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_807 = 7'h1e == index ? ram_0_30 : _GEN_806; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_808 = 7'h1f == index ? ram_0_31 : _GEN_807; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_809 = 7'h20 == index ? ram_0_32 : _GEN_808; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_810 = 7'h21 == index ? ram_0_33 : _GEN_809; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_811 = 7'h22 == index ? ram_0_34 : _GEN_810; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_812 = 7'h23 == index ? ram_0_35 : _GEN_811; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_813 = 7'h24 == index ? ram_0_36 : _GEN_812; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_814 = 7'h25 == index ? ram_0_37 : _GEN_813; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_815 = 7'h26 == index ? ram_0_38 : _GEN_814; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_816 = 7'h27 == index ? ram_0_39 : _GEN_815; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_817 = 7'h28 == index ? ram_0_40 : _GEN_816; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_818 = 7'h29 == index ? ram_0_41 : _GEN_817; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_819 = 7'h2a == index ? ram_0_42 : _GEN_818; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_820 = 7'h2b == index ? ram_0_43 : _GEN_819; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_821 = 7'h2c == index ? ram_0_44 : _GEN_820; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_822 = 7'h2d == index ? ram_0_45 : _GEN_821; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_823 = 7'h2e == index ? ram_0_46 : _GEN_822; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_824 = 7'h2f == index ? ram_0_47 : _GEN_823; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_825 = 7'h30 == index ? ram_0_48 : _GEN_824; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_826 = 7'h31 == index ? ram_0_49 : _GEN_825; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_827 = 7'h32 == index ? ram_0_50 : _GEN_826; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_828 = 7'h33 == index ? ram_0_51 : _GEN_827; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_829 = 7'h34 == index ? ram_0_52 : _GEN_828; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_830 = 7'h35 == index ? ram_0_53 : _GEN_829; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_831 = 7'h36 == index ? ram_0_54 : _GEN_830; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_832 = 7'h37 == index ? ram_0_55 : _GEN_831; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_833 = 7'h38 == index ? ram_0_56 : _GEN_832; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_834 = 7'h39 == index ? ram_0_57 : _GEN_833; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_835 = 7'h3a == index ? ram_0_58 : _GEN_834; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_836 = 7'h3b == index ? ram_0_59 : _GEN_835; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_837 = 7'h3c == index ? ram_0_60 : _GEN_836; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_838 = 7'h3d == index ? ram_0_61 : _GEN_837; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_839 = 7'h3e == index ? ram_0_62 : _GEN_838; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_840 = 7'h3f == index ? ram_0_63 : _GEN_839; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_841 = 7'h40 == index ? ram_0_64 : _GEN_840; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_842 = 7'h41 == index ? ram_0_65 : _GEN_841; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_843 = 7'h42 == index ? ram_0_66 : _GEN_842; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_844 = 7'h43 == index ? ram_0_67 : _GEN_843; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_845 = 7'h44 == index ? ram_0_68 : _GEN_844; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_846 = 7'h45 == index ? ram_0_69 : _GEN_845; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_847 = 7'h46 == index ? ram_0_70 : _GEN_846; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_848 = 7'h47 == index ? ram_0_71 : _GEN_847; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_849 = 7'h48 == index ? ram_0_72 : _GEN_848; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_850 = 7'h49 == index ? ram_0_73 : _GEN_849; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_851 = 7'h4a == index ? ram_0_74 : _GEN_850; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_852 = 7'h4b == index ? ram_0_75 : _GEN_851; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_853 = 7'h4c == index ? ram_0_76 : _GEN_852; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_854 = 7'h4d == index ? ram_0_77 : _GEN_853; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_855 = 7'h4e == index ? ram_0_78 : _GEN_854; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_856 = 7'h4f == index ? ram_0_79 : _GEN_855; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_857 = 7'h50 == index ? ram_0_80 : _GEN_856; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_858 = 7'h51 == index ? ram_0_81 : _GEN_857; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_859 = 7'h52 == index ? ram_0_82 : _GEN_858; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_860 = 7'h53 == index ? ram_0_83 : _GEN_859; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_861 = 7'h54 == index ? ram_0_84 : _GEN_860; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_862 = 7'h55 == index ? ram_0_85 : _GEN_861; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_863 = 7'h56 == index ? ram_0_86 : _GEN_862; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_864 = 7'h57 == index ? ram_0_87 : _GEN_863; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_865 = 7'h58 == index ? ram_0_88 : _GEN_864; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_866 = 7'h59 == index ? ram_0_89 : _GEN_865; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_867 = 7'h5a == index ? ram_0_90 : _GEN_866; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_868 = 7'h5b == index ? ram_0_91 : _GEN_867; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_869 = 7'h5c == index ? ram_0_92 : _GEN_868; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_870 = 7'h5d == index ? ram_0_93 : _GEN_869; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_871 = 7'h5e == index ? ram_0_94 : _GEN_870; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_872 = 7'h5f == index ? ram_0_95 : _GEN_871; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_873 = 7'h60 == index ? ram_0_96 : _GEN_872; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_874 = 7'h61 == index ? ram_0_97 : _GEN_873; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_875 = 7'h62 == index ? ram_0_98 : _GEN_874; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_876 = 7'h63 == index ? ram_0_99 : _GEN_875; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_877 = 7'h64 == index ? ram_0_100 : _GEN_876; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_878 = 7'h65 == index ? ram_0_101 : _GEN_877; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_879 = 7'h66 == index ? ram_0_102 : _GEN_878; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_880 = 7'h67 == index ? ram_0_103 : _GEN_879; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_881 = 7'h68 == index ? ram_0_104 : _GEN_880; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_882 = 7'h69 == index ? ram_0_105 : _GEN_881; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_883 = 7'h6a == index ? ram_0_106 : _GEN_882; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_884 = 7'h6b == index ? ram_0_107 : _GEN_883; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_885 = 7'h6c == index ? ram_0_108 : _GEN_884; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_886 = 7'h6d == index ? ram_0_109 : _GEN_885; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_887 = 7'h6e == index ? ram_0_110 : _GEN_886; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_888 = 7'h6f == index ? ram_0_111 : _GEN_887; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_889 = 7'h70 == index ? ram_0_112 : _GEN_888; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_890 = 7'h71 == index ? ram_0_113 : _GEN_889; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_891 = 7'h72 == index ? ram_0_114 : _GEN_890; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_892 = 7'h73 == index ? ram_0_115 : _GEN_891; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_893 = 7'h74 == index ? ram_0_116 : _GEN_892; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_894 = 7'h75 == index ? ram_0_117 : _GEN_893; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_895 = 7'h76 == index ? ram_0_118 : _GEN_894; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_896 = 7'h77 == index ? ram_0_119 : _GEN_895; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_897 = 7'h78 == index ? ram_0_120 : _GEN_896; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_898 = 7'h79 == index ? ram_0_121 : _GEN_897; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_899 = 7'h7a == index ? ram_0_122 : _GEN_898; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_900 = 7'h7b == index ? ram_0_123 : _GEN_899; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_901 = 7'h7c == index ? ram_0_124 : _GEN_900; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_902 = 7'h7d == index ? ram_0_125 : _GEN_901; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_903 = 7'h7e == index ? ram_0_126 : _GEN_902; // @[d_cache.scala 115:{92,92}]
  wire [63:0] _GEN_904 = 7'h7f == index ? ram_0_127 : _GEN_903; // @[d_cache.scala 115:{92,92}]
  wire [126:0] _GEN_19747 = {{63'd0}, _GEN_904}; // @[d_cache.scala 115:92]
  wire [126:0] _ram_0_T_4 = _GEN_19747 & _ram_0_T_3; // @[d_cache.scala 115:92]
  wire [126:0] _ram_0_T_5 = _ram_0_T_1 | _ram_0_T_4; // @[d_cache.scala 115:76]
  wire [63:0] _GEN_905 = 7'h0 == index ? _ram_0_T_5[63:0] : ram_0_0; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_906 = 7'h1 == index ? _ram_0_T_5[63:0] : ram_0_1; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_907 = 7'h2 == index ? _ram_0_T_5[63:0] : ram_0_2; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_908 = 7'h3 == index ? _ram_0_T_5[63:0] : ram_0_3; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_909 = 7'h4 == index ? _ram_0_T_5[63:0] : ram_0_4; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_910 = 7'h5 == index ? _ram_0_T_5[63:0] : ram_0_5; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_911 = 7'h6 == index ? _ram_0_T_5[63:0] : ram_0_6; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_912 = 7'h7 == index ? _ram_0_T_5[63:0] : ram_0_7; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_913 = 7'h8 == index ? _ram_0_T_5[63:0] : ram_0_8; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_914 = 7'h9 == index ? _ram_0_T_5[63:0] : ram_0_9; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_915 = 7'ha == index ? _ram_0_T_5[63:0] : ram_0_10; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_916 = 7'hb == index ? _ram_0_T_5[63:0] : ram_0_11; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_917 = 7'hc == index ? _ram_0_T_5[63:0] : ram_0_12; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_918 = 7'hd == index ? _ram_0_T_5[63:0] : ram_0_13; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_919 = 7'he == index ? _ram_0_T_5[63:0] : ram_0_14; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_920 = 7'hf == index ? _ram_0_T_5[63:0] : ram_0_15; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_921 = 7'h10 == index ? _ram_0_T_5[63:0] : ram_0_16; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_922 = 7'h11 == index ? _ram_0_T_5[63:0] : ram_0_17; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_923 = 7'h12 == index ? _ram_0_T_5[63:0] : ram_0_18; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_924 = 7'h13 == index ? _ram_0_T_5[63:0] : ram_0_19; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_925 = 7'h14 == index ? _ram_0_T_5[63:0] : ram_0_20; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_926 = 7'h15 == index ? _ram_0_T_5[63:0] : ram_0_21; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_927 = 7'h16 == index ? _ram_0_T_5[63:0] : ram_0_22; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_928 = 7'h17 == index ? _ram_0_T_5[63:0] : ram_0_23; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_929 = 7'h18 == index ? _ram_0_T_5[63:0] : ram_0_24; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_930 = 7'h19 == index ? _ram_0_T_5[63:0] : ram_0_25; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_931 = 7'h1a == index ? _ram_0_T_5[63:0] : ram_0_26; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_932 = 7'h1b == index ? _ram_0_T_5[63:0] : ram_0_27; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_933 = 7'h1c == index ? _ram_0_T_5[63:0] : ram_0_28; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_934 = 7'h1d == index ? _ram_0_T_5[63:0] : ram_0_29; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_935 = 7'h1e == index ? _ram_0_T_5[63:0] : ram_0_30; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_936 = 7'h1f == index ? _ram_0_T_5[63:0] : ram_0_31; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_937 = 7'h20 == index ? _ram_0_T_5[63:0] : ram_0_32; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_938 = 7'h21 == index ? _ram_0_T_5[63:0] : ram_0_33; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_939 = 7'h22 == index ? _ram_0_T_5[63:0] : ram_0_34; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_940 = 7'h23 == index ? _ram_0_T_5[63:0] : ram_0_35; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_941 = 7'h24 == index ? _ram_0_T_5[63:0] : ram_0_36; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_942 = 7'h25 == index ? _ram_0_T_5[63:0] : ram_0_37; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_943 = 7'h26 == index ? _ram_0_T_5[63:0] : ram_0_38; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_944 = 7'h27 == index ? _ram_0_T_5[63:0] : ram_0_39; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_945 = 7'h28 == index ? _ram_0_T_5[63:0] : ram_0_40; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_946 = 7'h29 == index ? _ram_0_T_5[63:0] : ram_0_41; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_947 = 7'h2a == index ? _ram_0_T_5[63:0] : ram_0_42; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_948 = 7'h2b == index ? _ram_0_T_5[63:0] : ram_0_43; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_949 = 7'h2c == index ? _ram_0_T_5[63:0] : ram_0_44; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_950 = 7'h2d == index ? _ram_0_T_5[63:0] : ram_0_45; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_951 = 7'h2e == index ? _ram_0_T_5[63:0] : ram_0_46; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_952 = 7'h2f == index ? _ram_0_T_5[63:0] : ram_0_47; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_953 = 7'h30 == index ? _ram_0_T_5[63:0] : ram_0_48; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_954 = 7'h31 == index ? _ram_0_T_5[63:0] : ram_0_49; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_955 = 7'h32 == index ? _ram_0_T_5[63:0] : ram_0_50; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_956 = 7'h33 == index ? _ram_0_T_5[63:0] : ram_0_51; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_957 = 7'h34 == index ? _ram_0_T_5[63:0] : ram_0_52; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_958 = 7'h35 == index ? _ram_0_T_5[63:0] : ram_0_53; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_959 = 7'h36 == index ? _ram_0_T_5[63:0] : ram_0_54; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_960 = 7'h37 == index ? _ram_0_T_5[63:0] : ram_0_55; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_961 = 7'h38 == index ? _ram_0_T_5[63:0] : ram_0_56; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_962 = 7'h39 == index ? _ram_0_T_5[63:0] : ram_0_57; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_963 = 7'h3a == index ? _ram_0_T_5[63:0] : ram_0_58; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_964 = 7'h3b == index ? _ram_0_T_5[63:0] : ram_0_59; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_965 = 7'h3c == index ? _ram_0_T_5[63:0] : ram_0_60; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_966 = 7'h3d == index ? _ram_0_T_5[63:0] : ram_0_61; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_967 = 7'h3e == index ? _ram_0_T_5[63:0] : ram_0_62; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_968 = 7'h3f == index ? _ram_0_T_5[63:0] : ram_0_63; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_969 = 7'h40 == index ? _ram_0_T_5[63:0] : ram_0_64; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_970 = 7'h41 == index ? _ram_0_T_5[63:0] : ram_0_65; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_971 = 7'h42 == index ? _ram_0_T_5[63:0] : ram_0_66; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_972 = 7'h43 == index ? _ram_0_T_5[63:0] : ram_0_67; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_973 = 7'h44 == index ? _ram_0_T_5[63:0] : ram_0_68; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_974 = 7'h45 == index ? _ram_0_T_5[63:0] : ram_0_69; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_975 = 7'h46 == index ? _ram_0_T_5[63:0] : ram_0_70; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_976 = 7'h47 == index ? _ram_0_T_5[63:0] : ram_0_71; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_977 = 7'h48 == index ? _ram_0_T_5[63:0] : ram_0_72; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_978 = 7'h49 == index ? _ram_0_T_5[63:0] : ram_0_73; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_979 = 7'h4a == index ? _ram_0_T_5[63:0] : ram_0_74; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_980 = 7'h4b == index ? _ram_0_T_5[63:0] : ram_0_75; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_981 = 7'h4c == index ? _ram_0_T_5[63:0] : ram_0_76; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_982 = 7'h4d == index ? _ram_0_T_5[63:0] : ram_0_77; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_983 = 7'h4e == index ? _ram_0_T_5[63:0] : ram_0_78; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_984 = 7'h4f == index ? _ram_0_T_5[63:0] : ram_0_79; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_985 = 7'h50 == index ? _ram_0_T_5[63:0] : ram_0_80; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_986 = 7'h51 == index ? _ram_0_T_5[63:0] : ram_0_81; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_987 = 7'h52 == index ? _ram_0_T_5[63:0] : ram_0_82; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_988 = 7'h53 == index ? _ram_0_T_5[63:0] : ram_0_83; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_989 = 7'h54 == index ? _ram_0_T_5[63:0] : ram_0_84; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_990 = 7'h55 == index ? _ram_0_T_5[63:0] : ram_0_85; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_991 = 7'h56 == index ? _ram_0_T_5[63:0] : ram_0_86; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_992 = 7'h57 == index ? _ram_0_T_5[63:0] : ram_0_87; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_993 = 7'h58 == index ? _ram_0_T_5[63:0] : ram_0_88; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_994 = 7'h59 == index ? _ram_0_T_5[63:0] : ram_0_89; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_995 = 7'h5a == index ? _ram_0_T_5[63:0] : ram_0_90; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_996 = 7'h5b == index ? _ram_0_T_5[63:0] : ram_0_91; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_997 = 7'h5c == index ? _ram_0_T_5[63:0] : ram_0_92; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_998 = 7'h5d == index ? _ram_0_T_5[63:0] : ram_0_93; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_999 = 7'h5e == index ? _ram_0_T_5[63:0] : ram_0_94; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1000 = 7'h5f == index ? _ram_0_T_5[63:0] : ram_0_95; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1001 = 7'h60 == index ? _ram_0_T_5[63:0] : ram_0_96; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1002 = 7'h61 == index ? _ram_0_T_5[63:0] : ram_0_97; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1003 = 7'h62 == index ? _ram_0_T_5[63:0] : ram_0_98; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1004 = 7'h63 == index ? _ram_0_T_5[63:0] : ram_0_99; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1005 = 7'h64 == index ? _ram_0_T_5[63:0] : ram_0_100; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1006 = 7'h65 == index ? _ram_0_T_5[63:0] : ram_0_101; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1007 = 7'h66 == index ? _ram_0_T_5[63:0] : ram_0_102; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1008 = 7'h67 == index ? _ram_0_T_5[63:0] : ram_0_103; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1009 = 7'h68 == index ? _ram_0_T_5[63:0] : ram_0_104; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1010 = 7'h69 == index ? _ram_0_T_5[63:0] : ram_0_105; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1011 = 7'h6a == index ? _ram_0_T_5[63:0] : ram_0_106; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1012 = 7'h6b == index ? _ram_0_T_5[63:0] : ram_0_107; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1013 = 7'h6c == index ? _ram_0_T_5[63:0] : ram_0_108; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1014 = 7'h6d == index ? _ram_0_T_5[63:0] : ram_0_109; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1015 = 7'h6e == index ? _ram_0_T_5[63:0] : ram_0_110; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1016 = 7'h6f == index ? _ram_0_T_5[63:0] : ram_0_111; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1017 = 7'h70 == index ? _ram_0_T_5[63:0] : ram_0_112; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1018 = 7'h71 == index ? _ram_0_T_5[63:0] : ram_0_113; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1019 = 7'h72 == index ? _ram_0_T_5[63:0] : ram_0_114; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1020 = 7'h73 == index ? _ram_0_T_5[63:0] : ram_0_115; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1021 = 7'h74 == index ? _ram_0_T_5[63:0] : ram_0_116; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1022 = 7'h75 == index ? _ram_0_T_5[63:0] : ram_0_117; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1023 = 7'h76 == index ? _ram_0_T_5[63:0] : ram_0_118; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1024 = 7'h77 == index ? _ram_0_T_5[63:0] : ram_0_119; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1025 = 7'h78 == index ? _ram_0_T_5[63:0] : ram_0_120; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1026 = 7'h79 == index ? _ram_0_T_5[63:0] : ram_0_121; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1027 = 7'h7a == index ? _ram_0_T_5[63:0] : ram_0_122; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1028 = 7'h7b == index ? _ram_0_T_5[63:0] : ram_0_123; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1029 = 7'h7c == index ? _ram_0_T_5[63:0] : ram_0_124; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1030 = 7'h7d == index ? _ram_0_T_5[63:0] : ram_0_125; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1031 = 7'h7e == index ? _ram_0_T_5[63:0] : ram_0_126; // @[d_cache.scala 115:{30,30} 19:24]
  wire [63:0] _GEN_1032 = 7'h7f == index ? _ram_0_T_5[63:0] : ram_0_127; // @[d_cache.scala 115:{30,30} 19:24]
  wire  _GEN_19748 = 7'h0 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1033 = 7'h0 == index | dirty_0_0; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19749 = 7'h1 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1034 = 7'h1 == index | dirty_0_1; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19750 = 7'h2 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1035 = 7'h2 == index | dirty_0_2; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19751 = 7'h3 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1036 = 7'h3 == index | dirty_0_3; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19752 = 7'h4 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1037 = 7'h4 == index | dirty_0_4; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19753 = 7'h5 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1038 = 7'h5 == index | dirty_0_5; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19754 = 7'h6 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1039 = 7'h6 == index | dirty_0_6; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19755 = 7'h7 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1040 = 7'h7 == index | dirty_0_7; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19756 = 7'h8 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1041 = 7'h8 == index | dirty_0_8; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19757 = 7'h9 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1042 = 7'h9 == index | dirty_0_9; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19758 = 7'ha == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1043 = 7'ha == index | dirty_0_10; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19759 = 7'hb == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1044 = 7'hb == index | dirty_0_11; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19760 = 7'hc == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1045 = 7'hc == index | dirty_0_12; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19761 = 7'hd == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1046 = 7'hd == index | dirty_0_13; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19762 = 7'he == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1047 = 7'he == index | dirty_0_14; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19763 = 7'hf == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1048 = 7'hf == index | dirty_0_15; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19764 = 7'h10 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1049 = 7'h10 == index | dirty_0_16; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19765 = 7'h11 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1050 = 7'h11 == index | dirty_0_17; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19766 = 7'h12 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1051 = 7'h12 == index | dirty_0_18; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19767 = 7'h13 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1052 = 7'h13 == index | dirty_0_19; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19768 = 7'h14 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1053 = 7'h14 == index | dirty_0_20; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19769 = 7'h15 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1054 = 7'h15 == index | dirty_0_21; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19770 = 7'h16 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1055 = 7'h16 == index | dirty_0_22; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19771 = 7'h17 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1056 = 7'h17 == index | dirty_0_23; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19772 = 7'h18 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1057 = 7'h18 == index | dirty_0_24; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19773 = 7'h19 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1058 = 7'h19 == index | dirty_0_25; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19774 = 7'h1a == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1059 = 7'h1a == index | dirty_0_26; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19775 = 7'h1b == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1060 = 7'h1b == index | dirty_0_27; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19776 = 7'h1c == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1061 = 7'h1c == index | dirty_0_28; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19777 = 7'h1d == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1062 = 7'h1d == index | dirty_0_29; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19778 = 7'h1e == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1063 = 7'h1e == index | dirty_0_30; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19779 = 7'h1f == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1064 = 7'h1f == index | dirty_0_31; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19780 = 7'h20 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1065 = 7'h20 == index | dirty_0_32; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19781 = 7'h21 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1066 = 7'h21 == index | dirty_0_33; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19782 = 7'h22 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1067 = 7'h22 == index | dirty_0_34; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19783 = 7'h23 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1068 = 7'h23 == index | dirty_0_35; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19784 = 7'h24 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1069 = 7'h24 == index | dirty_0_36; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19785 = 7'h25 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1070 = 7'h25 == index | dirty_0_37; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19786 = 7'h26 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1071 = 7'h26 == index | dirty_0_38; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19787 = 7'h27 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1072 = 7'h27 == index | dirty_0_39; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19788 = 7'h28 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1073 = 7'h28 == index | dirty_0_40; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19789 = 7'h29 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1074 = 7'h29 == index | dirty_0_41; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19790 = 7'h2a == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1075 = 7'h2a == index | dirty_0_42; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19791 = 7'h2b == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1076 = 7'h2b == index | dirty_0_43; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19792 = 7'h2c == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1077 = 7'h2c == index | dirty_0_44; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19793 = 7'h2d == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1078 = 7'h2d == index | dirty_0_45; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19794 = 7'h2e == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1079 = 7'h2e == index | dirty_0_46; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19795 = 7'h2f == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1080 = 7'h2f == index | dirty_0_47; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19796 = 7'h30 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1081 = 7'h30 == index | dirty_0_48; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19797 = 7'h31 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1082 = 7'h31 == index | dirty_0_49; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19798 = 7'h32 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1083 = 7'h32 == index | dirty_0_50; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19799 = 7'h33 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1084 = 7'h33 == index | dirty_0_51; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19800 = 7'h34 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1085 = 7'h34 == index | dirty_0_52; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19801 = 7'h35 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1086 = 7'h35 == index | dirty_0_53; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19802 = 7'h36 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1087 = 7'h36 == index | dirty_0_54; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19803 = 7'h37 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1088 = 7'h37 == index | dirty_0_55; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19804 = 7'h38 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1089 = 7'h38 == index | dirty_0_56; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19805 = 7'h39 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1090 = 7'h39 == index | dirty_0_57; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19806 = 7'h3a == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1091 = 7'h3a == index | dirty_0_58; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19807 = 7'h3b == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1092 = 7'h3b == index | dirty_0_59; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19808 = 7'h3c == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1093 = 7'h3c == index | dirty_0_60; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19809 = 7'h3d == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1094 = 7'h3d == index | dirty_0_61; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19810 = 7'h3e == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1095 = 7'h3e == index | dirty_0_62; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19811 = 7'h3f == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1096 = 7'h3f == index | dirty_0_63; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19812 = 7'h40 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1097 = 7'h40 == index | dirty_0_64; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19813 = 7'h41 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1098 = 7'h41 == index | dirty_0_65; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19814 = 7'h42 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1099 = 7'h42 == index | dirty_0_66; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19815 = 7'h43 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1100 = 7'h43 == index | dirty_0_67; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19816 = 7'h44 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1101 = 7'h44 == index | dirty_0_68; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19817 = 7'h45 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1102 = 7'h45 == index | dirty_0_69; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19818 = 7'h46 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1103 = 7'h46 == index | dirty_0_70; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19819 = 7'h47 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1104 = 7'h47 == index | dirty_0_71; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19820 = 7'h48 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1105 = 7'h48 == index | dirty_0_72; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19821 = 7'h49 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1106 = 7'h49 == index | dirty_0_73; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19822 = 7'h4a == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1107 = 7'h4a == index | dirty_0_74; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19823 = 7'h4b == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1108 = 7'h4b == index | dirty_0_75; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19824 = 7'h4c == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1109 = 7'h4c == index | dirty_0_76; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19825 = 7'h4d == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1110 = 7'h4d == index | dirty_0_77; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19826 = 7'h4e == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1111 = 7'h4e == index | dirty_0_78; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19827 = 7'h4f == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1112 = 7'h4f == index | dirty_0_79; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19828 = 7'h50 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1113 = 7'h50 == index | dirty_0_80; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19829 = 7'h51 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1114 = 7'h51 == index | dirty_0_81; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19830 = 7'h52 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1115 = 7'h52 == index | dirty_0_82; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19831 = 7'h53 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1116 = 7'h53 == index | dirty_0_83; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19832 = 7'h54 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1117 = 7'h54 == index | dirty_0_84; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19833 = 7'h55 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1118 = 7'h55 == index | dirty_0_85; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19834 = 7'h56 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1119 = 7'h56 == index | dirty_0_86; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19835 = 7'h57 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1120 = 7'h57 == index | dirty_0_87; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19836 = 7'h58 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1121 = 7'h58 == index | dirty_0_88; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19837 = 7'h59 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1122 = 7'h59 == index | dirty_0_89; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19838 = 7'h5a == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1123 = 7'h5a == index | dirty_0_90; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19839 = 7'h5b == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1124 = 7'h5b == index | dirty_0_91; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19840 = 7'h5c == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1125 = 7'h5c == index | dirty_0_92; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19841 = 7'h5d == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1126 = 7'h5d == index | dirty_0_93; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19842 = 7'h5e == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1127 = 7'h5e == index | dirty_0_94; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19843 = 7'h5f == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1128 = 7'h5f == index | dirty_0_95; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19844 = 7'h60 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1129 = 7'h60 == index | dirty_0_96; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19845 = 7'h61 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1130 = 7'h61 == index | dirty_0_97; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19846 = 7'h62 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1131 = 7'h62 == index | dirty_0_98; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19847 = 7'h63 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1132 = 7'h63 == index | dirty_0_99; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19848 = 7'h64 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1133 = 7'h64 == index | dirty_0_100; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19849 = 7'h65 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1134 = 7'h65 == index | dirty_0_101; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19850 = 7'h66 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1135 = 7'h66 == index | dirty_0_102; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19851 = 7'h67 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1136 = 7'h67 == index | dirty_0_103; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19852 = 7'h68 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1137 = 7'h68 == index | dirty_0_104; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19853 = 7'h69 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1138 = 7'h69 == index | dirty_0_105; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19854 = 7'h6a == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1139 = 7'h6a == index | dirty_0_106; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19855 = 7'h6b == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1140 = 7'h6b == index | dirty_0_107; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19856 = 7'h6c == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1141 = 7'h6c == index | dirty_0_108; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19857 = 7'h6d == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1142 = 7'h6d == index | dirty_0_109; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19858 = 7'h6e == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1143 = 7'h6e == index | dirty_0_110; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19859 = 7'h6f == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1144 = 7'h6f == index | dirty_0_111; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19860 = 7'h70 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1145 = 7'h70 == index | dirty_0_112; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19861 = 7'h71 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1146 = 7'h71 == index | dirty_0_113; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19862 = 7'h72 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1147 = 7'h72 == index | dirty_0_114; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19863 = 7'h73 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1148 = 7'h73 == index | dirty_0_115; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19864 = 7'h74 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1149 = 7'h74 == index | dirty_0_116; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19865 = 7'h75 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1150 = 7'h75 == index | dirty_0_117; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19866 = 7'h76 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1151 = 7'h76 == index | dirty_0_118; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19867 = 7'h77 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1152 = 7'h77 == index | dirty_0_119; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19868 = 7'h78 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1153 = 7'h78 == index | dirty_0_120; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19869 = 7'h79 == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1154 = 7'h79 == index | dirty_0_121; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19870 = 7'h7a == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1155 = 7'h7a == index | dirty_0_122; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19871 = 7'h7b == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1156 = 7'h7b == index | dirty_0_123; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19872 = 7'h7c == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1157 = 7'h7c == index | dirty_0_124; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19873 = 7'h7d == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1158 = 7'h7d == index | dirty_0_125; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19874 = 7'h7e == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1159 = 7'h7e == index | dirty_0_126; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_19875 = 7'h7f == index; // @[d_cache.scala 119:{32,32} 32:26]
  wire  _GEN_1160 = 7'h7f == index | dirty_0_127; // @[d_cache.scala 119:{32,32} 32:26]
  wire [63:0] _GEN_1290 = 7'h1 == index ? ram_1_1 : ram_1_0; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1291 = 7'h2 == index ? ram_1_2 : _GEN_1290; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1292 = 7'h3 == index ? ram_1_3 : _GEN_1291; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1293 = 7'h4 == index ? ram_1_4 : _GEN_1292; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1294 = 7'h5 == index ? ram_1_5 : _GEN_1293; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1295 = 7'h6 == index ? ram_1_6 : _GEN_1294; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1296 = 7'h7 == index ? ram_1_7 : _GEN_1295; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1297 = 7'h8 == index ? ram_1_8 : _GEN_1296; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1298 = 7'h9 == index ? ram_1_9 : _GEN_1297; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1299 = 7'ha == index ? ram_1_10 : _GEN_1298; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1300 = 7'hb == index ? ram_1_11 : _GEN_1299; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1301 = 7'hc == index ? ram_1_12 : _GEN_1300; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1302 = 7'hd == index ? ram_1_13 : _GEN_1301; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1303 = 7'he == index ? ram_1_14 : _GEN_1302; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1304 = 7'hf == index ? ram_1_15 : _GEN_1303; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1305 = 7'h10 == index ? ram_1_16 : _GEN_1304; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1306 = 7'h11 == index ? ram_1_17 : _GEN_1305; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1307 = 7'h12 == index ? ram_1_18 : _GEN_1306; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1308 = 7'h13 == index ? ram_1_19 : _GEN_1307; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1309 = 7'h14 == index ? ram_1_20 : _GEN_1308; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1310 = 7'h15 == index ? ram_1_21 : _GEN_1309; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1311 = 7'h16 == index ? ram_1_22 : _GEN_1310; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1312 = 7'h17 == index ? ram_1_23 : _GEN_1311; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1313 = 7'h18 == index ? ram_1_24 : _GEN_1312; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1314 = 7'h19 == index ? ram_1_25 : _GEN_1313; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1315 = 7'h1a == index ? ram_1_26 : _GEN_1314; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1316 = 7'h1b == index ? ram_1_27 : _GEN_1315; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1317 = 7'h1c == index ? ram_1_28 : _GEN_1316; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1318 = 7'h1d == index ? ram_1_29 : _GEN_1317; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1319 = 7'h1e == index ? ram_1_30 : _GEN_1318; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1320 = 7'h1f == index ? ram_1_31 : _GEN_1319; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1321 = 7'h20 == index ? ram_1_32 : _GEN_1320; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1322 = 7'h21 == index ? ram_1_33 : _GEN_1321; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1323 = 7'h22 == index ? ram_1_34 : _GEN_1322; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1324 = 7'h23 == index ? ram_1_35 : _GEN_1323; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1325 = 7'h24 == index ? ram_1_36 : _GEN_1324; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1326 = 7'h25 == index ? ram_1_37 : _GEN_1325; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1327 = 7'h26 == index ? ram_1_38 : _GEN_1326; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1328 = 7'h27 == index ? ram_1_39 : _GEN_1327; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1329 = 7'h28 == index ? ram_1_40 : _GEN_1328; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1330 = 7'h29 == index ? ram_1_41 : _GEN_1329; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1331 = 7'h2a == index ? ram_1_42 : _GEN_1330; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1332 = 7'h2b == index ? ram_1_43 : _GEN_1331; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1333 = 7'h2c == index ? ram_1_44 : _GEN_1332; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1334 = 7'h2d == index ? ram_1_45 : _GEN_1333; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1335 = 7'h2e == index ? ram_1_46 : _GEN_1334; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1336 = 7'h2f == index ? ram_1_47 : _GEN_1335; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1337 = 7'h30 == index ? ram_1_48 : _GEN_1336; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1338 = 7'h31 == index ? ram_1_49 : _GEN_1337; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1339 = 7'h32 == index ? ram_1_50 : _GEN_1338; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1340 = 7'h33 == index ? ram_1_51 : _GEN_1339; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1341 = 7'h34 == index ? ram_1_52 : _GEN_1340; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1342 = 7'h35 == index ? ram_1_53 : _GEN_1341; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1343 = 7'h36 == index ? ram_1_54 : _GEN_1342; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1344 = 7'h37 == index ? ram_1_55 : _GEN_1343; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1345 = 7'h38 == index ? ram_1_56 : _GEN_1344; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1346 = 7'h39 == index ? ram_1_57 : _GEN_1345; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1347 = 7'h3a == index ? ram_1_58 : _GEN_1346; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1348 = 7'h3b == index ? ram_1_59 : _GEN_1347; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1349 = 7'h3c == index ? ram_1_60 : _GEN_1348; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1350 = 7'h3d == index ? ram_1_61 : _GEN_1349; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1351 = 7'h3e == index ? ram_1_62 : _GEN_1350; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1352 = 7'h3f == index ? ram_1_63 : _GEN_1351; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1353 = 7'h40 == index ? ram_1_64 : _GEN_1352; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1354 = 7'h41 == index ? ram_1_65 : _GEN_1353; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1355 = 7'h42 == index ? ram_1_66 : _GEN_1354; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1356 = 7'h43 == index ? ram_1_67 : _GEN_1355; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1357 = 7'h44 == index ? ram_1_68 : _GEN_1356; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1358 = 7'h45 == index ? ram_1_69 : _GEN_1357; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1359 = 7'h46 == index ? ram_1_70 : _GEN_1358; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1360 = 7'h47 == index ? ram_1_71 : _GEN_1359; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1361 = 7'h48 == index ? ram_1_72 : _GEN_1360; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1362 = 7'h49 == index ? ram_1_73 : _GEN_1361; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1363 = 7'h4a == index ? ram_1_74 : _GEN_1362; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1364 = 7'h4b == index ? ram_1_75 : _GEN_1363; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1365 = 7'h4c == index ? ram_1_76 : _GEN_1364; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1366 = 7'h4d == index ? ram_1_77 : _GEN_1365; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1367 = 7'h4e == index ? ram_1_78 : _GEN_1366; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1368 = 7'h4f == index ? ram_1_79 : _GEN_1367; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1369 = 7'h50 == index ? ram_1_80 : _GEN_1368; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1370 = 7'h51 == index ? ram_1_81 : _GEN_1369; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1371 = 7'h52 == index ? ram_1_82 : _GEN_1370; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1372 = 7'h53 == index ? ram_1_83 : _GEN_1371; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1373 = 7'h54 == index ? ram_1_84 : _GEN_1372; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1374 = 7'h55 == index ? ram_1_85 : _GEN_1373; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1375 = 7'h56 == index ? ram_1_86 : _GEN_1374; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1376 = 7'h57 == index ? ram_1_87 : _GEN_1375; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1377 = 7'h58 == index ? ram_1_88 : _GEN_1376; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1378 = 7'h59 == index ? ram_1_89 : _GEN_1377; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1379 = 7'h5a == index ? ram_1_90 : _GEN_1378; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1380 = 7'h5b == index ? ram_1_91 : _GEN_1379; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1381 = 7'h5c == index ? ram_1_92 : _GEN_1380; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1382 = 7'h5d == index ? ram_1_93 : _GEN_1381; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1383 = 7'h5e == index ? ram_1_94 : _GEN_1382; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1384 = 7'h5f == index ? ram_1_95 : _GEN_1383; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1385 = 7'h60 == index ? ram_1_96 : _GEN_1384; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1386 = 7'h61 == index ? ram_1_97 : _GEN_1385; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1387 = 7'h62 == index ? ram_1_98 : _GEN_1386; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1388 = 7'h63 == index ? ram_1_99 : _GEN_1387; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1389 = 7'h64 == index ? ram_1_100 : _GEN_1388; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1390 = 7'h65 == index ? ram_1_101 : _GEN_1389; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1391 = 7'h66 == index ? ram_1_102 : _GEN_1390; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1392 = 7'h67 == index ? ram_1_103 : _GEN_1391; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1393 = 7'h68 == index ? ram_1_104 : _GEN_1392; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1394 = 7'h69 == index ? ram_1_105 : _GEN_1393; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1395 = 7'h6a == index ? ram_1_106 : _GEN_1394; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1396 = 7'h6b == index ? ram_1_107 : _GEN_1395; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1397 = 7'h6c == index ? ram_1_108 : _GEN_1396; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1398 = 7'h6d == index ? ram_1_109 : _GEN_1397; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1399 = 7'h6e == index ? ram_1_110 : _GEN_1398; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1400 = 7'h6f == index ? ram_1_111 : _GEN_1399; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1401 = 7'h70 == index ? ram_1_112 : _GEN_1400; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1402 = 7'h71 == index ? ram_1_113 : _GEN_1401; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1403 = 7'h72 == index ? ram_1_114 : _GEN_1402; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1404 = 7'h73 == index ? ram_1_115 : _GEN_1403; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1405 = 7'h74 == index ? ram_1_116 : _GEN_1404; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1406 = 7'h75 == index ? ram_1_117 : _GEN_1405; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1407 = 7'h76 == index ? ram_1_118 : _GEN_1406; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1408 = 7'h77 == index ? ram_1_119 : _GEN_1407; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1409 = 7'h78 == index ? ram_1_120 : _GEN_1408; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1410 = 7'h79 == index ? ram_1_121 : _GEN_1409; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1411 = 7'h7a == index ? ram_1_122 : _GEN_1410; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1412 = 7'h7b == index ? ram_1_123 : _GEN_1411; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1413 = 7'h7c == index ? ram_1_124 : _GEN_1412; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1414 = 7'h7d == index ? ram_1_125 : _GEN_1413; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1415 = 7'h7e == index ? ram_1_126 : _GEN_1414; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1416 = 7'h7f == index ? ram_1_127 : _GEN_1415; // @[d_cache.scala 123:{39,39}]
  wire [63:0] _GEN_1161 = 7'h0 == index ? _GEN_1416 : record_olddata_0; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1162 = 7'h1 == index ? _GEN_1416 : record_olddata_1; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1163 = 7'h2 == index ? _GEN_1416 : record_olddata_2; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1164 = 7'h3 == index ? _GEN_1416 : record_olddata_3; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1165 = 7'h4 == index ? _GEN_1416 : record_olddata_4; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1166 = 7'h5 == index ? _GEN_1416 : record_olddata_5; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1167 = 7'h6 == index ? _GEN_1416 : record_olddata_6; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1168 = 7'h7 == index ? _GEN_1416 : record_olddata_7; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1169 = 7'h8 == index ? _GEN_1416 : record_olddata_8; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1170 = 7'h9 == index ? _GEN_1416 : record_olddata_9; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1171 = 7'ha == index ? _GEN_1416 : record_olddata_10; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1172 = 7'hb == index ? _GEN_1416 : record_olddata_11; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1173 = 7'hc == index ? _GEN_1416 : record_olddata_12; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1174 = 7'hd == index ? _GEN_1416 : record_olddata_13; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1175 = 7'he == index ? _GEN_1416 : record_olddata_14; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1176 = 7'hf == index ? _GEN_1416 : record_olddata_15; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1177 = 7'h10 == index ? _GEN_1416 : record_olddata_16; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1178 = 7'h11 == index ? _GEN_1416 : record_olddata_17; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1179 = 7'h12 == index ? _GEN_1416 : record_olddata_18; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1180 = 7'h13 == index ? _GEN_1416 : record_olddata_19; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1181 = 7'h14 == index ? _GEN_1416 : record_olddata_20; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1182 = 7'h15 == index ? _GEN_1416 : record_olddata_21; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1183 = 7'h16 == index ? _GEN_1416 : record_olddata_22; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1184 = 7'h17 == index ? _GEN_1416 : record_olddata_23; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1185 = 7'h18 == index ? _GEN_1416 : record_olddata_24; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1186 = 7'h19 == index ? _GEN_1416 : record_olddata_25; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1187 = 7'h1a == index ? _GEN_1416 : record_olddata_26; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1188 = 7'h1b == index ? _GEN_1416 : record_olddata_27; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1189 = 7'h1c == index ? _GEN_1416 : record_olddata_28; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1190 = 7'h1d == index ? _GEN_1416 : record_olddata_29; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1191 = 7'h1e == index ? _GEN_1416 : record_olddata_30; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1192 = 7'h1f == index ? _GEN_1416 : record_olddata_31; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1193 = 7'h20 == index ? _GEN_1416 : record_olddata_32; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1194 = 7'h21 == index ? _GEN_1416 : record_olddata_33; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1195 = 7'h22 == index ? _GEN_1416 : record_olddata_34; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1196 = 7'h23 == index ? _GEN_1416 : record_olddata_35; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1197 = 7'h24 == index ? _GEN_1416 : record_olddata_36; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1198 = 7'h25 == index ? _GEN_1416 : record_olddata_37; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1199 = 7'h26 == index ? _GEN_1416 : record_olddata_38; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1200 = 7'h27 == index ? _GEN_1416 : record_olddata_39; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1201 = 7'h28 == index ? _GEN_1416 : record_olddata_40; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1202 = 7'h29 == index ? _GEN_1416 : record_olddata_41; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1203 = 7'h2a == index ? _GEN_1416 : record_olddata_42; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1204 = 7'h2b == index ? _GEN_1416 : record_olddata_43; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1205 = 7'h2c == index ? _GEN_1416 : record_olddata_44; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1206 = 7'h2d == index ? _GEN_1416 : record_olddata_45; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1207 = 7'h2e == index ? _GEN_1416 : record_olddata_46; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1208 = 7'h2f == index ? _GEN_1416 : record_olddata_47; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1209 = 7'h30 == index ? _GEN_1416 : record_olddata_48; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1210 = 7'h31 == index ? _GEN_1416 : record_olddata_49; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1211 = 7'h32 == index ? _GEN_1416 : record_olddata_50; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1212 = 7'h33 == index ? _GEN_1416 : record_olddata_51; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1213 = 7'h34 == index ? _GEN_1416 : record_olddata_52; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1214 = 7'h35 == index ? _GEN_1416 : record_olddata_53; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1215 = 7'h36 == index ? _GEN_1416 : record_olddata_54; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1216 = 7'h37 == index ? _GEN_1416 : record_olddata_55; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1217 = 7'h38 == index ? _GEN_1416 : record_olddata_56; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1218 = 7'h39 == index ? _GEN_1416 : record_olddata_57; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1219 = 7'h3a == index ? _GEN_1416 : record_olddata_58; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1220 = 7'h3b == index ? _GEN_1416 : record_olddata_59; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1221 = 7'h3c == index ? _GEN_1416 : record_olddata_60; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1222 = 7'h3d == index ? _GEN_1416 : record_olddata_61; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1223 = 7'h3e == index ? _GEN_1416 : record_olddata_62; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1224 = 7'h3f == index ? _GEN_1416 : record_olddata_63; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1225 = 7'h40 == index ? _GEN_1416 : record_olddata_64; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1226 = 7'h41 == index ? _GEN_1416 : record_olddata_65; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1227 = 7'h42 == index ? _GEN_1416 : record_olddata_66; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1228 = 7'h43 == index ? _GEN_1416 : record_olddata_67; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1229 = 7'h44 == index ? _GEN_1416 : record_olddata_68; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1230 = 7'h45 == index ? _GEN_1416 : record_olddata_69; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1231 = 7'h46 == index ? _GEN_1416 : record_olddata_70; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1232 = 7'h47 == index ? _GEN_1416 : record_olddata_71; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1233 = 7'h48 == index ? _GEN_1416 : record_olddata_72; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1234 = 7'h49 == index ? _GEN_1416 : record_olddata_73; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1235 = 7'h4a == index ? _GEN_1416 : record_olddata_74; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1236 = 7'h4b == index ? _GEN_1416 : record_olddata_75; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1237 = 7'h4c == index ? _GEN_1416 : record_olddata_76; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1238 = 7'h4d == index ? _GEN_1416 : record_olddata_77; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1239 = 7'h4e == index ? _GEN_1416 : record_olddata_78; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1240 = 7'h4f == index ? _GEN_1416 : record_olddata_79; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1241 = 7'h50 == index ? _GEN_1416 : record_olddata_80; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1242 = 7'h51 == index ? _GEN_1416 : record_olddata_81; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1243 = 7'h52 == index ? _GEN_1416 : record_olddata_82; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1244 = 7'h53 == index ? _GEN_1416 : record_olddata_83; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1245 = 7'h54 == index ? _GEN_1416 : record_olddata_84; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1246 = 7'h55 == index ? _GEN_1416 : record_olddata_85; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1247 = 7'h56 == index ? _GEN_1416 : record_olddata_86; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1248 = 7'h57 == index ? _GEN_1416 : record_olddata_87; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1249 = 7'h58 == index ? _GEN_1416 : record_olddata_88; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1250 = 7'h59 == index ? _GEN_1416 : record_olddata_89; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1251 = 7'h5a == index ? _GEN_1416 : record_olddata_90; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1252 = 7'h5b == index ? _GEN_1416 : record_olddata_91; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1253 = 7'h5c == index ? _GEN_1416 : record_olddata_92; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1254 = 7'h5d == index ? _GEN_1416 : record_olddata_93; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1255 = 7'h5e == index ? _GEN_1416 : record_olddata_94; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1256 = 7'h5f == index ? _GEN_1416 : record_olddata_95; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1257 = 7'h60 == index ? _GEN_1416 : record_olddata_96; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1258 = 7'h61 == index ? _GEN_1416 : record_olddata_97; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1259 = 7'h62 == index ? _GEN_1416 : record_olddata_98; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1260 = 7'h63 == index ? _GEN_1416 : record_olddata_99; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1261 = 7'h64 == index ? _GEN_1416 : record_olddata_100; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1262 = 7'h65 == index ? _GEN_1416 : record_olddata_101; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1263 = 7'h66 == index ? _GEN_1416 : record_olddata_102; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1264 = 7'h67 == index ? _GEN_1416 : record_olddata_103; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1265 = 7'h68 == index ? _GEN_1416 : record_olddata_104; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1266 = 7'h69 == index ? _GEN_1416 : record_olddata_105; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1267 = 7'h6a == index ? _GEN_1416 : record_olddata_106; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1268 = 7'h6b == index ? _GEN_1416 : record_olddata_107; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1269 = 7'h6c == index ? _GEN_1416 : record_olddata_108; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1270 = 7'h6d == index ? _GEN_1416 : record_olddata_109; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1271 = 7'h6e == index ? _GEN_1416 : record_olddata_110; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1272 = 7'h6f == index ? _GEN_1416 : record_olddata_111; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1273 = 7'h70 == index ? _GEN_1416 : record_olddata_112; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1274 = 7'h71 == index ? _GEN_1416 : record_olddata_113; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1275 = 7'h72 == index ? _GEN_1416 : record_olddata_114; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1276 = 7'h73 == index ? _GEN_1416 : record_olddata_115; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1277 = 7'h74 == index ? _GEN_1416 : record_olddata_116; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1278 = 7'h75 == index ? _GEN_1416 : record_olddata_117; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1279 = 7'h76 == index ? _GEN_1416 : record_olddata_118; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1280 = 7'h77 == index ? _GEN_1416 : record_olddata_119; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1281 = 7'h78 == index ? _GEN_1416 : record_olddata_120; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1282 = 7'h79 == index ? _GEN_1416 : record_olddata_121; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1283 = 7'h7a == index ? _GEN_1416 : record_olddata_122; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1284 = 7'h7b == index ? _GEN_1416 : record_olddata_123; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1285 = 7'h7c == index ? _GEN_1416 : record_olddata_124; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1286 = 7'h7d == index ? _GEN_1416 : record_olddata_125; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1287 = 7'h7e == index ? _GEN_1416 : record_olddata_126; // @[d_cache.scala 123:{39,39} 25:33]
  wire [63:0] _GEN_1288 = 7'h7f == index ? _GEN_1416 : record_olddata_127; // @[d_cache.scala 123:{39,39} 25:33]
  wire [126:0] _GEN_19876 = {{63'd0}, _GEN_1416}; // @[d_cache.scala 124:92]
  wire [126:0] _ram_1_T_4 = _GEN_19876 & _ram_0_T_3; // @[d_cache.scala 124:92]
  wire [126:0] _ram_1_T_5 = _ram_0_T_1 | _ram_1_T_4; // @[d_cache.scala 124:76]
  wire [63:0] _GEN_1417 = 7'h0 == index ? _ram_1_T_5[63:0] : ram_1_0; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1418 = 7'h1 == index ? _ram_1_T_5[63:0] : ram_1_1; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1419 = 7'h2 == index ? _ram_1_T_5[63:0] : ram_1_2; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1420 = 7'h3 == index ? _ram_1_T_5[63:0] : ram_1_3; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1421 = 7'h4 == index ? _ram_1_T_5[63:0] : ram_1_4; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1422 = 7'h5 == index ? _ram_1_T_5[63:0] : ram_1_5; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1423 = 7'h6 == index ? _ram_1_T_5[63:0] : ram_1_6; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1424 = 7'h7 == index ? _ram_1_T_5[63:0] : ram_1_7; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1425 = 7'h8 == index ? _ram_1_T_5[63:0] : ram_1_8; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1426 = 7'h9 == index ? _ram_1_T_5[63:0] : ram_1_9; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1427 = 7'ha == index ? _ram_1_T_5[63:0] : ram_1_10; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1428 = 7'hb == index ? _ram_1_T_5[63:0] : ram_1_11; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1429 = 7'hc == index ? _ram_1_T_5[63:0] : ram_1_12; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1430 = 7'hd == index ? _ram_1_T_5[63:0] : ram_1_13; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1431 = 7'he == index ? _ram_1_T_5[63:0] : ram_1_14; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1432 = 7'hf == index ? _ram_1_T_5[63:0] : ram_1_15; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1433 = 7'h10 == index ? _ram_1_T_5[63:0] : ram_1_16; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1434 = 7'h11 == index ? _ram_1_T_5[63:0] : ram_1_17; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1435 = 7'h12 == index ? _ram_1_T_5[63:0] : ram_1_18; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1436 = 7'h13 == index ? _ram_1_T_5[63:0] : ram_1_19; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1437 = 7'h14 == index ? _ram_1_T_5[63:0] : ram_1_20; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1438 = 7'h15 == index ? _ram_1_T_5[63:0] : ram_1_21; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1439 = 7'h16 == index ? _ram_1_T_5[63:0] : ram_1_22; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1440 = 7'h17 == index ? _ram_1_T_5[63:0] : ram_1_23; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1441 = 7'h18 == index ? _ram_1_T_5[63:0] : ram_1_24; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1442 = 7'h19 == index ? _ram_1_T_5[63:0] : ram_1_25; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1443 = 7'h1a == index ? _ram_1_T_5[63:0] : ram_1_26; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1444 = 7'h1b == index ? _ram_1_T_5[63:0] : ram_1_27; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1445 = 7'h1c == index ? _ram_1_T_5[63:0] : ram_1_28; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1446 = 7'h1d == index ? _ram_1_T_5[63:0] : ram_1_29; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1447 = 7'h1e == index ? _ram_1_T_5[63:0] : ram_1_30; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1448 = 7'h1f == index ? _ram_1_T_5[63:0] : ram_1_31; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1449 = 7'h20 == index ? _ram_1_T_5[63:0] : ram_1_32; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1450 = 7'h21 == index ? _ram_1_T_5[63:0] : ram_1_33; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1451 = 7'h22 == index ? _ram_1_T_5[63:0] : ram_1_34; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1452 = 7'h23 == index ? _ram_1_T_5[63:0] : ram_1_35; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1453 = 7'h24 == index ? _ram_1_T_5[63:0] : ram_1_36; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1454 = 7'h25 == index ? _ram_1_T_5[63:0] : ram_1_37; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1455 = 7'h26 == index ? _ram_1_T_5[63:0] : ram_1_38; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1456 = 7'h27 == index ? _ram_1_T_5[63:0] : ram_1_39; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1457 = 7'h28 == index ? _ram_1_T_5[63:0] : ram_1_40; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1458 = 7'h29 == index ? _ram_1_T_5[63:0] : ram_1_41; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1459 = 7'h2a == index ? _ram_1_T_5[63:0] : ram_1_42; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1460 = 7'h2b == index ? _ram_1_T_5[63:0] : ram_1_43; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1461 = 7'h2c == index ? _ram_1_T_5[63:0] : ram_1_44; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1462 = 7'h2d == index ? _ram_1_T_5[63:0] : ram_1_45; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1463 = 7'h2e == index ? _ram_1_T_5[63:0] : ram_1_46; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1464 = 7'h2f == index ? _ram_1_T_5[63:0] : ram_1_47; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1465 = 7'h30 == index ? _ram_1_T_5[63:0] : ram_1_48; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1466 = 7'h31 == index ? _ram_1_T_5[63:0] : ram_1_49; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1467 = 7'h32 == index ? _ram_1_T_5[63:0] : ram_1_50; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1468 = 7'h33 == index ? _ram_1_T_5[63:0] : ram_1_51; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1469 = 7'h34 == index ? _ram_1_T_5[63:0] : ram_1_52; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1470 = 7'h35 == index ? _ram_1_T_5[63:0] : ram_1_53; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1471 = 7'h36 == index ? _ram_1_T_5[63:0] : ram_1_54; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1472 = 7'h37 == index ? _ram_1_T_5[63:0] : ram_1_55; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1473 = 7'h38 == index ? _ram_1_T_5[63:0] : ram_1_56; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1474 = 7'h39 == index ? _ram_1_T_5[63:0] : ram_1_57; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1475 = 7'h3a == index ? _ram_1_T_5[63:0] : ram_1_58; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1476 = 7'h3b == index ? _ram_1_T_5[63:0] : ram_1_59; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1477 = 7'h3c == index ? _ram_1_T_5[63:0] : ram_1_60; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1478 = 7'h3d == index ? _ram_1_T_5[63:0] : ram_1_61; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1479 = 7'h3e == index ? _ram_1_T_5[63:0] : ram_1_62; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1480 = 7'h3f == index ? _ram_1_T_5[63:0] : ram_1_63; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1481 = 7'h40 == index ? _ram_1_T_5[63:0] : ram_1_64; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1482 = 7'h41 == index ? _ram_1_T_5[63:0] : ram_1_65; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1483 = 7'h42 == index ? _ram_1_T_5[63:0] : ram_1_66; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1484 = 7'h43 == index ? _ram_1_T_5[63:0] : ram_1_67; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1485 = 7'h44 == index ? _ram_1_T_5[63:0] : ram_1_68; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1486 = 7'h45 == index ? _ram_1_T_5[63:0] : ram_1_69; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1487 = 7'h46 == index ? _ram_1_T_5[63:0] : ram_1_70; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1488 = 7'h47 == index ? _ram_1_T_5[63:0] : ram_1_71; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1489 = 7'h48 == index ? _ram_1_T_5[63:0] : ram_1_72; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1490 = 7'h49 == index ? _ram_1_T_5[63:0] : ram_1_73; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1491 = 7'h4a == index ? _ram_1_T_5[63:0] : ram_1_74; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1492 = 7'h4b == index ? _ram_1_T_5[63:0] : ram_1_75; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1493 = 7'h4c == index ? _ram_1_T_5[63:0] : ram_1_76; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1494 = 7'h4d == index ? _ram_1_T_5[63:0] : ram_1_77; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1495 = 7'h4e == index ? _ram_1_T_5[63:0] : ram_1_78; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1496 = 7'h4f == index ? _ram_1_T_5[63:0] : ram_1_79; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1497 = 7'h50 == index ? _ram_1_T_5[63:0] : ram_1_80; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1498 = 7'h51 == index ? _ram_1_T_5[63:0] : ram_1_81; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1499 = 7'h52 == index ? _ram_1_T_5[63:0] : ram_1_82; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1500 = 7'h53 == index ? _ram_1_T_5[63:0] : ram_1_83; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1501 = 7'h54 == index ? _ram_1_T_5[63:0] : ram_1_84; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1502 = 7'h55 == index ? _ram_1_T_5[63:0] : ram_1_85; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1503 = 7'h56 == index ? _ram_1_T_5[63:0] : ram_1_86; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1504 = 7'h57 == index ? _ram_1_T_5[63:0] : ram_1_87; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1505 = 7'h58 == index ? _ram_1_T_5[63:0] : ram_1_88; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1506 = 7'h59 == index ? _ram_1_T_5[63:0] : ram_1_89; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1507 = 7'h5a == index ? _ram_1_T_5[63:0] : ram_1_90; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1508 = 7'h5b == index ? _ram_1_T_5[63:0] : ram_1_91; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1509 = 7'h5c == index ? _ram_1_T_5[63:0] : ram_1_92; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1510 = 7'h5d == index ? _ram_1_T_5[63:0] : ram_1_93; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1511 = 7'h5e == index ? _ram_1_T_5[63:0] : ram_1_94; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1512 = 7'h5f == index ? _ram_1_T_5[63:0] : ram_1_95; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1513 = 7'h60 == index ? _ram_1_T_5[63:0] : ram_1_96; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1514 = 7'h61 == index ? _ram_1_T_5[63:0] : ram_1_97; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1515 = 7'h62 == index ? _ram_1_T_5[63:0] : ram_1_98; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1516 = 7'h63 == index ? _ram_1_T_5[63:0] : ram_1_99; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1517 = 7'h64 == index ? _ram_1_T_5[63:0] : ram_1_100; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1518 = 7'h65 == index ? _ram_1_T_5[63:0] : ram_1_101; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1519 = 7'h66 == index ? _ram_1_T_5[63:0] : ram_1_102; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1520 = 7'h67 == index ? _ram_1_T_5[63:0] : ram_1_103; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1521 = 7'h68 == index ? _ram_1_T_5[63:0] : ram_1_104; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1522 = 7'h69 == index ? _ram_1_T_5[63:0] : ram_1_105; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1523 = 7'h6a == index ? _ram_1_T_5[63:0] : ram_1_106; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1524 = 7'h6b == index ? _ram_1_T_5[63:0] : ram_1_107; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1525 = 7'h6c == index ? _ram_1_T_5[63:0] : ram_1_108; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1526 = 7'h6d == index ? _ram_1_T_5[63:0] : ram_1_109; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1527 = 7'h6e == index ? _ram_1_T_5[63:0] : ram_1_110; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1528 = 7'h6f == index ? _ram_1_T_5[63:0] : ram_1_111; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1529 = 7'h70 == index ? _ram_1_T_5[63:0] : ram_1_112; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1530 = 7'h71 == index ? _ram_1_T_5[63:0] : ram_1_113; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1531 = 7'h72 == index ? _ram_1_T_5[63:0] : ram_1_114; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1532 = 7'h73 == index ? _ram_1_T_5[63:0] : ram_1_115; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1533 = 7'h74 == index ? _ram_1_T_5[63:0] : ram_1_116; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1534 = 7'h75 == index ? _ram_1_T_5[63:0] : ram_1_117; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1535 = 7'h76 == index ? _ram_1_T_5[63:0] : ram_1_118; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1536 = 7'h77 == index ? _ram_1_T_5[63:0] : ram_1_119; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1537 = 7'h78 == index ? _ram_1_T_5[63:0] : ram_1_120; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1538 = 7'h79 == index ? _ram_1_T_5[63:0] : ram_1_121; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1539 = 7'h7a == index ? _ram_1_T_5[63:0] : ram_1_122; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1540 = 7'h7b == index ? _ram_1_T_5[63:0] : ram_1_123; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1541 = 7'h7c == index ? _ram_1_T_5[63:0] : ram_1_124; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1542 = 7'h7d == index ? _ram_1_T_5[63:0] : ram_1_125; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1543 = 7'h7e == index ? _ram_1_T_5[63:0] : ram_1_126; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1544 = 7'h7f == index ? _ram_1_T_5[63:0] : ram_1_127; // @[d_cache.scala 124:{30,30} 20:24]
  wire [63:0] _GEN_1545 = 7'h0 == index ? io_from_lsu_wdata : record_wdata1_0; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1546 = 7'h1 == index ? io_from_lsu_wdata : record_wdata1_1; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1547 = 7'h2 == index ? io_from_lsu_wdata : record_wdata1_2; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1548 = 7'h3 == index ? io_from_lsu_wdata : record_wdata1_3; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1549 = 7'h4 == index ? io_from_lsu_wdata : record_wdata1_4; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1550 = 7'h5 == index ? io_from_lsu_wdata : record_wdata1_5; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1551 = 7'h6 == index ? io_from_lsu_wdata : record_wdata1_6; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1552 = 7'h7 == index ? io_from_lsu_wdata : record_wdata1_7; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1553 = 7'h8 == index ? io_from_lsu_wdata : record_wdata1_8; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1554 = 7'h9 == index ? io_from_lsu_wdata : record_wdata1_9; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1555 = 7'ha == index ? io_from_lsu_wdata : record_wdata1_10; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1556 = 7'hb == index ? io_from_lsu_wdata : record_wdata1_11; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1557 = 7'hc == index ? io_from_lsu_wdata : record_wdata1_12; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1558 = 7'hd == index ? io_from_lsu_wdata : record_wdata1_13; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1559 = 7'he == index ? io_from_lsu_wdata : record_wdata1_14; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1560 = 7'hf == index ? io_from_lsu_wdata : record_wdata1_15; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1561 = 7'h10 == index ? io_from_lsu_wdata : record_wdata1_16; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1562 = 7'h11 == index ? io_from_lsu_wdata : record_wdata1_17; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1563 = 7'h12 == index ? io_from_lsu_wdata : record_wdata1_18; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1564 = 7'h13 == index ? io_from_lsu_wdata : record_wdata1_19; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1565 = 7'h14 == index ? io_from_lsu_wdata : record_wdata1_20; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1566 = 7'h15 == index ? io_from_lsu_wdata : record_wdata1_21; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1567 = 7'h16 == index ? io_from_lsu_wdata : record_wdata1_22; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1568 = 7'h17 == index ? io_from_lsu_wdata : record_wdata1_23; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1569 = 7'h18 == index ? io_from_lsu_wdata : record_wdata1_24; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1570 = 7'h19 == index ? io_from_lsu_wdata : record_wdata1_25; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1571 = 7'h1a == index ? io_from_lsu_wdata : record_wdata1_26; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1572 = 7'h1b == index ? io_from_lsu_wdata : record_wdata1_27; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1573 = 7'h1c == index ? io_from_lsu_wdata : record_wdata1_28; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1574 = 7'h1d == index ? io_from_lsu_wdata : record_wdata1_29; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1575 = 7'h1e == index ? io_from_lsu_wdata : record_wdata1_30; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1576 = 7'h1f == index ? io_from_lsu_wdata : record_wdata1_31; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1577 = 7'h20 == index ? io_from_lsu_wdata : record_wdata1_32; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1578 = 7'h21 == index ? io_from_lsu_wdata : record_wdata1_33; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1579 = 7'h22 == index ? io_from_lsu_wdata : record_wdata1_34; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1580 = 7'h23 == index ? io_from_lsu_wdata : record_wdata1_35; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1581 = 7'h24 == index ? io_from_lsu_wdata : record_wdata1_36; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1582 = 7'h25 == index ? io_from_lsu_wdata : record_wdata1_37; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1583 = 7'h26 == index ? io_from_lsu_wdata : record_wdata1_38; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1584 = 7'h27 == index ? io_from_lsu_wdata : record_wdata1_39; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1585 = 7'h28 == index ? io_from_lsu_wdata : record_wdata1_40; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1586 = 7'h29 == index ? io_from_lsu_wdata : record_wdata1_41; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1587 = 7'h2a == index ? io_from_lsu_wdata : record_wdata1_42; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1588 = 7'h2b == index ? io_from_lsu_wdata : record_wdata1_43; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1589 = 7'h2c == index ? io_from_lsu_wdata : record_wdata1_44; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1590 = 7'h2d == index ? io_from_lsu_wdata : record_wdata1_45; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1591 = 7'h2e == index ? io_from_lsu_wdata : record_wdata1_46; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1592 = 7'h2f == index ? io_from_lsu_wdata : record_wdata1_47; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1593 = 7'h30 == index ? io_from_lsu_wdata : record_wdata1_48; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1594 = 7'h31 == index ? io_from_lsu_wdata : record_wdata1_49; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1595 = 7'h32 == index ? io_from_lsu_wdata : record_wdata1_50; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1596 = 7'h33 == index ? io_from_lsu_wdata : record_wdata1_51; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1597 = 7'h34 == index ? io_from_lsu_wdata : record_wdata1_52; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1598 = 7'h35 == index ? io_from_lsu_wdata : record_wdata1_53; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1599 = 7'h36 == index ? io_from_lsu_wdata : record_wdata1_54; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1600 = 7'h37 == index ? io_from_lsu_wdata : record_wdata1_55; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1601 = 7'h38 == index ? io_from_lsu_wdata : record_wdata1_56; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1602 = 7'h39 == index ? io_from_lsu_wdata : record_wdata1_57; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1603 = 7'h3a == index ? io_from_lsu_wdata : record_wdata1_58; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1604 = 7'h3b == index ? io_from_lsu_wdata : record_wdata1_59; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1605 = 7'h3c == index ? io_from_lsu_wdata : record_wdata1_60; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1606 = 7'h3d == index ? io_from_lsu_wdata : record_wdata1_61; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1607 = 7'h3e == index ? io_from_lsu_wdata : record_wdata1_62; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1608 = 7'h3f == index ? io_from_lsu_wdata : record_wdata1_63; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1609 = 7'h40 == index ? io_from_lsu_wdata : record_wdata1_64; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1610 = 7'h41 == index ? io_from_lsu_wdata : record_wdata1_65; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1611 = 7'h42 == index ? io_from_lsu_wdata : record_wdata1_66; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1612 = 7'h43 == index ? io_from_lsu_wdata : record_wdata1_67; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1613 = 7'h44 == index ? io_from_lsu_wdata : record_wdata1_68; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1614 = 7'h45 == index ? io_from_lsu_wdata : record_wdata1_69; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1615 = 7'h46 == index ? io_from_lsu_wdata : record_wdata1_70; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1616 = 7'h47 == index ? io_from_lsu_wdata : record_wdata1_71; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1617 = 7'h48 == index ? io_from_lsu_wdata : record_wdata1_72; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1618 = 7'h49 == index ? io_from_lsu_wdata : record_wdata1_73; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1619 = 7'h4a == index ? io_from_lsu_wdata : record_wdata1_74; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1620 = 7'h4b == index ? io_from_lsu_wdata : record_wdata1_75; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1621 = 7'h4c == index ? io_from_lsu_wdata : record_wdata1_76; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1622 = 7'h4d == index ? io_from_lsu_wdata : record_wdata1_77; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1623 = 7'h4e == index ? io_from_lsu_wdata : record_wdata1_78; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1624 = 7'h4f == index ? io_from_lsu_wdata : record_wdata1_79; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1625 = 7'h50 == index ? io_from_lsu_wdata : record_wdata1_80; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1626 = 7'h51 == index ? io_from_lsu_wdata : record_wdata1_81; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1627 = 7'h52 == index ? io_from_lsu_wdata : record_wdata1_82; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1628 = 7'h53 == index ? io_from_lsu_wdata : record_wdata1_83; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1629 = 7'h54 == index ? io_from_lsu_wdata : record_wdata1_84; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1630 = 7'h55 == index ? io_from_lsu_wdata : record_wdata1_85; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1631 = 7'h56 == index ? io_from_lsu_wdata : record_wdata1_86; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1632 = 7'h57 == index ? io_from_lsu_wdata : record_wdata1_87; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1633 = 7'h58 == index ? io_from_lsu_wdata : record_wdata1_88; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1634 = 7'h59 == index ? io_from_lsu_wdata : record_wdata1_89; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1635 = 7'h5a == index ? io_from_lsu_wdata : record_wdata1_90; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1636 = 7'h5b == index ? io_from_lsu_wdata : record_wdata1_91; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1637 = 7'h5c == index ? io_from_lsu_wdata : record_wdata1_92; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1638 = 7'h5d == index ? io_from_lsu_wdata : record_wdata1_93; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1639 = 7'h5e == index ? io_from_lsu_wdata : record_wdata1_94; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1640 = 7'h5f == index ? io_from_lsu_wdata : record_wdata1_95; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1641 = 7'h60 == index ? io_from_lsu_wdata : record_wdata1_96; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1642 = 7'h61 == index ? io_from_lsu_wdata : record_wdata1_97; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1643 = 7'h62 == index ? io_from_lsu_wdata : record_wdata1_98; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1644 = 7'h63 == index ? io_from_lsu_wdata : record_wdata1_99; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1645 = 7'h64 == index ? io_from_lsu_wdata : record_wdata1_100; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1646 = 7'h65 == index ? io_from_lsu_wdata : record_wdata1_101; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1647 = 7'h66 == index ? io_from_lsu_wdata : record_wdata1_102; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1648 = 7'h67 == index ? io_from_lsu_wdata : record_wdata1_103; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1649 = 7'h68 == index ? io_from_lsu_wdata : record_wdata1_104; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1650 = 7'h69 == index ? io_from_lsu_wdata : record_wdata1_105; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1651 = 7'h6a == index ? io_from_lsu_wdata : record_wdata1_106; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1652 = 7'h6b == index ? io_from_lsu_wdata : record_wdata1_107; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1653 = 7'h6c == index ? io_from_lsu_wdata : record_wdata1_108; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1654 = 7'h6d == index ? io_from_lsu_wdata : record_wdata1_109; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1655 = 7'h6e == index ? io_from_lsu_wdata : record_wdata1_110; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1656 = 7'h6f == index ? io_from_lsu_wdata : record_wdata1_111; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1657 = 7'h70 == index ? io_from_lsu_wdata : record_wdata1_112; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1658 = 7'h71 == index ? io_from_lsu_wdata : record_wdata1_113; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1659 = 7'h72 == index ? io_from_lsu_wdata : record_wdata1_114; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1660 = 7'h73 == index ? io_from_lsu_wdata : record_wdata1_115; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1661 = 7'h74 == index ? io_from_lsu_wdata : record_wdata1_116; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1662 = 7'h75 == index ? io_from_lsu_wdata : record_wdata1_117; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1663 = 7'h76 == index ? io_from_lsu_wdata : record_wdata1_118; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1664 = 7'h77 == index ? io_from_lsu_wdata : record_wdata1_119; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1665 = 7'h78 == index ? io_from_lsu_wdata : record_wdata1_120; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1666 = 7'h79 == index ? io_from_lsu_wdata : record_wdata1_121; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1667 = 7'h7a == index ? io_from_lsu_wdata : record_wdata1_122; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1668 = 7'h7b == index ? io_from_lsu_wdata : record_wdata1_123; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1669 = 7'h7c == index ? io_from_lsu_wdata : record_wdata1_124; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1670 = 7'h7d == index ? io_from_lsu_wdata : record_wdata1_125; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1671 = 7'h7e == index ? io_from_lsu_wdata : record_wdata1_126; // @[d_cache.scala 125:{38,38} 21:32]
  wire [63:0] _GEN_1672 = 7'h7f == index ? io_from_lsu_wdata : record_wdata1_127; // @[d_cache.scala 125:{38,38} 21:32]
  wire [7:0] _GEN_1673 = 7'h0 == index ? io_from_lsu_wstrb : record_wstrb1_0; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1674 = 7'h1 == index ? io_from_lsu_wstrb : record_wstrb1_1; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1675 = 7'h2 == index ? io_from_lsu_wstrb : record_wstrb1_2; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1676 = 7'h3 == index ? io_from_lsu_wstrb : record_wstrb1_3; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1677 = 7'h4 == index ? io_from_lsu_wstrb : record_wstrb1_4; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1678 = 7'h5 == index ? io_from_lsu_wstrb : record_wstrb1_5; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1679 = 7'h6 == index ? io_from_lsu_wstrb : record_wstrb1_6; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1680 = 7'h7 == index ? io_from_lsu_wstrb : record_wstrb1_7; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1681 = 7'h8 == index ? io_from_lsu_wstrb : record_wstrb1_8; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1682 = 7'h9 == index ? io_from_lsu_wstrb : record_wstrb1_9; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1683 = 7'ha == index ? io_from_lsu_wstrb : record_wstrb1_10; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1684 = 7'hb == index ? io_from_lsu_wstrb : record_wstrb1_11; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1685 = 7'hc == index ? io_from_lsu_wstrb : record_wstrb1_12; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1686 = 7'hd == index ? io_from_lsu_wstrb : record_wstrb1_13; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1687 = 7'he == index ? io_from_lsu_wstrb : record_wstrb1_14; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1688 = 7'hf == index ? io_from_lsu_wstrb : record_wstrb1_15; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1689 = 7'h10 == index ? io_from_lsu_wstrb : record_wstrb1_16; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1690 = 7'h11 == index ? io_from_lsu_wstrb : record_wstrb1_17; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1691 = 7'h12 == index ? io_from_lsu_wstrb : record_wstrb1_18; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1692 = 7'h13 == index ? io_from_lsu_wstrb : record_wstrb1_19; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1693 = 7'h14 == index ? io_from_lsu_wstrb : record_wstrb1_20; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1694 = 7'h15 == index ? io_from_lsu_wstrb : record_wstrb1_21; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1695 = 7'h16 == index ? io_from_lsu_wstrb : record_wstrb1_22; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1696 = 7'h17 == index ? io_from_lsu_wstrb : record_wstrb1_23; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1697 = 7'h18 == index ? io_from_lsu_wstrb : record_wstrb1_24; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1698 = 7'h19 == index ? io_from_lsu_wstrb : record_wstrb1_25; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1699 = 7'h1a == index ? io_from_lsu_wstrb : record_wstrb1_26; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1700 = 7'h1b == index ? io_from_lsu_wstrb : record_wstrb1_27; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1701 = 7'h1c == index ? io_from_lsu_wstrb : record_wstrb1_28; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1702 = 7'h1d == index ? io_from_lsu_wstrb : record_wstrb1_29; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1703 = 7'h1e == index ? io_from_lsu_wstrb : record_wstrb1_30; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1704 = 7'h1f == index ? io_from_lsu_wstrb : record_wstrb1_31; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1705 = 7'h20 == index ? io_from_lsu_wstrb : record_wstrb1_32; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1706 = 7'h21 == index ? io_from_lsu_wstrb : record_wstrb1_33; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1707 = 7'h22 == index ? io_from_lsu_wstrb : record_wstrb1_34; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1708 = 7'h23 == index ? io_from_lsu_wstrb : record_wstrb1_35; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1709 = 7'h24 == index ? io_from_lsu_wstrb : record_wstrb1_36; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1710 = 7'h25 == index ? io_from_lsu_wstrb : record_wstrb1_37; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1711 = 7'h26 == index ? io_from_lsu_wstrb : record_wstrb1_38; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1712 = 7'h27 == index ? io_from_lsu_wstrb : record_wstrb1_39; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1713 = 7'h28 == index ? io_from_lsu_wstrb : record_wstrb1_40; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1714 = 7'h29 == index ? io_from_lsu_wstrb : record_wstrb1_41; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1715 = 7'h2a == index ? io_from_lsu_wstrb : record_wstrb1_42; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1716 = 7'h2b == index ? io_from_lsu_wstrb : record_wstrb1_43; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1717 = 7'h2c == index ? io_from_lsu_wstrb : record_wstrb1_44; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1718 = 7'h2d == index ? io_from_lsu_wstrb : record_wstrb1_45; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1719 = 7'h2e == index ? io_from_lsu_wstrb : record_wstrb1_46; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1720 = 7'h2f == index ? io_from_lsu_wstrb : record_wstrb1_47; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1721 = 7'h30 == index ? io_from_lsu_wstrb : record_wstrb1_48; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1722 = 7'h31 == index ? io_from_lsu_wstrb : record_wstrb1_49; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1723 = 7'h32 == index ? io_from_lsu_wstrb : record_wstrb1_50; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1724 = 7'h33 == index ? io_from_lsu_wstrb : record_wstrb1_51; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1725 = 7'h34 == index ? io_from_lsu_wstrb : record_wstrb1_52; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1726 = 7'h35 == index ? io_from_lsu_wstrb : record_wstrb1_53; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1727 = 7'h36 == index ? io_from_lsu_wstrb : record_wstrb1_54; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1728 = 7'h37 == index ? io_from_lsu_wstrb : record_wstrb1_55; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1729 = 7'h38 == index ? io_from_lsu_wstrb : record_wstrb1_56; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1730 = 7'h39 == index ? io_from_lsu_wstrb : record_wstrb1_57; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1731 = 7'h3a == index ? io_from_lsu_wstrb : record_wstrb1_58; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1732 = 7'h3b == index ? io_from_lsu_wstrb : record_wstrb1_59; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1733 = 7'h3c == index ? io_from_lsu_wstrb : record_wstrb1_60; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1734 = 7'h3d == index ? io_from_lsu_wstrb : record_wstrb1_61; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1735 = 7'h3e == index ? io_from_lsu_wstrb : record_wstrb1_62; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1736 = 7'h3f == index ? io_from_lsu_wstrb : record_wstrb1_63; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1737 = 7'h40 == index ? io_from_lsu_wstrb : record_wstrb1_64; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1738 = 7'h41 == index ? io_from_lsu_wstrb : record_wstrb1_65; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1739 = 7'h42 == index ? io_from_lsu_wstrb : record_wstrb1_66; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1740 = 7'h43 == index ? io_from_lsu_wstrb : record_wstrb1_67; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1741 = 7'h44 == index ? io_from_lsu_wstrb : record_wstrb1_68; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1742 = 7'h45 == index ? io_from_lsu_wstrb : record_wstrb1_69; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1743 = 7'h46 == index ? io_from_lsu_wstrb : record_wstrb1_70; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1744 = 7'h47 == index ? io_from_lsu_wstrb : record_wstrb1_71; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1745 = 7'h48 == index ? io_from_lsu_wstrb : record_wstrb1_72; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1746 = 7'h49 == index ? io_from_lsu_wstrb : record_wstrb1_73; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1747 = 7'h4a == index ? io_from_lsu_wstrb : record_wstrb1_74; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1748 = 7'h4b == index ? io_from_lsu_wstrb : record_wstrb1_75; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1749 = 7'h4c == index ? io_from_lsu_wstrb : record_wstrb1_76; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1750 = 7'h4d == index ? io_from_lsu_wstrb : record_wstrb1_77; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1751 = 7'h4e == index ? io_from_lsu_wstrb : record_wstrb1_78; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1752 = 7'h4f == index ? io_from_lsu_wstrb : record_wstrb1_79; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1753 = 7'h50 == index ? io_from_lsu_wstrb : record_wstrb1_80; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1754 = 7'h51 == index ? io_from_lsu_wstrb : record_wstrb1_81; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1755 = 7'h52 == index ? io_from_lsu_wstrb : record_wstrb1_82; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1756 = 7'h53 == index ? io_from_lsu_wstrb : record_wstrb1_83; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1757 = 7'h54 == index ? io_from_lsu_wstrb : record_wstrb1_84; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1758 = 7'h55 == index ? io_from_lsu_wstrb : record_wstrb1_85; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1759 = 7'h56 == index ? io_from_lsu_wstrb : record_wstrb1_86; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1760 = 7'h57 == index ? io_from_lsu_wstrb : record_wstrb1_87; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1761 = 7'h58 == index ? io_from_lsu_wstrb : record_wstrb1_88; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1762 = 7'h59 == index ? io_from_lsu_wstrb : record_wstrb1_89; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1763 = 7'h5a == index ? io_from_lsu_wstrb : record_wstrb1_90; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1764 = 7'h5b == index ? io_from_lsu_wstrb : record_wstrb1_91; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1765 = 7'h5c == index ? io_from_lsu_wstrb : record_wstrb1_92; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1766 = 7'h5d == index ? io_from_lsu_wstrb : record_wstrb1_93; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1767 = 7'h5e == index ? io_from_lsu_wstrb : record_wstrb1_94; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1768 = 7'h5f == index ? io_from_lsu_wstrb : record_wstrb1_95; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1769 = 7'h60 == index ? io_from_lsu_wstrb : record_wstrb1_96; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1770 = 7'h61 == index ? io_from_lsu_wstrb : record_wstrb1_97; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1771 = 7'h62 == index ? io_from_lsu_wstrb : record_wstrb1_98; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1772 = 7'h63 == index ? io_from_lsu_wstrb : record_wstrb1_99; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1773 = 7'h64 == index ? io_from_lsu_wstrb : record_wstrb1_100; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1774 = 7'h65 == index ? io_from_lsu_wstrb : record_wstrb1_101; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1775 = 7'h66 == index ? io_from_lsu_wstrb : record_wstrb1_102; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1776 = 7'h67 == index ? io_from_lsu_wstrb : record_wstrb1_103; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1777 = 7'h68 == index ? io_from_lsu_wstrb : record_wstrb1_104; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1778 = 7'h69 == index ? io_from_lsu_wstrb : record_wstrb1_105; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1779 = 7'h6a == index ? io_from_lsu_wstrb : record_wstrb1_106; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1780 = 7'h6b == index ? io_from_lsu_wstrb : record_wstrb1_107; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1781 = 7'h6c == index ? io_from_lsu_wstrb : record_wstrb1_108; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1782 = 7'h6d == index ? io_from_lsu_wstrb : record_wstrb1_109; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1783 = 7'h6e == index ? io_from_lsu_wstrb : record_wstrb1_110; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1784 = 7'h6f == index ? io_from_lsu_wstrb : record_wstrb1_111; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1785 = 7'h70 == index ? io_from_lsu_wstrb : record_wstrb1_112; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1786 = 7'h71 == index ? io_from_lsu_wstrb : record_wstrb1_113; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1787 = 7'h72 == index ? io_from_lsu_wstrb : record_wstrb1_114; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1788 = 7'h73 == index ? io_from_lsu_wstrb : record_wstrb1_115; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1789 = 7'h74 == index ? io_from_lsu_wstrb : record_wstrb1_116; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1790 = 7'h75 == index ? io_from_lsu_wstrb : record_wstrb1_117; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1791 = 7'h76 == index ? io_from_lsu_wstrb : record_wstrb1_118; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1792 = 7'h77 == index ? io_from_lsu_wstrb : record_wstrb1_119; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1793 = 7'h78 == index ? io_from_lsu_wstrb : record_wstrb1_120; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1794 = 7'h79 == index ? io_from_lsu_wstrb : record_wstrb1_121; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1795 = 7'h7a == index ? io_from_lsu_wstrb : record_wstrb1_122; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1796 = 7'h7b == index ? io_from_lsu_wstrb : record_wstrb1_123; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1797 = 7'h7c == index ? io_from_lsu_wstrb : record_wstrb1_124; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1798 = 7'h7d == index ? io_from_lsu_wstrb : record_wstrb1_125; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1799 = 7'h7e == index ? io_from_lsu_wstrb : record_wstrb1_126; // @[d_cache.scala 126:{38,38} 22:32]
  wire [7:0] _GEN_1800 = 7'h7f == index ? io_from_lsu_wstrb : record_wstrb1_127; // @[d_cache.scala 126:{38,38} 22:32]
  wire [63:0] _GEN_1801 = 7'h0 == index ? io_pc_now : record_pc_0; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1802 = 7'h1 == index ? io_pc_now : record_pc_1; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1803 = 7'h2 == index ? io_pc_now : record_pc_2; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1804 = 7'h3 == index ? io_pc_now : record_pc_3; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1805 = 7'h4 == index ? io_pc_now : record_pc_4; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1806 = 7'h5 == index ? io_pc_now : record_pc_5; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1807 = 7'h6 == index ? io_pc_now : record_pc_6; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1808 = 7'h7 == index ? io_pc_now : record_pc_7; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1809 = 7'h8 == index ? io_pc_now : record_pc_8; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1810 = 7'h9 == index ? io_pc_now : record_pc_9; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1811 = 7'ha == index ? io_pc_now : record_pc_10; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1812 = 7'hb == index ? io_pc_now : record_pc_11; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1813 = 7'hc == index ? io_pc_now : record_pc_12; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1814 = 7'hd == index ? io_pc_now : record_pc_13; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1815 = 7'he == index ? io_pc_now : record_pc_14; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1816 = 7'hf == index ? io_pc_now : record_pc_15; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1817 = 7'h10 == index ? io_pc_now : record_pc_16; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1818 = 7'h11 == index ? io_pc_now : record_pc_17; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1819 = 7'h12 == index ? io_pc_now : record_pc_18; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1820 = 7'h13 == index ? io_pc_now : record_pc_19; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1821 = 7'h14 == index ? io_pc_now : record_pc_20; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1822 = 7'h15 == index ? io_pc_now : record_pc_21; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1823 = 7'h16 == index ? io_pc_now : record_pc_22; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1824 = 7'h17 == index ? io_pc_now : record_pc_23; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1825 = 7'h18 == index ? io_pc_now : record_pc_24; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1826 = 7'h19 == index ? io_pc_now : record_pc_25; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1827 = 7'h1a == index ? io_pc_now : record_pc_26; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1828 = 7'h1b == index ? io_pc_now : record_pc_27; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1829 = 7'h1c == index ? io_pc_now : record_pc_28; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1830 = 7'h1d == index ? io_pc_now : record_pc_29; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1831 = 7'h1e == index ? io_pc_now : record_pc_30; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1832 = 7'h1f == index ? io_pc_now : record_pc_31; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1833 = 7'h20 == index ? io_pc_now : record_pc_32; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1834 = 7'h21 == index ? io_pc_now : record_pc_33; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1835 = 7'h22 == index ? io_pc_now : record_pc_34; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1836 = 7'h23 == index ? io_pc_now : record_pc_35; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1837 = 7'h24 == index ? io_pc_now : record_pc_36; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1838 = 7'h25 == index ? io_pc_now : record_pc_37; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1839 = 7'h26 == index ? io_pc_now : record_pc_38; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1840 = 7'h27 == index ? io_pc_now : record_pc_39; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1841 = 7'h28 == index ? io_pc_now : record_pc_40; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1842 = 7'h29 == index ? io_pc_now : record_pc_41; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1843 = 7'h2a == index ? io_pc_now : record_pc_42; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1844 = 7'h2b == index ? io_pc_now : record_pc_43; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1845 = 7'h2c == index ? io_pc_now : record_pc_44; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1846 = 7'h2d == index ? io_pc_now : record_pc_45; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1847 = 7'h2e == index ? io_pc_now : record_pc_46; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1848 = 7'h2f == index ? io_pc_now : record_pc_47; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1849 = 7'h30 == index ? io_pc_now : record_pc_48; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1850 = 7'h31 == index ? io_pc_now : record_pc_49; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1851 = 7'h32 == index ? io_pc_now : record_pc_50; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1852 = 7'h33 == index ? io_pc_now : record_pc_51; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1853 = 7'h34 == index ? io_pc_now : record_pc_52; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1854 = 7'h35 == index ? io_pc_now : record_pc_53; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1855 = 7'h36 == index ? io_pc_now : record_pc_54; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1856 = 7'h37 == index ? io_pc_now : record_pc_55; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1857 = 7'h38 == index ? io_pc_now : record_pc_56; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1858 = 7'h39 == index ? io_pc_now : record_pc_57; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1859 = 7'h3a == index ? io_pc_now : record_pc_58; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1860 = 7'h3b == index ? io_pc_now : record_pc_59; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1861 = 7'h3c == index ? io_pc_now : record_pc_60; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1862 = 7'h3d == index ? io_pc_now : record_pc_61; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1863 = 7'h3e == index ? io_pc_now : record_pc_62; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1864 = 7'h3f == index ? io_pc_now : record_pc_63; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1865 = 7'h40 == index ? io_pc_now : record_pc_64; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1866 = 7'h41 == index ? io_pc_now : record_pc_65; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1867 = 7'h42 == index ? io_pc_now : record_pc_66; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1868 = 7'h43 == index ? io_pc_now : record_pc_67; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1869 = 7'h44 == index ? io_pc_now : record_pc_68; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1870 = 7'h45 == index ? io_pc_now : record_pc_69; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1871 = 7'h46 == index ? io_pc_now : record_pc_70; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1872 = 7'h47 == index ? io_pc_now : record_pc_71; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1873 = 7'h48 == index ? io_pc_now : record_pc_72; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1874 = 7'h49 == index ? io_pc_now : record_pc_73; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1875 = 7'h4a == index ? io_pc_now : record_pc_74; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1876 = 7'h4b == index ? io_pc_now : record_pc_75; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1877 = 7'h4c == index ? io_pc_now : record_pc_76; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1878 = 7'h4d == index ? io_pc_now : record_pc_77; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1879 = 7'h4e == index ? io_pc_now : record_pc_78; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1880 = 7'h4f == index ? io_pc_now : record_pc_79; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1881 = 7'h50 == index ? io_pc_now : record_pc_80; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1882 = 7'h51 == index ? io_pc_now : record_pc_81; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1883 = 7'h52 == index ? io_pc_now : record_pc_82; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1884 = 7'h53 == index ? io_pc_now : record_pc_83; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1885 = 7'h54 == index ? io_pc_now : record_pc_84; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1886 = 7'h55 == index ? io_pc_now : record_pc_85; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1887 = 7'h56 == index ? io_pc_now : record_pc_86; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1888 = 7'h57 == index ? io_pc_now : record_pc_87; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1889 = 7'h58 == index ? io_pc_now : record_pc_88; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1890 = 7'h59 == index ? io_pc_now : record_pc_89; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1891 = 7'h5a == index ? io_pc_now : record_pc_90; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1892 = 7'h5b == index ? io_pc_now : record_pc_91; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1893 = 7'h5c == index ? io_pc_now : record_pc_92; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1894 = 7'h5d == index ? io_pc_now : record_pc_93; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1895 = 7'h5e == index ? io_pc_now : record_pc_94; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1896 = 7'h5f == index ? io_pc_now : record_pc_95; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1897 = 7'h60 == index ? io_pc_now : record_pc_96; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1898 = 7'h61 == index ? io_pc_now : record_pc_97; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1899 = 7'h62 == index ? io_pc_now : record_pc_98; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1900 = 7'h63 == index ? io_pc_now : record_pc_99; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1901 = 7'h64 == index ? io_pc_now : record_pc_100; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1902 = 7'h65 == index ? io_pc_now : record_pc_101; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1903 = 7'h66 == index ? io_pc_now : record_pc_102; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1904 = 7'h67 == index ? io_pc_now : record_pc_103; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1905 = 7'h68 == index ? io_pc_now : record_pc_104; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1906 = 7'h69 == index ? io_pc_now : record_pc_105; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1907 = 7'h6a == index ? io_pc_now : record_pc_106; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1908 = 7'h6b == index ? io_pc_now : record_pc_107; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1909 = 7'h6c == index ? io_pc_now : record_pc_108; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1910 = 7'h6d == index ? io_pc_now : record_pc_109; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1911 = 7'h6e == index ? io_pc_now : record_pc_110; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1912 = 7'h6f == index ? io_pc_now : record_pc_111; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1913 = 7'h70 == index ? io_pc_now : record_pc_112; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1914 = 7'h71 == index ? io_pc_now : record_pc_113; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1915 = 7'h72 == index ? io_pc_now : record_pc_114; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1916 = 7'h73 == index ? io_pc_now : record_pc_115; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1917 = 7'h74 == index ? io_pc_now : record_pc_116; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1918 = 7'h75 == index ? io_pc_now : record_pc_117; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1919 = 7'h76 == index ? io_pc_now : record_pc_118; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1920 = 7'h77 == index ? io_pc_now : record_pc_119; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1921 = 7'h78 == index ? io_pc_now : record_pc_120; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1922 = 7'h79 == index ? io_pc_now : record_pc_121; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1923 = 7'h7a == index ? io_pc_now : record_pc_122; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1924 = 7'h7b == index ? io_pc_now : record_pc_123; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1925 = 7'h7c == index ? io_pc_now : record_pc_124; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1926 = 7'h7d == index ? io_pc_now : record_pc_125; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1927 = 7'h7e == index ? io_pc_now : record_pc_126; // @[d_cache.scala 127:{34,34} 23:28]
  wire [63:0] _GEN_1928 = 7'h7f == index ? io_pc_now : record_pc_127; // @[d_cache.scala 127:{34,34} 23:28]
  wire [31:0] _GEN_1929 = 7'h0 == index ? io_from_lsu_awaddr : record_addr_0; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1930 = 7'h1 == index ? io_from_lsu_awaddr : record_addr_1; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1931 = 7'h2 == index ? io_from_lsu_awaddr : record_addr_2; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1932 = 7'h3 == index ? io_from_lsu_awaddr : record_addr_3; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1933 = 7'h4 == index ? io_from_lsu_awaddr : record_addr_4; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1934 = 7'h5 == index ? io_from_lsu_awaddr : record_addr_5; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1935 = 7'h6 == index ? io_from_lsu_awaddr : record_addr_6; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1936 = 7'h7 == index ? io_from_lsu_awaddr : record_addr_7; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1937 = 7'h8 == index ? io_from_lsu_awaddr : record_addr_8; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1938 = 7'h9 == index ? io_from_lsu_awaddr : record_addr_9; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1939 = 7'ha == index ? io_from_lsu_awaddr : record_addr_10; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1940 = 7'hb == index ? io_from_lsu_awaddr : record_addr_11; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1941 = 7'hc == index ? io_from_lsu_awaddr : record_addr_12; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1942 = 7'hd == index ? io_from_lsu_awaddr : record_addr_13; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1943 = 7'he == index ? io_from_lsu_awaddr : record_addr_14; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1944 = 7'hf == index ? io_from_lsu_awaddr : record_addr_15; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1945 = 7'h10 == index ? io_from_lsu_awaddr : record_addr_16; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1946 = 7'h11 == index ? io_from_lsu_awaddr : record_addr_17; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1947 = 7'h12 == index ? io_from_lsu_awaddr : record_addr_18; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1948 = 7'h13 == index ? io_from_lsu_awaddr : record_addr_19; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1949 = 7'h14 == index ? io_from_lsu_awaddr : record_addr_20; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1950 = 7'h15 == index ? io_from_lsu_awaddr : record_addr_21; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1951 = 7'h16 == index ? io_from_lsu_awaddr : record_addr_22; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1952 = 7'h17 == index ? io_from_lsu_awaddr : record_addr_23; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1953 = 7'h18 == index ? io_from_lsu_awaddr : record_addr_24; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1954 = 7'h19 == index ? io_from_lsu_awaddr : record_addr_25; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1955 = 7'h1a == index ? io_from_lsu_awaddr : record_addr_26; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1956 = 7'h1b == index ? io_from_lsu_awaddr : record_addr_27; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1957 = 7'h1c == index ? io_from_lsu_awaddr : record_addr_28; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1958 = 7'h1d == index ? io_from_lsu_awaddr : record_addr_29; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1959 = 7'h1e == index ? io_from_lsu_awaddr : record_addr_30; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1960 = 7'h1f == index ? io_from_lsu_awaddr : record_addr_31; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1961 = 7'h20 == index ? io_from_lsu_awaddr : record_addr_32; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1962 = 7'h21 == index ? io_from_lsu_awaddr : record_addr_33; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1963 = 7'h22 == index ? io_from_lsu_awaddr : record_addr_34; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1964 = 7'h23 == index ? io_from_lsu_awaddr : record_addr_35; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1965 = 7'h24 == index ? io_from_lsu_awaddr : record_addr_36; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1966 = 7'h25 == index ? io_from_lsu_awaddr : record_addr_37; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1967 = 7'h26 == index ? io_from_lsu_awaddr : record_addr_38; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1968 = 7'h27 == index ? io_from_lsu_awaddr : record_addr_39; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1969 = 7'h28 == index ? io_from_lsu_awaddr : record_addr_40; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1970 = 7'h29 == index ? io_from_lsu_awaddr : record_addr_41; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1971 = 7'h2a == index ? io_from_lsu_awaddr : record_addr_42; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1972 = 7'h2b == index ? io_from_lsu_awaddr : record_addr_43; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1973 = 7'h2c == index ? io_from_lsu_awaddr : record_addr_44; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1974 = 7'h2d == index ? io_from_lsu_awaddr : record_addr_45; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1975 = 7'h2e == index ? io_from_lsu_awaddr : record_addr_46; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1976 = 7'h2f == index ? io_from_lsu_awaddr : record_addr_47; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1977 = 7'h30 == index ? io_from_lsu_awaddr : record_addr_48; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1978 = 7'h31 == index ? io_from_lsu_awaddr : record_addr_49; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1979 = 7'h32 == index ? io_from_lsu_awaddr : record_addr_50; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1980 = 7'h33 == index ? io_from_lsu_awaddr : record_addr_51; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1981 = 7'h34 == index ? io_from_lsu_awaddr : record_addr_52; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1982 = 7'h35 == index ? io_from_lsu_awaddr : record_addr_53; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1983 = 7'h36 == index ? io_from_lsu_awaddr : record_addr_54; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1984 = 7'h37 == index ? io_from_lsu_awaddr : record_addr_55; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1985 = 7'h38 == index ? io_from_lsu_awaddr : record_addr_56; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1986 = 7'h39 == index ? io_from_lsu_awaddr : record_addr_57; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1987 = 7'h3a == index ? io_from_lsu_awaddr : record_addr_58; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1988 = 7'h3b == index ? io_from_lsu_awaddr : record_addr_59; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1989 = 7'h3c == index ? io_from_lsu_awaddr : record_addr_60; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1990 = 7'h3d == index ? io_from_lsu_awaddr : record_addr_61; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1991 = 7'h3e == index ? io_from_lsu_awaddr : record_addr_62; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1992 = 7'h3f == index ? io_from_lsu_awaddr : record_addr_63; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1993 = 7'h40 == index ? io_from_lsu_awaddr : record_addr_64; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1994 = 7'h41 == index ? io_from_lsu_awaddr : record_addr_65; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1995 = 7'h42 == index ? io_from_lsu_awaddr : record_addr_66; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1996 = 7'h43 == index ? io_from_lsu_awaddr : record_addr_67; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1997 = 7'h44 == index ? io_from_lsu_awaddr : record_addr_68; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1998 = 7'h45 == index ? io_from_lsu_awaddr : record_addr_69; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_1999 = 7'h46 == index ? io_from_lsu_awaddr : record_addr_70; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2000 = 7'h47 == index ? io_from_lsu_awaddr : record_addr_71; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2001 = 7'h48 == index ? io_from_lsu_awaddr : record_addr_72; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2002 = 7'h49 == index ? io_from_lsu_awaddr : record_addr_73; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2003 = 7'h4a == index ? io_from_lsu_awaddr : record_addr_74; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2004 = 7'h4b == index ? io_from_lsu_awaddr : record_addr_75; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2005 = 7'h4c == index ? io_from_lsu_awaddr : record_addr_76; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2006 = 7'h4d == index ? io_from_lsu_awaddr : record_addr_77; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2007 = 7'h4e == index ? io_from_lsu_awaddr : record_addr_78; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2008 = 7'h4f == index ? io_from_lsu_awaddr : record_addr_79; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2009 = 7'h50 == index ? io_from_lsu_awaddr : record_addr_80; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2010 = 7'h51 == index ? io_from_lsu_awaddr : record_addr_81; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2011 = 7'h52 == index ? io_from_lsu_awaddr : record_addr_82; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2012 = 7'h53 == index ? io_from_lsu_awaddr : record_addr_83; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2013 = 7'h54 == index ? io_from_lsu_awaddr : record_addr_84; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2014 = 7'h55 == index ? io_from_lsu_awaddr : record_addr_85; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2015 = 7'h56 == index ? io_from_lsu_awaddr : record_addr_86; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2016 = 7'h57 == index ? io_from_lsu_awaddr : record_addr_87; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2017 = 7'h58 == index ? io_from_lsu_awaddr : record_addr_88; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2018 = 7'h59 == index ? io_from_lsu_awaddr : record_addr_89; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2019 = 7'h5a == index ? io_from_lsu_awaddr : record_addr_90; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2020 = 7'h5b == index ? io_from_lsu_awaddr : record_addr_91; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2021 = 7'h5c == index ? io_from_lsu_awaddr : record_addr_92; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2022 = 7'h5d == index ? io_from_lsu_awaddr : record_addr_93; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2023 = 7'h5e == index ? io_from_lsu_awaddr : record_addr_94; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2024 = 7'h5f == index ? io_from_lsu_awaddr : record_addr_95; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2025 = 7'h60 == index ? io_from_lsu_awaddr : record_addr_96; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2026 = 7'h61 == index ? io_from_lsu_awaddr : record_addr_97; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2027 = 7'h62 == index ? io_from_lsu_awaddr : record_addr_98; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2028 = 7'h63 == index ? io_from_lsu_awaddr : record_addr_99; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2029 = 7'h64 == index ? io_from_lsu_awaddr : record_addr_100; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2030 = 7'h65 == index ? io_from_lsu_awaddr : record_addr_101; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2031 = 7'h66 == index ? io_from_lsu_awaddr : record_addr_102; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2032 = 7'h67 == index ? io_from_lsu_awaddr : record_addr_103; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2033 = 7'h68 == index ? io_from_lsu_awaddr : record_addr_104; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2034 = 7'h69 == index ? io_from_lsu_awaddr : record_addr_105; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2035 = 7'h6a == index ? io_from_lsu_awaddr : record_addr_106; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2036 = 7'h6b == index ? io_from_lsu_awaddr : record_addr_107; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2037 = 7'h6c == index ? io_from_lsu_awaddr : record_addr_108; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2038 = 7'h6d == index ? io_from_lsu_awaddr : record_addr_109; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2039 = 7'h6e == index ? io_from_lsu_awaddr : record_addr_110; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2040 = 7'h6f == index ? io_from_lsu_awaddr : record_addr_111; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2041 = 7'h70 == index ? io_from_lsu_awaddr : record_addr_112; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2042 = 7'h71 == index ? io_from_lsu_awaddr : record_addr_113; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2043 = 7'h72 == index ? io_from_lsu_awaddr : record_addr_114; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2044 = 7'h73 == index ? io_from_lsu_awaddr : record_addr_115; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2045 = 7'h74 == index ? io_from_lsu_awaddr : record_addr_116; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2046 = 7'h75 == index ? io_from_lsu_awaddr : record_addr_117; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2047 = 7'h76 == index ? io_from_lsu_awaddr : record_addr_118; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2048 = 7'h77 == index ? io_from_lsu_awaddr : record_addr_119; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2049 = 7'h78 == index ? io_from_lsu_awaddr : record_addr_120; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2050 = 7'h79 == index ? io_from_lsu_awaddr : record_addr_121; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2051 = 7'h7a == index ? io_from_lsu_awaddr : record_addr_122; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2052 = 7'h7b == index ? io_from_lsu_awaddr : record_addr_123; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2053 = 7'h7c == index ? io_from_lsu_awaddr : record_addr_124; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2054 = 7'h7d == index ? io_from_lsu_awaddr : record_addr_125; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2055 = 7'h7e == index ? io_from_lsu_awaddr : record_addr_126; // @[d_cache.scala 128:{36,36} 24:30]
  wire [31:0] _GEN_2056 = 7'h7f == index ? io_from_lsu_awaddr : record_addr_127; // @[d_cache.scala 128:{36,36} 24:30]
  wire  _GEN_2057 = _GEN_19748 | dirty_1_0; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2058 = _GEN_19749 | dirty_1_1; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2059 = _GEN_19750 | dirty_1_2; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2060 = _GEN_19751 | dirty_1_3; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2061 = _GEN_19752 | dirty_1_4; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2062 = _GEN_19753 | dirty_1_5; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2063 = _GEN_19754 | dirty_1_6; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2064 = _GEN_19755 | dirty_1_7; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2065 = _GEN_19756 | dirty_1_8; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2066 = _GEN_19757 | dirty_1_9; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2067 = _GEN_19758 | dirty_1_10; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2068 = _GEN_19759 | dirty_1_11; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2069 = _GEN_19760 | dirty_1_12; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2070 = _GEN_19761 | dirty_1_13; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2071 = _GEN_19762 | dirty_1_14; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2072 = _GEN_19763 | dirty_1_15; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2073 = _GEN_19764 | dirty_1_16; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2074 = _GEN_19765 | dirty_1_17; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2075 = _GEN_19766 | dirty_1_18; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2076 = _GEN_19767 | dirty_1_19; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2077 = _GEN_19768 | dirty_1_20; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2078 = _GEN_19769 | dirty_1_21; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2079 = _GEN_19770 | dirty_1_22; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2080 = _GEN_19771 | dirty_1_23; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2081 = _GEN_19772 | dirty_1_24; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2082 = _GEN_19773 | dirty_1_25; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2083 = _GEN_19774 | dirty_1_26; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2084 = _GEN_19775 | dirty_1_27; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2085 = _GEN_19776 | dirty_1_28; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2086 = _GEN_19777 | dirty_1_29; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2087 = _GEN_19778 | dirty_1_30; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2088 = _GEN_19779 | dirty_1_31; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2089 = _GEN_19780 | dirty_1_32; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2090 = _GEN_19781 | dirty_1_33; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2091 = _GEN_19782 | dirty_1_34; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2092 = _GEN_19783 | dirty_1_35; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2093 = _GEN_19784 | dirty_1_36; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2094 = _GEN_19785 | dirty_1_37; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2095 = _GEN_19786 | dirty_1_38; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2096 = _GEN_19787 | dirty_1_39; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2097 = _GEN_19788 | dirty_1_40; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2098 = _GEN_19789 | dirty_1_41; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2099 = _GEN_19790 | dirty_1_42; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2100 = _GEN_19791 | dirty_1_43; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2101 = _GEN_19792 | dirty_1_44; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2102 = _GEN_19793 | dirty_1_45; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2103 = _GEN_19794 | dirty_1_46; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2104 = _GEN_19795 | dirty_1_47; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2105 = _GEN_19796 | dirty_1_48; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2106 = _GEN_19797 | dirty_1_49; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2107 = _GEN_19798 | dirty_1_50; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2108 = _GEN_19799 | dirty_1_51; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2109 = _GEN_19800 | dirty_1_52; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2110 = _GEN_19801 | dirty_1_53; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2111 = _GEN_19802 | dirty_1_54; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2112 = _GEN_19803 | dirty_1_55; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2113 = _GEN_19804 | dirty_1_56; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2114 = _GEN_19805 | dirty_1_57; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2115 = _GEN_19806 | dirty_1_58; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2116 = _GEN_19807 | dirty_1_59; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2117 = _GEN_19808 | dirty_1_60; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2118 = _GEN_19809 | dirty_1_61; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2119 = _GEN_19810 | dirty_1_62; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2120 = _GEN_19811 | dirty_1_63; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2121 = _GEN_19812 | dirty_1_64; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2122 = _GEN_19813 | dirty_1_65; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2123 = _GEN_19814 | dirty_1_66; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2124 = _GEN_19815 | dirty_1_67; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2125 = _GEN_19816 | dirty_1_68; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2126 = _GEN_19817 | dirty_1_69; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2127 = _GEN_19818 | dirty_1_70; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2128 = _GEN_19819 | dirty_1_71; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2129 = _GEN_19820 | dirty_1_72; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2130 = _GEN_19821 | dirty_1_73; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2131 = _GEN_19822 | dirty_1_74; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2132 = _GEN_19823 | dirty_1_75; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2133 = _GEN_19824 | dirty_1_76; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2134 = _GEN_19825 | dirty_1_77; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2135 = _GEN_19826 | dirty_1_78; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2136 = _GEN_19827 | dirty_1_79; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2137 = _GEN_19828 | dirty_1_80; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2138 = _GEN_19829 | dirty_1_81; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2139 = _GEN_19830 | dirty_1_82; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2140 = _GEN_19831 | dirty_1_83; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2141 = _GEN_19832 | dirty_1_84; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2142 = _GEN_19833 | dirty_1_85; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2143 = _GEN_19834 | dirty_1_86; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2144 = _GEN_19835 | dirty_1_87; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2145 = _GEN_19836 | dirty_1_88; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2146 = _GEN_19837 | dirty_1_89; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2147 = _GEN_19838 | dirty_1_90; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2148 = _GEN_19839 | dirty_1_91; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2149 = _GEN_19840 | dirty_1_92; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2150 = _GEN_19841 | dirty_1_93; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2151 = _GEN_19842 | dirty_1_94; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2152 = _GEN_19843 | dirty_1_95; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2153 = _GEN_19844 | dirty_1_96; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2154 = _GEN_19845 | dirty_1_97; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2155 = _GEN_19846 | dirty_1_98; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2156 = _GEN_19847 | dirty_1_99; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2157 = _GEN_19848 | dirty_1_100; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2158 = _GEN_19849 | dirty_1_101; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2159 = _GEN_19850 | dirty_1_102; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2160 = _GEN_19851 | dirty_1_103; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2161 = _GEN_19852 | dirty_1_104; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2162 = _GEN_19853 | dirty_1_105; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2163 = _GEN_19854 | dirty_1_106; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2164 = _GEN_19855 | dirty_1_107; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2165 = _GEN_19856 | dirty_1_108; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2166 = _GEN_19857 | dirty_1_109; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2167 = _GEN_19858 | dirty_1_110; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2168 = _GEN_19859 | dirty_1_111; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2169 = _GEN_19860 | dirty_1_112; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2170 = _GEN_19861 | dirty_1_113; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2171 = _GEN_19862 | dirty_1_114; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2172 = _GEN_19863 | dirty_1_115; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2173 = _GEN_19864 | dirty_1_116; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2174 = _GEN_19865 | dirty_1_117; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2175 = _GEN_19866 | dirty_1_118; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2176 = _GEN_19867 | dirty_1_119; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2177 = _GEN_19868 | dirty_1_120; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2178 = _GEN_19869 | dirty_1_121; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2179 = _GEN_19870 | dirty_1_122; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2180 = _GEN_19871 | dirty_1_123; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2181 = _GEN_19872 | dirty_1_124; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2182 = _GEN_19873 | dirty_1_125; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2183 = _GEN_19874 | dirty_1_126; // @[d_cache.scala 131:{32,32} 33:26]
  wire  _GEN_2184 = _GEN_19875 | dirty_1_127; // @[d_cache.scala 131:{32,32} 33:26]
  wire [2:0] _GEN_2185 = way1_hit ? 3'h0 : 3'h4; // @[d_cache.scala 121:33 122:23 133:23]
  wire [63:0] _GEN_2186 = way1_hit ? _GEN_1161 : record_olddata_0; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2187 = way1_hit ? _GEN_1162 : record_olddata_1; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2188 = way1_hit ? _GEN_1163 : record_olddata_2; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2189 = way1_hit ? _GEN_1164 : record_olddata_3; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2190 = way1_hit ? _GEN_1165 : record_olddata_4; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2191 = way1_hit ? _GEN_1166 : record_olddata_5; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2192 = way1_hit ? _GEN_1167 : record_olddata_6; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2193 = way1_hit ? _GEN_1168 : record_olddata_7; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2194 = way1_hit ? _GEN_1169 : record_olddata_8; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2195 = way1_hit ? _GEN_1170 : record_olddata_9; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2196 = way1_hit ? _GEN_1171 : record_olddata_10; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2197 = way1_hit ? _GEN_1172 : record_olddata_11; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2198 = way1_hit ? _GEN_1173 : record_olddata_12; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2199 = way1_hit ? _GEN_1174 : record_olddata_13; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2200 = way1_hit ? _GEN_1175 : record_olddata_14; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2201 = way1_hit ? _GEN_1176 : record_olddata_15; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2202 = way1_hit ? _GEN_1177 : record_olddata_16; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2203 = way1_hit ? _GEN_1178 : record_olddata_17; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2204 = way1_hit ? _GEN_1179 : record_olddata_18; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2205 = way1_hit ? _GEN_1180 : record_olddata_19; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2206 = way1_hit ? _GEN_1181 : record_olddata_20; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2207 = way1_hit ? _GEN_1182 : record_olddata_21; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2208 = way1_hit ? _GEN_1183 : record_olddata_22; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2209 = way1_hit ? _GEN_1184 : record_olddata_23; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2210 = way1_hit ? _GEN_1185 : record_olddata_24; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2211 = way1_hit ? _GEN_1186 : record_olddata_25; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2212 = way1_hit ? _GEN_1187 : record_olddata_26; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2213 = way1_hit ? _GEN_1188 : record_olddata_27; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2214 = way1_hit ? _GEN_1189 : record_olddata_28; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2215 = way1_hit ? _GEN_1190 : record_olddata_29; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2216 = way1_hit ? _GEN_1191 : record_olddata_30; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2217 = way1_hit ? _GEN_1192 : record_olddata_31; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2218 = way1_hit ? _GEN_1193 : record_olddata_32; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2219 = way1_hit ? _GEN_1194 : record_olddata_33; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2220 = way1_hit ? _GEN_1195 : record_olddata_34; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2221 = way1_hit ? _GEN_1196 : record_olddata_35; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2222 = way1_hit ? _GEN_1197 : record_olddata_36; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2223 = way1_hit ? _GEN_1198 : record_olddata_37; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2224 = way1_hit ? _GEN_1199 : record_olddata_38; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2225 = way1_hit ? _GEN_1200 : record_olddata_39; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2226 = way1_hit ? _GEN_1201 : record_olddata_40; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2227 = way1_hit ? _GEN_1202 : record_olddata_41; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2228 = way1_hit ? _GEN_1203 : record_olddata_42; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2229 = way1_hit ? _GEN_1204 : record_olddata_43; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2230 = way1_hit ? _GEN_1205 : record_olddata_44; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2231 = way1_hit ? _GEN_1206 : record_olddata_45; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2232 = way1_hit ? _GEN_1207 : record_olddata_46; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2233 = way1_hit ? _GEN_1208 : record_olddata_47; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2234 = way1_hit ? _GEN_1209 : record_olddata_48; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2235 = way1_hit ? _GEN_1210 : record_olddata_49; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2236 = way1_hit ? _GEN_1211 : record_olddata_50; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2237 = way1_hit ? _GEN_1212 : record_olddata_51; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2238 = way1_hit ? _GEN_1213 : record_olddata_52; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2239 = way1_hit ? _GEN_1214 : record_olddata_53; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2240 = way1_hit ? _GEN_1215 : record_olddata_54; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2241 = way1_hit ? _GEN_1216 : record_olddata_55; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2242 = way1_hit ? _GEN_1217 : record_olddata_56; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2243 = way1_hit ? _GEN_1218 : record_olddata_57; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2244 = way1_hit ? _GEN_1219 : record_olddata_58; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2245 = way1_hit ? _GEN_1220 : record_olddata_59; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2246 = way1_hit ? _GEN_1221 : record_olddata_60; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2247 = way1_hit ? _GEN_1222 : record_olddata_61; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2248 = way1_hit ? _GEN_1223 : record_olddata_62; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2249 = way1_hit ? _GEN_1224 : record_olddata_63; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2250 = way1_hit ? _GEN_1225 : record_olddata_64; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2251 = way1_hit ? _GEN_1226 : record_olddata_65; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2252 = way1_hit ? _GEN_1227 : record_olddata_66; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2253 = way1_hit ? _GEN_1228 : record_olddata_67; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2254 = way1_hit ? _GEN_1229 : record_olddata_68; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2255 = way1_hit ? _GEN_1230 : record_olddata_69; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2256 = way1_hit ? _GEN_1231 : record_olddata_70; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2257 = way1_hit ? _GEN_1232 : record_olddata_71; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2258 = way1_hit ? _GEN_1233 : record_olddata_72; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2259 = way1_hit ? _GEN_1234 : record_olddata_73; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2260 = way1_hit ? _GEN_1235 : record_olddata_74; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2261 = way1_hit ? _GEN_1236 : record_olddata_75; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2262 = way1_hit ? _GEN_1237 : record_olddata_76; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2263 = way1_hit ? _GEN_1238 : record_olddata_77; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2264 = way1_hit ? _GEN_1239 : record_olddata_78; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2265 = way1_hit ? _GEN_1240 : record_olddata_79; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2266 = way1_hit ? _GEN_1241 : record_olddata_80; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2267 = way1_hit ? _GEN_1242 : record_olddata_81; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2268 = way1_hit ? _GEN_1243 : record_olddata_82; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2269 = way1_hit ? _GEN_1244 : record_olddata_83; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2270 = way1_hit ? _GEN_1245 : record_olddata_84; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2271 = way1_hit ? _GEN_1246 : record_olddata_85; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2272 = way1_hit ? _GEN_1247 : record_olddata_86; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2273 = way1_hit ? _GEN_1248 : record_olddata_87; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2274 = way1_hit ? _GEN_1249 : record_olddata_88; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2275 = way1_hit ? _GEN_1250 : record_olddata_89; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2276 = way1_hit ? _GEN_1251 : record_olddata_90; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2277 = way1_hit ? _GEN_1252 : record_olddata_91; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2278 = way1_hit ? _GEN_1253 : record_olddata_92; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2279 = way1_hit ? _GEN_1254 : record_olddata_93; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2280 = way1_hit ? _GEN_1255 : record_olddata_94; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2281 = way1_hit ? _GEN_1256 : record_olddata_95; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2282 = way1_hit ? _GEN_1257 : record_olddata_96; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2283 = way1_hit ? _GEN_1258 : record_olddata_97; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2284 = way1_hit ? _GEN_1259 : record_olddata_98; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2285 = way1_hit ? _GEN_1260 : record_olddata_99; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2286 = way1_hit ? _GEN_1261 : record_olddata_100; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2287 = way1_hit ? _GEN_1262 : record_olddata_101; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2288 = way1_hit ? _GEN_1263 : record_olddata_102; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2289 = way1_hit ? _GEN_1264 : record_olddata_103; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2290 = way1_hit ? _GEN_1265 : record_olddata_104; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2291 = way1_hit ? _GEN_1266 : record_olddata_105; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2292 = way1_hit ? _GEN_1267 : record_olddata_106; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2293 = way1_hit ? _GEN_1268 : record_olddata_107; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2294 = way1_hit ? _GEN_1269 : record_olddata_108; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2295 = way1_hit ? _GEN_1270 : record_olddata_109; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2296 = way1_hit ? _GEN_1271 : record_olddata_110; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2297 = way1_hit ? _GEN_1272 : record_olddata_111; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2298 = way1_hit ? _GEN_1273 : record_olddata_112; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2299 = way1_hit ? _GEN_1274 : record_olddata_113; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2300 = way1_hit ? _GEN_1275 : record_olddata_114; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2301 = way1_hit ? _GEN_1276 : record_olddata_115; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2302 = way1_hit ? _GEN_1277 : record_olddata_116; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2303 = way1_hit ? _GEN_1278 : record_olddata_117; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2304 = way1_hit ? _GEN_1279 : record_olddata_118; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2305 = way1_hit ? _GEN_1280 : record_olddata_119; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2306 = way1_hit ? _GEN_1281 : record_olddata_120; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2307 = way1_hit ? _GEN_1282 : record_olddata_121; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2308 = way1_hit ? _GEN_1283 : record_olddata_122; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2309 = way1_hit ? _GEN_1284 : record_olddata_123; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2310 = way1_hit ? _GEN_1285 : record_olddata_124; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2311 = way1_hit ? _GEN_1286 : record_olddata_125; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2312 = way1_hit ? _GEN_1287 : record_olddata_126; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2313 = way1_hit ? _GEN_1288 : record_olddata_127; // @[d_cache.scala 121:33 25:33]
  wire [63:0] _GEN_2314 = way1_hit ? _GEN_1417 : ram_1_0; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2315 = way1_hit ? _GEN_1418 : ram_1_1; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2316 = way1_hit ? _GEN_1419 : ram_1_2; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2317 = way1_hit ? _GEN_1420 : ram_1_3; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2318 = way1_hit ? _GEN_1421 : ram_1_4; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2319 = way1_hit ? _GEN_1422 : ram_1_5; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2320 = way1_hit ? _GEN_1423 : ram_1_6; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2321 = way1_hit ? _GEN_1424 : ram_1_7; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2322 = way1_hit ? _GEN_1425 : ram_1_8; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2323 = way1_hit ? _GEN_1426 : ram_1_9; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2324 = way1_hit ? _GEN_1427 : ram_1_10; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2325 = way1_hit ? _GEN_1428 : ram_1_11; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2326 = way1_hit ? _GEN_1429 : ram_1_12; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2327 = way1_hit ? _GEN_1430 : ram_1_13; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2328 = way1_hit ? _GEN_1431 : ram_1_14; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2329 = way1_hit ? _GEN_1432 : ram_1_15; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2330 = way1_hit ? _GEN_1433 : ram_1_16; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2331 = way1_hit ? _GEN_1434 : ram_1_17; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2332 = way1_hit ? _GEN_1435 : ram_1_18; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2333 = way1_hit ? _GEN_1436 : ram_1_19; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2334 = way1_hit ? _GEN_1437 : ram_1_20; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2335 = way1_hit ? _GEN_1438 : ram_1_21; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2336 = way1_hit ? _GEN_1439 : ram_1_22; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2337 = way1_hit ? _GEN_1440 : ram_1_23; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2338 = way1_hit ? _GEN_1441 : ram_1_24; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2339 = way1_hit ? _GEN_1442 : ram_1_25; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2340 = way1_hit ? _GEN_1443 : ram_1_26; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2341 = way1_hit ? _GEN_1444 : ram_1_27; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2342 = way1_hit ? _GEN_1445 : ram_1_28; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2343 = way1_hit ? _GEN_1446 : ram_1_29; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2344 = way1_hit ? _GEN_1447 : ram_1_30; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2345 = way1_hit ? _GEN_1448 : ram_1_31; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2346 = way1_hit ? _GEN_1449 : ram_1_32; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2347 = way1_hit ? _GEN_1450 : ram_1_33; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2348 = way1_hit ? _GEN_1451 : ram_1_34; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2349 = way1_hit ? _GEN_1452 : ram_1_35; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2350 = way1_hit ? _GEN_1453 : ram_1_36; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2351 = way1_hit ? _GEN_1454 : ram_1_37; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2352 = way1_hit ? _GEN_1455 : ram_1_38; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2353 = way1_hit ? _GEN_1456 : ram_1_39; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2354 = way1_hit ? _GEN_1457 : ram_1_40; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2355 = way1_hit ? _GEN_1458 : ram_1_41; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2356 = way1_hit ? _GEN_1459 : ram_1_42; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2357 = way1_hit ? _GEN_1460 : ram_1_43; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2358 = way1_hit ? _GEN_1461 : ram_1_44; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2359 = way1_hit ? _GEN_1462 : ram_1_45; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2360 = way1_hit ? _GEN_1463 : ram_1_46; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2361 = way1_hit ? _GEN_1464 : ram_1_47; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2362 = way1_hit ? _GEN_1465 : ram_1_48; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2363 = way1_hit ? _GEN_1466 : ram_1_49; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2364 = way1_hit ? _GEN_1467 : ram_1_50; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2365 = way1_hit ? _GEN_1468 : ram_1_51; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2366 = way1_hit ? _GEN_1469 : ram_1_52; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2367 = way1_hit ? _GEN_1470 : ram_1_53; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2368 = way1_hit ? _GEN_1471 : ram_1_54; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2369 = way1_hit ? _GEN_1472 : ram_1_55; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2370 = way1_hit ? _GEN_1473 : ram_1_56; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2371 = way1_hit ? _GEN_1474 : ram_1_57; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2372 = way1_hit ? _GEN_1475 : ram_1_58; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2373 = way1_hit ? _GEN_1476 : ram_1_59; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2374 = way1_hit ? _GEN_1477 : ram_1_60; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2375 = way1_hit ? _GEN_1478 : ram_1_61; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2376 = way1_hit ? _GEN_1479 : ram_1_62; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2377 = way1_hit ? _GEN_1480 : ram_1_63; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2378 = way1_hit ? _GEN_1481 : ram_1_64; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2379 = way1_hit ? _GEN_1482 : ram_1_65; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2380 = way1_hit ? _GEN_1483 : ram_1_66; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2381 = way1_hit ? _GEN_1484 : ram_1_67; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2382 = way1_hit ? _GEN_1485 : ram_1_68; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2383 = way1_hit ? _GEN_1486 : ram_1_69; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2384 = way1_hit ? _GEN_1487 : ram_1_70; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2385 = way1_hit ? _GEN_1488 : ram_1_71; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2386 = way1_hit ? _GEN_1489 : ram_1_72; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2387 = way1_hit ? _GEN_1490 : ram_1_73; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2388 = way1_hit ? _GEN_1491 : ram_1_74; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2389 = way1_hit ? _GEN_1492 : ram_1_75; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2390 = way1_hit ? _GEN_1493 : ram_1_76; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2391 = way1_hit ? _GEN_1494 : ram_1_77; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2392 = way1_hit ? _GEN_1495 : ram_1_78; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2393 = way1_hit ? _GEN_1496 : ram_1_79; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2394 = way1_hit ? _GEN_1497 : ram_1_80; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2395 = way1_hit ? _GEN_1498 : ram_1_81; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2396 = way1_hit ? _GEN_1499 : ram_1_82; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2397 = way1_hit ? _GEN_1500 : ram_1_83; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2398 = way1_hit ? _GEN_1501 : ram_1_84; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2399 = way1_hit ? _GEN_1502 : ram_1_85; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2400 = way1_hit ? _GEN_1503 : ram_1_86; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2401 = way1_hit ? _GEN_1504 : ram_1_87; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2402 = way1_hit ? _GEN_1505 : ram_1_88; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2403 = way1_hit ? _GEN_1506 : ram_1_89; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2404 = way1_hit ? _GEN_1507 : ram_1_90; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2405 = way1_hit ? _GEN_1508 : ram_1_91; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2406 = way1_hit ? _GEN_1509 : ram_1_92; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2407 = way1_hit ? _GEN_1510 : ram_1_93; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2408 = way1_hit ? _GEN_1511 : ram_1_94; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2409 = way1_hit ? _GEN_1512 : ram_1_95; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2410 = way1_hit ? _GEN_1513 : ram_1_96; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2411 = way1_hit ? _GEN_1514 : ram_1_97; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2412 = way1_hit ? _GEN_1515 : ram_1_98; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2413 = way1_hit ? _GEN_1516 : ram_1_99; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2414 = way1_hit ? _GEN_1517 : ram_1_100; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2415 = way1_hit ? _GEN_1518 : ram_1_101; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2416 = way1_hit ? _GEN_1519 : ram_1_102; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2417 = way1_hit ? _GEN_1520 : ram_1_103; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2418 = way1_hit ? _GEN_1521 : ram_1_104; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2419 = way1_hit ? _GEN_1522 : ram_1_105; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2420 = way1_hit ? _GEN_1523 : ram_1_106; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2421 = way1_hit ? _GEN_1524 : ram_1_107; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2422 = way1_hit ? _GEN_1525 : ram_1_108; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2423 = way1_hit ? _GEN_1526 : ram_1_109; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2424 = way1_hit ? _GEN_1527 : ram_1_110; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2425 = way1_hit ? _GEN_1528 : ram_1_111; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2426 = way1_hit ? _GEN_1529 : ram_1_112; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2427 = way1_hit ? _GEN_1530 : ram_1_113; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2428 = way1_hit ? _GEN_1531 : ram_1_114; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2429 = way1_hit ? _GEN_1532 : ram_1_115; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2430 = way1_hit ? _GEN_1533 : ram_1_116; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2431 = way1_hit ? _GEN_1534 : ram_1_117; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2432 = way1_hit ? _GEN_1535 : ram_1_118; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2433 = way1_hit ? _GEN_1536 : ram_1_119; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2434 = way1_hit ? _GEN_1537 : ram_1_120; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2435 = way1_hit ? _GEN_1538 : ram_1_121; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2436 = way1_hit ? _GEN_1539 : ram_1_122; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2437 = way1_hit ? _GEN_1540 : ram_1_123; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2438 = way1_hit ? _GEN_1541 : ram_1_124; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2439 = way1_hit ? _GEN_1542 : ram_1_125; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2440 = way1_hit ? _GEN_1543 : ram_1_126; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2441 = way1_hit ? _GEN_1544 : ram_1_127; // @[d_cache.scala 121:33 20:24]
  wire [63:0] _GEN_2442 = way1_hit ? _GEN_1545 : record_wdata1_0; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2443 = way1_hit ? _GEN_1546 : record_wdata1_1; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2444 = way1_hit ? _GEN_1547 : record_wdata1_2; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2445 = way1_hit ? _GEN_1548 : record_wdata1_3; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2446 = way1_hit ? _GEN_1549 : record_wdata1_4; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2447 = way1_hit ? _GEN_1550 : record_wdata1_5; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2448 = way1_hit ? _GEN_1551 : record_wdata1_6; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2449 = way1_hit ? _GEN_1552 : record_wdata1_7; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2450 = way1_hit ? _GEN_1553 : record_wdata1_8; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2451 = way1_hit ? _GEN_1554 : record_wdata1_9; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2452 = way1_hit ? _GEN_1555 : record_wdata1_10; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2453 = way1_hit ? _GEN_1556 : record_wdata1_11; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2454 = way1_hit ? _GEN_1557 : record_wdata1_12; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2455 = way1_hit ? _GEN_1558 : record_wdata1_13; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2456 = way1_hit ? _GEN_1559 : record_wdata1_14; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2457 = way1_hit ? _GEN_1560 : record_wdata1_15; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2458 = way1_hit ? _GEN_1561 : record_wdata1_16; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2459 = way1_hit ? _GEN_1562 : record_wdata1_17; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2460 = way1_hit ? _GEN_1563 : record_wdata1_18; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2461 = way1_hit ? _GEN_1564 : record_wdata1_19; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2462 = way1_hit ? _GEN_1565 : record_wdata1_20; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2463 = way1_hit ? _GEN_1566 : record_wdata1_21; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2464 = way1_hit ? _GEN_1567 : record_wdata1_22; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2465 = way1_hit ? _GEN_1568 : record_wdata1_23; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2466 = way1_hit ? _GEN_1569 : record_wdata1_24; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2467 = way1_hit ? _GEN_1570 : record_wdata1_25; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2468 = way1_hit ? _GEN_1571 : record_wdata1_26; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2469 = way1_hit ? _GEN_1572 : record_wdata1_27; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2470 = way1_hit ? _GEN_1573 : record_wdata1_28; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2471 = way1_hit ? _GEN_1574 : record_wdata1_29; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2472 = way1_hit ? _GEN_1575 : record_wdata1_30; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2473 = way1_hit ? _GEN_1576 : record_wdata1_31; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2474 = way1_hit ? _GEN_1577 : record_wdata1_32; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2475 = way1_hit ? _GEN_1578 : record_wdata1_33; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2476 = way1_hit ? _GEN_1579 : record_wdata1_34; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2477 = way1_hit ? _GEN_1580 : record_wdata1_35; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2478 = way1_hit ? _GEN_1581 : record_wdata1_36; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2479 = way1_hit ? _GEN_1582 : record_wdata1_37; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2480 = way1_hit ? _GEN_1583 : record_wdata1_38; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2481 = way1_hit ? _GEN_1584 : record_wdata1_39; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2482 = way1_hit ? _GEN_1585 : record_wdata1_40; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2483 = way1_hit ? _GEN_1586 : record_wdata1_41; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2484 = way1_hit ? _GEN_1587 : record_wdata1_42; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2485 = way1_hit ? _GEN_1588 : record_wdata1_43; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2486 = way1_hit ? _GEN_1589 : record_wdata1_44; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2487 = way1_hit ? _GEN_1590 : record_wdata1_45; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2488 = way1_hit ? _GEN_1591 : record_wdata1_46; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2489 = way1_hit ? _GEN_1592 : record_wdata1_47; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2490 = way1_hit ? _GEN_1593 : record_wdata1_48; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2491 = way1_hit ? _GEN_1594 : record_wdata1_49; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2492 = way1_hit ? _GEN_1595 : record_wdata1_50; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2493 = way1_hit ? _GEN_1596 : record_wdata1_51; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2494 = way1_hit ? _GEN_1597 : record_wdata1_52; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2495 = way1_hit ? _GEN_1598 : record_wdata1_53; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2496 = way1_hit ? _GEN_1599 : record_wdata1_54; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2497 = way1_hit ? _GEN_1600 : record_wdata1_55; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2498 = way1_hit ? _GEN_1601 : record_wdata1_56; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2499 = way1_hit ? _GEN_1602 : record_wdata1_57; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2500 = way1_hit ? _GEN_1603 : record_wdata1_58; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2501 = way1_hit ? _GEN_1604 : record_wdata1_59; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2502 = way1_hit ? _GEN_1605 : record_wdata1_60; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2503 = way1_hit ? _GEN_1606 : record_wdata1_61; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2504 = way1_hit ? _GEN_1607 : record_wdata1_62; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2505 = way1_hit ? _GEN_1608 : record_wdata1_63; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2506 = way1_hit ? _GEN_1609 : record_wdata1_64; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2507 = way1_hit ? _GEN_1610 : record_wdata1_65; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2508 = way1_hit ? _GEN_1611 : record_wdata1_66; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2509 = way1_hit ? _GEN_1612 : record_wdata1_67; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2510 = way1_hit ? _GEN_1613 : record_wdata1_68; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2511 = way1_hit ? _GEN_1614 : record_wdata1_69; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2512 = way1_hit ? _GEN_1615 : record_wdata1_70; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2513 = way1_hit ? _GEN_1616 : record_wdata1_71; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2514 = way1_hit ? _GEN_1617 : record_wdata1_72; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2515 = way1_hit ? _GEN_1618 : record_wdata1_73; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2516 = way1_hit ? _GEN_1619 : record_wdata1_74; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2517 = way1_hit ? _GEN_1620 : record_wdata1_75; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2518 = way1_hit ? _GEN_1621 : record_wdata1_76; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2519 = way1_hit ? _GEN_1622 : record_wdata1_77; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2520 = way1_hit ? _GEN_1623 : record_wdata1_78; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2521 = way1_hit ? _GEN_1624 : record_wdata1_79; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2522 = way1_hit ? _GEN_1625 : record_wdata1_80; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2523 = way1_hit ? _GEN_1626 : record_wdata1_81; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2524 = way1_hit ? _GEN_1627 : record_wdata1_82; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2525 = way1_hit ? _GEN_1628 : record_wdata1_83; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2526 = way1_hit ? _GEN_1629 : record_wdata1_84; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2527 = way1_hit ? _GEN_1630 : record_wdata1_85; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2528 = way1_hit ? _GEN_1631 : record_wdata1_86; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2529 = way1_hit ? _GEN_1632 : record_wdata1_87; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2530 = way1_hit ? _GEN_1633 : record_wdata1_88; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2531 = way1_hit ? _GEN_1634 : record_wdata1_89; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2532 = way1_hit ? _GEN_1635 : record_wdata1_90; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2533 = way1_hit ? _GEN_1636 : record_wdata1_91; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2534 = way1_hit ? _GEN_1637 : record_wdata1_92; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2535 = way1_hit ? _GEN_1638 : record_wdata1_93; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2536 = way1_hit ? _GEN_1639 : record_wdata1_94; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2537 = way1_hit ? _GEN_1640 : record_wdata1_95; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2538 = way1_hit ? _GEN_1641 : record_wdata1_96; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2539 = way1_hit ? _GEN_1642 : record_wdata1_97; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2540 = way1_hit ? _GEN_1643 : record_wdata1_98; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2541 = way1_hit ? _GEN_1644 : record_wdata1_99; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2542 = way1_hit ? _GEN_1645 : record_wdata1_100; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2543 = way1_hit ? _GEN_1646 : record_wdata1_101; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2544 = way1_hit ? _GEN_1647 : record_wdata1_102; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2545 = way1_hit ? _GEN_1648 : record_wdata1_103; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2546 = way1_hit ? _GEN_1649 : record_wdata1_104; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2547 = way1_hit ? _GEN_1650 : record_wdata1_105; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2548 = way1_hit ? _GEN_1651 : record_wdata1_106; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2549 = way1_hit ? _GEN_1652 : record_wdata1_107; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2550 = way1_hit ? _GEN_1653 : record_wdata1_108; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2551 = way1_hit ? _GEN_1654 : record_wdata1_109; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2552 = way1_hit ? _GEN_1655 : record_wdata1_110; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2553 = way1_hit ? _GEN_1656 : record_wdata1_111; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2554 = way1_hit ? _GEN_1657 : record_wdata1_112; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2555 = way1_hit ? _GEN_1658 : record_wdata1_113; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2556 = way1_hit ? _GEN_1659 : record_wdata1_114; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2557 = way1_hit ? _GEN_1660 : record_wdata1_115; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2558 = way1_hit ? _GEN_1661 : record_wdata1_116; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2559 = way1_hit ? _GEN_1662 : record_wdata1_117; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2560 = way1_hit ? _GEN_1663 : record_wdata1_118; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2561 = way1_hit ? _GEN_1664 : record_wdata1_119; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2562 = way1_hit ? _GEN_1665 : record_wdata1_120; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2563 = way1_hit ? _GEN_1666 : record_wdata1_121; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2564 = way1_hit ? _GEN_1667 : record_wdata1_122; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2565 = way1_hit ? _GEN_1668 : record_wdata1_123; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2566 = way1_hit ? _GEN_1669 : record_wdata1_124; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2567 = way1_hit ? _GEN_1670 : record_wdata1_125; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2568 = way1_hit ? _GEN_1671 : record_wdata1_126; // @[d_cache.scala 121:33 21:32]
  wire [63:0] _GEN_2569 = way1_hit ? _GEN_1672 : record_wdata1_127; // @[d_cache.scala 121:33 21:32]
  wire [7:0] _GEN_2570 = way1_hit ? _GEN_1673 : record_wstrb1_0; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2571 = way1_hit ? _GEN_1674 : record_wstrb1_1; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2572 = way1_hit ? _GEN_1675 : record_wstrb1_2; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2573 = way1_hit ? _GEN_1676 : record_wstrb1_3; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2574 = way1_hit ? _GEN_1677 : record_wstrb1_4; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2575 = way1_hit ? _GEN_1678 : record_wstrb1_5; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2576 = way1_hit ? _GEN_1679 : record_wstrb1_6; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2577 = way1_hit ? _GEN_1680 : record_wstrb1_7; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2578 = way1_hit ? _GEN_1681 : record_wstrb1_8; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2579 = way1_hit ? _GEN_1682 : record_wstrb1_9; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2580 = way1_hit ? _GEN_1683 : record_wstrb1_10; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2581 = way1_hit ? _GEN_1684 : record_wstrb1_11; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2582 = way1_hit ? _GEN_1685 : record_wstrb1_12; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2583 = way1_hit ? _GEN_1686 : record_wstrb1_13; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2584 = way1_hit ? _GEN_1687 : record_wstrb1_14; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2585 = way1_hit ? _GEN_1688 : record_wstrb1_15; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2586 = way1_hit ? _GEN_1689 : record_wstrb1_16; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2587 = way1_hit ? _GEN_1690 : record_wstrb1_17; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2588 = way1_hit ? _GEN_1691 : record_wstrb1_18; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2589 = way1_hit ? _GEN_1692 : record_wstrb1_19; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2590 = way1_hit ? _GEN_1693 : record_wstrb1_20; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2591 = way1_hit ? _GEN_1694 : record_wstrb1_21; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2592 = way1_hit ? _GEN_1695 : record_wstrb1_22; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2593 = way1_hit ? _GEN_1696 : record_wstrb1_23; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2594 = way1_hit ? _GEN_1697 : record_wstrb1_24; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2595 = way1_hit ? _GEN_1698 : record_wstrb1_25; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2596 = way1_hit ? _GEN_1699 : record_wstrb1_26; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2597 = way1_hit ? _GEN_1700 : record_wstrb1_27; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2598 = way1_hit ? _GEN_1701 : record_wstrb1_28; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2599 = way1_hit ? _GEN_1702 : record_wstrb1_29; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2600 = way1_hit ? _GEN_1703 : record_wstrb1_30; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2601 = way1_hit ? _GEN_1704 : record_wstrb1_31; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2602 = way1_hit ? _GEN_1705 : record_wstrb1_32; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2603 = way1_hit ? _GEN_1706 : record_wstrb1_33; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2604 = way1_hit ? _GEN_1707 : record_wstrb1_34; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2605 = way1_hit ? _GEN_1708 : record_wstrb1_35; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2606 = way1_hit ? _GEN_1709 : record_wstrb1_36; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2607 = way1_hit ? _GEN_1710 : record_wstrb1_37; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2608 = way1_hit ? _GEN_1711 : record_wstrb1_38; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2609 = way1_hit ? _GEN_1712 : record_wstrb1_39; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2610 = way1_hit ? _GEN_1713 : record_wstrb1_40; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2611 = way1_hit ? _GEN_1714 : record_wstrb1_41; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2612 = way1_hit ? _GEN_1715 : record_wstrb1_42; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2613 = way1_hit ? _GEN_1716 : record_wstrb1_43; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2614 = way1_hit ? _GEN_1717 : record_wstrb1_44; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2615 = way1_hit ? _GEN_1718 : record_wstrb1_45; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2616 = way1_hit ? _GEN_1719 : record_wstrb1_46; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2617 = way1_hit ? _GEN_1720 : record_wstrb1_47; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2618 = way1_hit ? _GEN_1721 : record_wstrb1_48; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2619 = way1_hit ? _GEN_1722 : record_wstrb1_49; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2620 = way1_hit ? _GEN_1723 : record_wstrb1_50; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2621 = way1_hit ? _GEN_1724 : record_wstrb1_51; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2622 = way1_hit ? _GEN_1725 : record_wstrb1_52; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2623 = way1_hit ? _GEN_1726 : record_wstrb1_53; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2624 = way1_hit ? _GEN_1727 : record_wstrb1_54; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2625 = way1_hit ? _GEN_1728 : record_wstrb1_55; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2626 = way1_hit ? _GEN_1729 : record_wstrb1_56; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2627 = way1_hit ? _GEN_1730 : record_wstrb1_57; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2628 = way1_hit ? _GEN_1731 : record_wstrb1_58; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2629 = way1_hit ? _GEN_1732 : record_wstrb1_59; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2630 = way1_hit ? _GEN_1733 : record_wstrb1_60; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2631 = way1_hit ? _GEN_1734 : record_wstrb1_61; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2632 = way1_hit ? _GEN_1735 : record_wstrb1_62; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2633 = way1_hit ? _GEN_1736 : record_wstrb1_63; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2634 = way1_hit ? _GEN_1737 : record_wstrb1_64; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2635 = way1_hit ? _GEN_1738 : record_wstrb1_65; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2636 = way1_hit ? _GEN_1739 : record_wstrb1_66; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2637 = way1_hit ? _GEN_1740 : record_wstrb1_67; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2638 = way1_hit ? _GEN_1741 : record_wstrb1_68; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2639 = way1_hit ? _GEN_1742 : record_wstrb1_69; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2640 = way1_hit ? _GEN_1743 : record_wstrb1_70; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2641 = way1_hit ? _GEN_1744 : record_wstrb1_71; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2642 = way1_hit ? _GEN_1745 : record_wstrb1_72; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2643 = way1_hit ? _GEN_1746 : record_wstrb1_73; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2644 = way1_hit ? _GEN_1747 : record_wstrb1_74; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2645 = way1_hit ? _GEN_1748 : record_wstrb1_75; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2646 = way1_hit ? _GEN_1749 : record_wstrb1_76; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2647 = way1_hit ? _GEN_1750 : record_wstrb1_77; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2648 = way1_hit ? _GEN_1751 : record_wstrb1_78; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2649 = way1_hit ? _GEN_1752 : record_wstrb1_79; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2650 = way1_hit ? _GEN_1753 : record_wstrb1_80; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2651 = way1_hit ? _GEN_1754 : record_wstrb1_81; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2652 = way1_hit ? _GEN_1755 : record_wstrb1_82; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2653 = way1_hit ? _GEN_1756 : record_wstrb1_83; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2654 = way1_hit ? _GEN_1757 : record_wstrb1_84; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2655 = way1_hit ? _GEN_1758 : record_wstrb1_85; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2656 = way1_hit ? _GEN_1759 : record_wstrb1_86; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2657 = way1_hit ? _GEN_1760 : record_wstrb1_87; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2658 = way1_hit ? _GEN_1761 : record_wstrb1_88; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2659 = way1_hit ? _GEN_1762 : record_wstrb1_89; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2660 = way1_hit ? _GEN_1763 : record_wstrb1_90; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2661 = way1_hit ? _GEN_1764 : record_wstrb1_91; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2662 = way1_hit ? _GEN_1765 : record_wstrb1_92; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2663 = way1_hit ? _GEN_1766 : record_wstrb1_93; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2664 = way1_hit ? _GEN_1767 : record_wstrb1_94; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2665 = way1_hit ? _GEN_1768 : record_wstrb1_95; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2666 = way1_hit ? _GEN_1769 : record_wstrb1_96; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2667 = way1_hit ? _GEN_1770 : record_wstrb1_97; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2668 = way1_hit ? _GEN_1771 : record_wstrb1_98; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2669 = way1_hit ? _GEN_1772 : record_wstrb1_99; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2670 = way1_hit ? _GEN_1773 : record_wstrb1_100; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2671 = way1_hit ? _GEN_1774 : record_wstrb1_101; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2672 = way1_hit ? _GEN_1775 : record_wstrb1_102; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2673 = way1_hit ? _GEN_1776 : record_wstrb1_103; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2674 = way1_hit ? _GEN_1777 : record_wstrb1_104; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2675 = way1_hit ? _GEN_1778 : record_wstrb1_105; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2676 = way1_hit ? _GEN_1779 : record_wstrb1_106; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2677 = way1_hit ? _GEN_1780 : record_wstrb1_107; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2678 = way1_hit ? _GEN_1781 : record_wstrb1_108; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2679 = way1_hit ? _GEN_1782 : record_wstrb1_109; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2680 = way1_hit ? _GEN_1783 : record_wstrb1_110; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2681 = way1_hit ? _GEN_1784 : record_wstrb1_111; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2682 = way1_hit ? _GEN_1785 : record_wstrb1_112; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2683 = way1_hit ? _GEN_1786 : record_wstrb1_113; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2684 = way1_hit ? _GEN_1787 : record_wstrb1_114; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2685 = way1_hit ? _GEN_1788 : record_wstrb1_115; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2686 = way1_hit ? _GEN_1789 : record_wstrb1_116; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2687 = way1_hit ? _GEN_1790 : record_wstrb1_117; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2688 = way1_hit ? _GEN_1791 : record_wstrb1_118; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2689 = way1_hit ? _GEN_1792 : record_wstrb1_119; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2690 = way1_hit ? _GEN_1793 : record_wstrb1_120; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2691 = way1_hit ? _GEN_1794 : record_wstrb1_121; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2692 = way1_hit ? _GEN_1795 : record_wstrb1_122; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2693 = way1_hit ? _GEN_1796 : record_wstrb1_123; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2694 = way1_hit ? _GEN_1797 : record_wstrb1_124; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2695 = way1_hit ? _GEN_1798 : record_wstrb1_125; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2696 = way1_hit ? _GEN_1799 : record_wstrb1_126; // @[d_cache.scala 121:33 22:32]
  wire [7:0] _GEN_2697 = way1_hit ? _GEN_1800 : record_wstrb1_127; // @[d_cache.scala 121:33 22:32]
  wire [63:0] _GEN_2698 = way1_hit ? _GEN_1801 : record_pc_0; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2699 = way1_hit ? _GEN_1802 : record_pc_1; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2700 = way1_hit ? _GEN_1803 : record_pc_2; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2701 = way1_hit ? _GEN_1804 : record_pc_3; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2702 = way1_hit ? _GEN_1805 : record_pc_4; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2703 = way1_hit ? _GEN_1806 : record_pc_5; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2704 = way1_hit ? _GEN_1807 : record_pc_6; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2705 = way1_hit ? _GEN_1808 : record_pc_7; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2706 = way1_hit ? _GEN_1809 : record_pc_8; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2707 = way1_hit ? _GEN_1810 : record_pc_9; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2708 = way1_hit ? _GEN_1811 : record_pc_10; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2709 = way1_hit ? _GEN_1812 : record_pc_11; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2710 = way1_hit ? _GEN_1813 : record_pc_12; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2711 = way1_hit ? _GEN_1814 : record_pc_13; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2712 = way1_hit ? _GEN_1815 : record_pc_14; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2713 = way1_hit ? _GEN_1816 : record_pc_15; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2714 = way1_hit ? _GEN_1817 : record_pc_16; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2715 = way1_hit ? _GEN_1818 : record_pc_17; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2716 = way1_hit ? _GEN_1819 : record_pc_18; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2717 = way1_hit ? _GEN_1820 : record_pc_19; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2718 = way1_hit ? _GEN_1821 : record_pc_20; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2719 = way1_hit ? _GEN_1822 : record_pc_21; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2720 = way1_hit ? _GEN_1823 : record_pc_22; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2721 = way1_hit ? _GEN_1824 : record_pc_23; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2722 = way1_hit ? _GEN_1825 : record_pc_24; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2723 = way1_hit ? _GEN_1826 : record_pc_25; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2724 = way1_hit ? _GEN_1827 : record_pc_26; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2725 = way1_hit ? _GEN_1828 : record_pc_27; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2726 = way1_hit ? _GEN_1829 : record_pc_28; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2727 = way1_hit ? _GEN_1830 : record_pc_29; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2728 = way1_hit ? _GEN_1831 : record_pc_30; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2729 = way1_hit ? _GEN_1832 : record_pc_31; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2730 = way1_hit ? _GEN_1833 : record_pc_32; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2731 = way1_hit ? _GEN_1834 : record_pc_33; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2732 = way1_hit ? _GEN_1835 : record_pc_34; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2733 = way1_hit ? _GEN_1836 : record_pc_35; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2734 = way1_hit ? _GEN_1837 : record_pc_36; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2735 = way1_hit ? _GEN_1838 : record_pc_37; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2736 = way1_hit ? _GEN_1839 : record_pc_38; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2737 = way1_hit ? _GEN_1840 : record_pc_39; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2738 = way1_hit ? _GEN_1841 : record_pc_40; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2739 = way1_hit ? _GEN_1842 : record_pc_41; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2740 = way1_hit ? _GEN_1843 : record_pc_42; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2741 = way1_hit ? _GEN_1844 : record_pc_43; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2742 = way1_hit ? _GEN_1845 : record_pc_44; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2743 = way1_hit ? _GEN_1846 : record_pc_45; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2744 = way1_hit ? _GEN_1847 : record_pc_46; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2745 = way1_hit ? _GEN_1848 : record_pc_47; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2746 = way1_hit ? _GEN_1849 : record_pc_48; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2747 = way1_hit ? _GEN_1850 : record_pc_49; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2748 = way1_hit ? _GEN_1851 : record_pc_50; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2749 = way1_hit ? _GEN_1852 : record_pc_51; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2750 = way1_hit ? _GEN_1853 : record_pc_52; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2751 = way1_hit ? _GEN_1854 : record_pc_53; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2752 = way1_hit ? _GEN_1855 : record_pc_54; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2753 = way1_hit ? _GEN_1856 : record_pc_55; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2754 = way1_hit ? _GEN_1857 : record_pc_56; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2755 = way1_hit ? _GEN_1858 : record_pc_57; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2756 = way1_hit ? _GEN_1859 : record_pc_58; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2757 = way1_hit ? _GEN_1860 : record_pc_59; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2758 = way1_hit ? _GEN_1861 : record_pc_60; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2759 = way1_hit ? _GEN_1862 : record_pc_61; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2760 = way1_hit ? _GEN_1863 : record_pc_62; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2761 = way1_hit ? _GEN_1864 : record_pc_63; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2762 = way1_hit ? _GEN_1865 : record_pc_64; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2763 = way1_hit ? _GEN_1866 : record_pc_65; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2764 = way1_hit ? _GEN_1867 : record_pc_66; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2765 = way1_hit ? _GEN_1868 : record_pc_67; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2766 = way1_hit ? _GEN_1869 : record_pc_68; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2767 = way1_hit ? _GEN_1870 : record_pc_69; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2768 = way1_hit ? _GEN_1871 : record_pc_70; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2769 = way1_hit ? _GEN_1872 : record_pc_71; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2770 = way1_hit ? _GEN_1873 : record_pc_72; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2771 = way1_hit ? _GEN_1874 : record_pc_73; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2772 = way1_hit ? _GEN_1875 : record_pc_74; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2773 = way1_hit ? _GEN_1876 : record_pc_75; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2774 = way1_hit ? _GEN_1877 : record_pc_76; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2775 = way1_hit ? _GEN_1878 : record_pc_77; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2776 = way1_hit ? _GEN_1879 : record_pc_78; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2777 = way1_hit ? _GEN_1880 : record_pc_79; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2778 = way1_hit ? _GEN_1881 : record_pc_80; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2779 = way1_hit ? _GEN_1882 : record_pc_81; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2780 = way1_hit ? _GEN_1883 : record_pc_82; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2781 = way1_hit ? _GEN_1884 : record_pc_83; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2782 = way1_hit ? _GEN_1885 : record_pc_84; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2783 = way1_hit ? _GEN_1886 : record_pc_85; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2784 = way1_hit ? _GEN_1887 : record_pc_86; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2785 = way1_hit ? _GEN_1888 : record_pc_87; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2786 = way1_hit ? _GEN_1889 : record_pc_88; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2787 = way1_hit ? _GEN_1890 : record_pc_89; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2788 = way1_hit ? _GEN_1891 : record_pc_90; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2789 = way1_hit ? _GEN_1892 : record_pc_91; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2790 = way1_hit ? _GEN_1893 : record_pc_92; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2791 = way1_hit ? _GEN_1894 : record_pc_93; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2792 = way1_hit ? _GEN_1895 : record_pc_94; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2793 = way1_hit ? _GEN_1896 : record_pc_95; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2794 = way1_hit ? _GEN_1897 : record_pc_96; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2795 = way1_hit ? _GEN_1898 : record_pc_97; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2796 = way1_hit ? _GEN_1899 : record_pc_98; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2797 = way1_hit ? _GEN_1900 : record_pc_99; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2798 = way1_hit ? _GEN_1901 : record_pc_100; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2799 = way1_hit ? _GEN_1902 : record_pc_101; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2800 = way1_hit ? _GEN_1903 : record_pc_102; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2801 = way1_hit ? _GEN_1904 : record_pc_103; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2802 = way1_hit ? _GEN_1905 : record_pc_104; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2803 = way1_hit ? _GEN_1906 : record_pc_105; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2804 = way1_hit ? _GEN_1907 : record_pc_106; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2805 = way1_hit ? _GEN_1908 : record_pc_107; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2806 = way1_hit ? _GEN_1909 : record_pc_108; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2807 = way1_hit ? _GEN_1910 : record_pc_109; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2808 = way1_hit ? _GEN_1911 : record_pc_110; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2809 = way1_hit ? _GEN_1912 : record_pc_111; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2810 = way1_hit ? _GEN_1913 : record_pc_112; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2811 = way1_hit ? _GEN_1914 : record_pc_113; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2812 = way1_hit ? _GEN_1915 : record_pc_114; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2813 = way1_hit ? _GEN_1916 : record_pc_115; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2814 = way1_hit ? _GEN_1917 : record_pc_116; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2815 = way1_hit ? _GEN_1918 : record_pc_117; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2816 = way1_hit ? _GEN_1919 : record_pc_118; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2817 = way1_hit ? _GEN_1920 : record_pc_119; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2818 = way1_hit ? _GEN_1921 : record_pc_120; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2819 = way1_hit ? _GEN_1922 : record_pc_121; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2820 = way1_hit ? _GEN_1923 : record_pc_122; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2821 = way1_hit ? _GEN_1924 : record_pc_123; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2822 = way1_hit ? _GEN_1925 : record_pc_124; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2823 = way1_hit ? _GEN_1926 : record_pc_125; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2824 = way1_hit ? _GEN_1927 : record_pc_126; // @[d_cache.scala 121:33 23:28]
  wire [63:0] _GEN_2825 = way1_hit ? _GEN_1928 : record_pc_127; // @[d_cache.scala 121:33 23:28]
  wire [31:0] _GEN_2826 = way1_hit ? _GEN_1929 : record_addr_0; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2827 = way1_hit ? _GEN_1930 : record_addr_1; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2828 = way1_hit ? _GEN_1931 : record_addr_2; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2829 = way1_hit ? _GEN_1932 : record_addr_3; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2830 = way1_hit ? _GEN_1933 : record_addr_4; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2831 = way1_hit ? _GEN_1934 : record_addr_5; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2832 = way1_hit ? _GEN_1935 : record_addr_6; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2833 = way1_hit ? _GEN_1936 : record_addr_7; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2834 = way1_hit ? _GEN_1937 : record_addr_8; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2835 = way1_hit ? _GEN_1938 : record_addr_9; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2836 = way1_hit ? _GEN_1939 : record_addr_10; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2837 = way1_hit ? _GEN_1940 : record_addr_11; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2838 = way1_hit ? _GEN_1941 : record_addr_12; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2839 = way1_hit ? _GEN_1942 : record_addr_13; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2840 = way1_hit ? _GEN_1943 : record_addr_14; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2841 = way1_hit ? _GEN_1944 : record_addr_15; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2842 = way1_hit ? _GEN_1945 : record_addr_16; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2843 = way1_hit ? _GEN_1946 : record_addr_17; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2844 = way1_hit ? _GEN_1947 : record_addr_18; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2845 = way1_hit ? _GEN_1948 : record_addr_19; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2846 = way1_hit ? _GEN_1949 : record_addr_20; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2847 = way1_hit ? _GEN_1950 : record_addr_21; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2848 = way1_hit ? _GEN_1951 : record_addr_22; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2849 = way1_hit ? _GEN_1952 : record_addr_23; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2850 = way1_hit ? _GEN_1953 : record_addr_24; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2851 = way1_hit ? _GEN_1954 : record_addr_25; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2852 = way1_hit ? _GEN_1955 : record_addr_26; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2853 = way1_hit ? _GEN_1956 : record_addr_27; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2854 = way1_hit ? _GEN_1957 : record_addr_28; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2855 = way1_hit ? _GEN_1958 : record_addr_29; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2856 = way1_hit ? _GEN_1959 : record_addr_30; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2857 = way1_hit ? _GEN_1960 : record_addr_31; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2858 = way1_hit ? _GEN_1961 : record_addr_32; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2859 = way1_hit ? _GEN_1962 : record_addr_33; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2860 = way1_hit ? _GEN_1963 : record_addr_34; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2861 = way1_hit ? _GEN_1964 : record_addr_35; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2862 = way1_hit ? _GEN_1965 : record_addr_36; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2863 = way1_hit ? _GEN_1966 : record_addr_37; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2864 = way1_hit ? _GEN_1967 : record_addr_38; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2865 = way1_hit ? _GEN_1968 : record_addr_39; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2866 = way1_hit ? _GEN_1969 : record_addr_40; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2867 = way1_hit ? _GEN_1970 : record_addr_41; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2868 = way1_hit ? _GEN_1971 : record_addr_42; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2869 = way1_hit ? _GEN_1972 : record_addr_43; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2870 = way1_hit ? _GEN_1973 : record_addr_44; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2871 = way1_hit ? _GEN_1974 : record_addr_45; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2872 = way1_hit ? _GEN_1975 : record_addr_46; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2873 = way1_hit ? _GEN_1976 : record_addr_47; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2874 = way1_hit ? _GEN_1977 : record_addr_48; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2875 = way1_hit ? _GEN_1978 : record_addr_49; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2876 = way1_hit ? _GEN_1979 : record_addr_50; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2877 = way1_hit ? _GEN_1980 : record_addr_51; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2878 = way1_hit ? _GEN_1981 : record_addr_52; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2879 = way1_hit ? _GEN_1982 : record_addr_53; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2880 = way1_hit ? _GEN_1983 : record_addr_54; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2881 = way1_hit ? _GEN_1984 : record_addr_55; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2882 = way1_hit ? _GEN_1985 : record_addr_56; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2883 = way1_hit ? _GEN_1986 : record_addr_57; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2884 = way1_hit ? _GEN_1987 : record_addr_58; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2885 = way1_hit ? _GEN_1988 : record_addr_59; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2886 = way1_hit ? _GEN_1989 : record_addr_60; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2887 = way1_hit ? _GEN_1990 : record_addr_61; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2888 = way1_hit ? _GEN_1991 : record_addr_62; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2889 = way1_hit ? _GEN_1992 : record_addr_63; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2890 = way1_hit ? _GEN_1993 : record_addr_64; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2891 = way1_hit ? _GEN_1994 : record_addr_65; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2892 = way1_hit ? _GEN_1995 : record_addr_66; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2893 = way1_hit ? _GEN_1996 : record_addr_67; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2894 = way1_hit ? _GEN_1997 : record_addr_68; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2895 = way1_hit ? _GEN_1998 : record_addr_69; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2896 = way1_hit ? _GEN_1999 : record_addr_70; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2897 = way1_hit ? _GEN_2000 : record_addr_71; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2898 = way1_hit ? _GEN_2001 : record_addr_72; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2899 = way1_hit ? _GEN_2002 : record_addr_73; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2900 = way1_hit ? _GEN_2003 : record_addr_74; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2901 = way1_hit ? _GEN_2004 : record_addr_75; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2902 = way1_hit ? _GEN_2005 : record_addr_76; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2903 = way1_hit ? _GEN_2006 : record_addr_77; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2904 = way1_hit ? _GEN_2007 : record_addr_78; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2905 = way1_hit ? _GEN_2008 : record_addr_79; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2906 = way1_hit ? _GEN_2009 : record_addr_80; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2907 = way1_hit ? _GEN_2010 : record_addr_81; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2908 = way1_hit ? _GEN_2011 : record_addr_82; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2909 = way1_hit ? _GEN_2012 : record_addr_83; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2910 = way1_hit ? _GEN_2013 : record_addr_84; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2911 = way1_hit ? _GEN_2014 : record_addr_85; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2912 = way1_hit ? _GEN_2015 : record_addr_86; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2913 = way1_hit ? _GEN_2016 : record_addr_87; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2914 = way1_hit ? _GEN_2017 : record_addr_88; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2915 = way1_hit ? _GEN_2018 : record_addr_89; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2916 = way1_hit ? _GEN_2019 : record_addr_90; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2917 = way1_hit ? _GEN_2020 : record_addr_91; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2918 = way1_hit ? _GEN_2021 : record_addr_92; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2919 = way1_hit ? _GEN_2022 : record_addr_93; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2920 = way1_hit ? _GEN_2023 : record_addr_94; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2921 = way1_hit ? _GEN_2024 : record_addr_95; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2922 = way1_hit ? _GEN_2025 : record_addr_96; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2923 = way1_hit ? _GEN_2026 : record_addr_97; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2924 = way1_hit ? _GEN_2027 : record_addr_98; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2925 = way1_hit ? _GEN_2028 : record_addr_99; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2926 = way1_hit ? _GEN_2029 : record_addr_100; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2927 = way1_hit ? _GEN_2030 : record_addr_101; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2928 = way1_hit ? _GEN_2031 : record_addr_102; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2929 = way1_hit ? _GEN_2032 : record_addr_103; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2930 = way1_hit ? _GEN_2033 : record_addr_104; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2931 = way1_hit ? _GEN_2034 : record_addr_105; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2932 = way1_hit ? _GEN_2035 : record_addr_106; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2933 = way1_hit ? _GEN_2036 : record_addr_107; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2934 = way1_hit ? _GEN_2037 : record_addr_108; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2935 = way1_hit ? _GEN_2038 : record_addr_109; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2936 = way1_hit ? _GEN_2039 : record_addr_110; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2937 = way1_hit ? _GEN_2040 : record_addr_111; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2938 = way1_hit ? _GEN_2041 : record_addr_112; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2939 = way1_hit ? _GEN_2042 : record_addr_113; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2940 = way1_hit ? _GEN_2043 : record_addr_114; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2941 = way1_hit ? _GEN_2044 : record_addr_115; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2942 = way1_hit ? _GEN_2045 : record_addr_116; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2943 = way1_hit ? _GEN_2046 : record_addr_117; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2944 = way1_hit ? _GEN_2047 : record_addr_118; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2945 = way1_hit ? _GEN_2048 : record_addr_119; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2946 = way1_hit ? _GEN_2049 : record_addr_120; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2947 = way1_hit ? _GEN_2050 : record_addr_121; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2948 = way1_hit ? _GEN_2051 : record_addr_122; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2949 = way1_hit ? _GEN_2052 : record_addr_123; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2950 = way1_hit ? _GEN_2053 : record_addr_124; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2951 = way1_hit ? _GEN_2054 : record_addr_125; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2952 = way1_hit ? _GEN_2055 : record_addr_126; // @[d_cache.scala 121:33 24:30]
  wire [31:0] _GEN_2953 = way1_hit ? _GEN_2056 : record_addr_127; // @[d_cache.scala 121:33 24:30]
  wire  _GEN_2954 = way1_hit ? _GEN_2057 : dirty_1_0; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2955 = way1_hit ? _GEN_2058 : dirty_1_1; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2956 = way1_hit ? _GEN_2059 : dirty_1_2; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2957 = way1_hit ? _GEN_2060 : dirty_1_3; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2958 = way1_hit ? _GEN_2061 : dirty_1_4; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2959 = way1_hit ? _GEN_2062 : dirty_1_5; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2960 = way1_hit ? _GEN_2063 : dirty_1_6; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2961 = way1_hit ? _GEN_2064 : dirty_1_7; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2962 = way1_hit ? _GEN_2065 : dirty_1_8; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2963 = way1_hit ? _GEN_2066 : dirty_1_9; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2964 = way1_hit ? _GEN_2067 : dirty_1_10; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2965 = way1_hit ? _GEN_2068 : dirty_1_11; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2966 = way1_hit ? _GEN_2069 : dirty_1_12; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2967 = way1_hit ? _GEN_2070 : dirty_1_13; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2968 = way1_hit ? _GEN_2071 : dirty_1_14; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2969 = way1_hit ? _GEN_2072 : dirty_1_15; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2970 = way1_hit ? _GEN_2073 : dirty_1_16; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2971 = way1_hit ? _GEN_2074 : dirty_1_17; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2972 = way1_hit ? _GEN_2075 : dirty_1_18; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2973 = way1_hit ? _GEN_2076 : dirty_1_19; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2974 = way1_hit ? _GEN_2077 : dirty_1_20; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2975 = way1_hit ? _GEN_2078 : dirty_1_21; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2976 = way1_hit ? _GEN_2079 : dirty_1_22; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2977 = way1_hit ? _GEN_2080 : dirty_1_23; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2978 = way1_hit ? _GEN_2081 : dirty_1_24; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2979 = way1_hit ? _GEN_2082 : dirty_1_25; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2980 = way1_hit ? _GEN_2083 : dirty_1_26; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2981 = way1_hit ? _GEN_2084 : dirty_1_27; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2982 = way1_hit ? _GEN_2085 : dirty_1_28; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2983 = way1_hit ? _GEN_2086 : dirty_1_29; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2984 = way1_hit ? _GEN_2087 : dirty_1_30; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2985 = way1_hit ? _GEN_2088 : dirty_1_31; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2986 = way1_hit ? _GEN_2089 : dirty_1_32; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2987 = way1_hit ? _GEN_2090 : dirty_1_33; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2988 = way1_hit ? _GEN_2091 : dirty_1_34; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2989 = way1_hit ? _GEN_2092 : dirty_1_35; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2990 = way1_hit ? _GEN_2093 : dirty_1_36; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2991 = way1_hit ? _GEN_2094 : dirty_1_37; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2992 = way1_hit ? _GEN_2095 : dirty_1_38; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2993 = way1_hit ? _GEN_2096 : dirty_1_39; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2994 = way1_hit ? _GEN_2097 : dirty_1_40; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2995 = way1_hit ? _GEN_2098 : dirty_1_41; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2996 = way1_hit ? _GEN_2099 : dirty_1_42; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2997 = way1_hit ? _GEN_2100 : dirty_1_43; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2998 = way1_hit ? _GEN_2101 : dirty_1_44; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_2999 = way1_hit ? _GEN_2102 : dirty_1_45; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3000 = way1_hit ? _GEN_2103 : dirty_1_46; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3001 = way1_hit ? _GEN_2104 : dirty_1_47; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3002 = way1_hit ? _GEN_2105 : dirty_1_48; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3003 = way1_hit ? _GEN_2106 : dirty_1_49; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3004 = way1_hit ? _GEN_2107 : dirty_1_50; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3005 = way1_hit ? _GEN_2108 : dirty_1_51; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3006 = way1_hit ? _GEN_2109 : dirty_1_52; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3007 = way1_hit ? _GEN_2110 : dirty_1_53; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3008 = way1_hit ? _GEN_2111 : dirty_1_54; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3009 = way1_hit ? _GEN_2112 : dirty_1_55; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3010 = way1_hit ? _GEN_2113 : dirty_1_56; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3011 = way1_hit ? _GEN_2114 : dirty_1_57; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3012 = way1_hit ? _GEN_2115 : dirty_1_58; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3013 = way1_hit ? _GEN_2116 : dirty_1_59; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3014 = way1_hit ? _GEN_2117 : dirty_1_60; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3015 = way1_hit ? _GEN_2118 : dirty_1_61; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3016 = way1_hit ? _GEN_2119 : dirty_1_62; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3017 = way1_hit ? _GEN_2120 : dirty_1_63; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3018 = way1_hit ? _GEN_2121 : dirty_1_64; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3019 = way1_hit ? _GEN_2122 : dirty_1_65; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3020 = way1_hit ? _GEN_2123 : dirty_1_66; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3021 = way1_hit ? _GEN_2124 : dirty_1_67; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3022 = way1_hit ? _GEN_2125 : dirty_1_68; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3023 = way1_hit ? _GEN_2126 : dirty_1_69; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3024 = way1_hit ? _GEN_2127 : dirty_1_70; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3025 = way1_hit ? _GEN_2128 : dirty_1_71; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3026 = way1_hit ? _GEN_2129 : dirty_1_72; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3027 = way1_hit ? _GEN_2130 : dirty_1_73; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3028 = way1_hit ? _GEN_2131 : dirty_1_74; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3029 = way1_hit ? _GEN_2132 : dirty_1_75; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3030 = way1_hit ? _GEN_2133 : dirty_1_76; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3031 = way1_hit ? _GEN_2134 : dirty_1_77; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3032 = way1_hit ? _GEN_2135 : dirty_1_78; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3033 = way1_hit ? _GEN_2136 : dirty_1_79; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3034 = way1_hit ? _GEN_2137 : dirty_1_80; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3035 = way1_hit ? _GEN_2138 : dirty_1_81; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3036 = way1_hit ? _GEN_2139 : dirty_1_82; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3037 = way1_hit ? _GEN_2140 : dirty_1_83; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3038 = way1_hit ? _GEN_2141 : dirty_1_84; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3039 = way1_hit ? _GEN_2142 : dirty_1_85; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3040 = way1_hit ? _GEN_2143 : dirty_1_86; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3041 = way1_hit ? _GEN_2144 : dirty_1_87; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3042 = way1_hit ? _GEN_2145 : dirty_1_88; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3043 = way1_hit ? _GEN_2146 : dirty_1_89; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3044 = way1_hit ? _GEN_2147 : dirty_1_90; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3045 = way1_hit ? _GEN_2148 : dirty_1_91; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3046 = way1_hit ? _GEN_2149 : dirty_1_92; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3047 = way1_hit ? _GEN_2150 : dirty_1_93; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3048 = way1_hit ? _GEN_2151 : dirty_1_94; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3049 = way1_hit ? _GEN_2152 : dirty_1_95; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3050 = way1_hit ? _GEN_2153 : dirty_1_96; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3051 = way1_hit ? _GEN_2154 : dirty_1_97; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3052 = way1_hit ? _GEN_2155 : dirty_1_98; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3053 = way1_hit ? _GEN_2156 : dirty_1_99; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3054 = way1_hit ? _GEN_2157 : dirty_1_100; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3055 = way1_hit ? _GEN_2158 : dirty_1_101; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3056 = way1_hit ? _GEN_2159 : dirty_1_102; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3057 = way1_hit ? _GEN_2160 : dirty_1_103; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3058 = way1_hit ? _GEN_2161 : dirty_1_104; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3059 = way1_hit ? _GEN_2162 : dirty_1_105; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3060 = way1_hit ? _GEN_2163 : dirty_1_106; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3061 = way1_hit ? _GEN_2164 : dirty_1_107; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3062 = way1_hit ? _GEN_2165 : dirty_1_108; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3063 = way1_hit ? _GEN_2166 : dirty_1_109; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3064 = way1_hit ? _GEN_2167 : dirty_1_110; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3065 = way1_hit ? _GEN_2168 : dirty_1_111; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3066 = way1_hit ? _GEN_2169 : dirty_1_112; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3067 = way1_hit ? _GEN_2170 : dirty_1_113; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3068 = way1_hit ? _GEN_2171 : dirty_1_114; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3069 = way1_hit ? _GEN_2172 : dirty_1_115; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3070 = way1_hit ? _GEN_2173 : dirty_1_116; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3071 = way1_hit ? _GEN_2174 : dirty_1_117; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3072 = way1_hit ? _GEN_2175 : dirty_1_118; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3073 = way1_hit ? _GEN_2176 : dirty_1_119; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3074 = way1_hit ? _GEN_2177 : dirty_1_120; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3075 = way1_hit ? _GEN_2178 : dirty_1_121; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3076 = way1_hit ? _GEN_2179 : dirty_1_122; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3077 = way1_hit ? _GEN_2180 : dirty_1_123; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3078 = way1_hit ? _GEN_2181 : dirty_1_124; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3079 = way1_hit ? _GEN_2182 : dirty_1_125; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3080 = way1_hit ? _GEN_2183 : dirty_1_126; // @[d_cache.scala 121:33 33:26]
  wire  _GEN_3081 = way1_hit ? _GEN_2184 : dirty_1_127; // @[d_cache.scala 121:33 33:26]
  wire [2:0] _GEN_3082 = way0_hit ? 3'h0 : _GEN_2185; // @[d_cache.scala 113:27 114:23]
  wire [63:0] _GEN_3083 = way0_hit ? _GEN_905 : ram_0_0; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3084 = way0_hit ? _GEN_906 : ram_0_1; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3085 = way0_hit ? _GEN_907 : ram_0_2; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3086 = way0_hit ? _GEN_908 : ram_0_3; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3087 = way0_hit ? _GEN_909 : ram_0_4; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3088 = way0_hit ? _GEN_910 : ram_0_5; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3089 = way0_hit ? _GEN_911 : ram_0_6; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3090 = way0_hit ? _GEN_912 : ram_0_7; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3091 = way0_hit ? _GEN_913 : ram_0_8; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3092 = way0_hit ? _GEN_914 : ram_0_9; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3093 = way0_hit ? _GEN_915 : ram_0_10; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3094 = way0_hit ? _GEN_916 : ram_0_11; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3095 = way0_hit ? _GEN_917 : ram_0_12; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3096 = way0_hit ? _GEN_918 : ram_0_13; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3097 = way0_hit ? _GEN_919 : ram_0_14; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3098 = way0_hit ? _GEN_920 : ram_0_15; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3099 = way0_hit ? _GEN_921 : ram_0_16; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3100 = way0_hit ? _GEN_922 : ram_0_17; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3101 = way0_hit ? _GEN_923 : ram_0_18; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3102 = way0_hit ? _GEN_924 : ram_0_19; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3103 = way0_hit ? _GEN_925 : ram_0_20; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3104 = way0_hit ? _GEN_926 : ram_0_21; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3105 = way0_hit ? _GEN_927 : ram_0_22; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3106 = way0_hit ? _GEN_928 : ram_0_23; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3107 = way0_hit ? _GEN_929 : ram_0_24; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3108 = way0_hit ? _GEN_930 : ram_0_25; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3109 = way0_hit ? _GEN_931 : ram_0_26; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3110 = way0_hit ? _GEN_932 : ram_0_27; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3111 = way0_hit ? _GEN_933 : ram_0_28; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3112 = way0_hit ? _GEN_934 : ram_0_29; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3113 = way0_hit ? _GEN_935 : ram_0_30; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3114 = way0_hit ? _GEN_936 : ram_0_31; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3115 = way0_hit ? _GEN_937 : ram_0_32; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3116 = way0_hit ? _GEN_938 : ram_0_33; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3117 = way0_hit ? _GEN_939 : ram_0_34; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3118 = way0_hit ? _GEN_940 : ram_0_35; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3119 = way0_hit ? _GEN_941 : ram_0_36; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3120 = way0_hit ? _GEN_942 : ram_0_37; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3121 = way0_hit ? _GEN_943 : ram_0_38; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3122 = way0_hit ? _GEN_944 : ram_0_39; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3123 = way0_hit ? _GEN_945 : ram_0_40; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3124 = way0_hit ? _GEN_946 : ram_0_41; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3125 = way0_hit ? _GEN_947 : ram_0_42; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3126 = way0_hit ? _GEN_948 : ram_0_43; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3127 = way0_hit ? _GEN_949 : ram_0_44; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3128 = way0_hit ? _GEN_950 : ram_0_45; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3129 = way0_hit ? _GEN_951 : ram_0_46; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3130 = way0_hit ? _GEN_952 : ram_0_47; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3131 = way0_hit ? _GEN_953 : ram_0_48; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3132 = way0_hit ? _GEN_954 : ram_0_49; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3133 = way0_hit ? _GEN_955 : ram_0_50; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3134 = way0_hit ? _GEN_956 : ram_0_51; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3135 = way0_hit ? _GEN_957 : ram_0_52; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3136 = way0_hit ? _GEN_958 : ram_0_53; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3137 = way0_hit ? _GEN_959 : ram_0_54; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3138 = way0_hit ? _GEN_960 : ram_0_55; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3139 = way0_hit ? _GEN_961 : ram_0_56; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3140 = way0_hit ? _GEN_962 : ram_0_57; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3141 = way0_hit ? _GEN_963 : ram_0_58; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3142 = way0_hit ? _GEN_964 : ram_0_59; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3143 = way0_hit ? _GEN_965 : ram_0_60; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3144 = way0_hit ? _GEN_966 : ram_0_61; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3145 = way0_hit ? _GEN_967 : ram_0_62; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3146 = way0_hit ? _GEN_968 : ram_0_63; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3147 = way0_hit ? _GEN_969 : ram_0_64; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3148 = way0_hit ? _GEN_970 : ram_0_65; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3149 = way0_hit ? _GEN_971 : ram_0_66; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3150 = way0_hit ? _GEN_972 : ram_0_67; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3151 = way0_hit ? _GEN_973 : ram_0_68; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3152 = way0_hit ? _GEN_974 : ram_0_69; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3153 = way0_hit ? _GEN_975 : ram_0_70; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3154 = way0_hit ? _GEN_976 : ram_0_71; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3155 = way0_hit ? _GEN_977 : ram_0_72; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3156 = way0_hit ? _GEN_978 : ram_0_73; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3157 = way0_hit ? _GEN_979 : ram_0_74; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3158 = way0_hit ? _GEN_980 : ram_0_75; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3159 = way0_hit ? _GEN_981 : ram_0_76; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3160 = way0_hit ? _GEN_982 : ram_0_77; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3161 = way0_hit ? _GEN_983 : ram_0_78; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3162 = way0_hit ? _GEN_984 : ram_0_79; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3163 = way0_hit ? _GEN_985 : ram_0_80; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3164 = way0_hit ? _GEN_986 : ram_0_81; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3165 = way0_hit ? _GEN_987 : ram_0_82; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3166 = way0_hit ? _GEN_988 : ram_0_83; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3167 = way0_hit ? _GEN_989 : ram_0_84; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3168 = way0_hit ? _GEN_990 : ram_0_85; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3169 = way0_hit ? _GEN_991 : ram_0_86; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3170 = way0_hit ? _GEN_992 : ram_0_87; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3171 = way0_hit ? _GEN_993 : ram_0_88; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3172 = way0_hit ? _GEN_994 : ram_0_89; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3173 = way0_hit ? _GEN_995 : ram_0_90; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3174 = way0_hit ? _GEN_996 : ram_0_91; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3175 = way0_hit ? _GEN_997 : ram_0_92; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3176 = way0_hit ? _GEN_998 : ram_0_93; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3177 = way0_hit ? _GEN_999 : ram_0_94; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3178 = way0_hit ? _GEN_1000 : ram_0_95; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3179 = way0_hit ? _GEN_1001 : ram_0_96; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3180 = way0_hit ? _GEN_1002 : ram_0_97; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3181 = way0_hit ? _GEN_1003 : ram_0_98; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3182 = way0_hit ? _GEN_1004 : ram_0_99; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3183 = way0_hit ? _GEN_1005 : ram_0_100; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3184 = way0_hit ? _GEN_1006 : ram_0_101; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3185 = way0_hit ? _GEN_1007 : ram_0_102; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3186 = way0_hit ? _GEN_1008 : ram_0_103; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3187 = way0_hit ? _GEN_1009 : ram_0_104; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3188 = way0_hit ? _GEN_1010 : ram_0_105; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3189 = way0_hit ? _GEN_1011 : ram_0_106; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3190 = way0_hit ? _GEN_1012 : ram_0_107; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3191 = way0_hit ? _GEN_1013 : ram_0_108; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3192 = way0_hit ? _GEN_1014 : ram_0_109; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3193 = way0_hit ? _GEN_1015 : ram_0_110; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3194 = way0_hit ? _GEN_1016 : ram_0_111; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3195 = way0_hit ? _GEN_1017 : ram_0_112; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3196 = way0_hit ? _GEN_1018 : ram_0_113; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3197 = way0_hit ? _GEN_1019 : ram_0_114; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3198 = way0_hit ? _GEN_1020 : ram_0_115; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3199 = way0_hit ? _GEN_1021 : ram_0_116; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3200 = way0_hit ? _GEN_1022 : ram_0_117; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3201 = way0_hit ? _GEN_1023 : ram_0_118; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3202 = way0_hit ? _GEN_1024 : ram_0_119; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3203 = way0_hit ? _GEN_1025 : ram_0_120; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3204 = way0_hit ? _GEN_1026 : ram_0_121; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3205 = way0_hit ? _GEN_1027 : ram_0_122; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3206 = way0_hit ? _GEN_1028 : ram_0_123; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3207 = way0_hit ? _GEN_1029 : ram_0_124; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3208 = way0_hit ? _GEN_1030 : ram_0_125; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3209 = way0_hit ? _GEN_1031 : ram_0_126; // @[d_cache.scala 113:27 19:24]
  wire [63:0] _GEN_3210 = way0_hit ? _GEN_1032 : ram_0_127; // @[d_cache.scala 113:27 19:24]
  wire  _GEN_3211 = way0_hit ? _GEN_1033 : dirty_0_0; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3212 = way0_hit ? _GEN_1034 : dirty_0_1; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3213 = way0_hit ? _GEN_1035 : dirty_0_2; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3214 = way0_hit ? _GEN_1036 : dirty_0_3; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3215 = way0_hit ? _GEN_1037 : dirty_0_4; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3216 = way0_hit ? _GEN_1038 : dirty_0_5; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3217 = way0_hit ? _GEN_1039 : dirty_0_6; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3218 = way0_hit ? _GEN_1040 : dirty_0_7; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3219 = way0_hit ? _GEN_1041 : dirty_0_8; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3220 = way0_hit ? _GEN_1042 : dirty_0_9; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3221 = way0_hit ? _GEN_1043 : dirty_0_10; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3222 = way0_hit ? _GEN_1044 : dirty_0_11; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3223 = way0_hit ? _GEN_1045 : dirty_0_12; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3224 = way0_hit ? _GEN_1046 : dirty_0_13; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3225 = way0_hit ? _GEN_1047 : dirty_0_14; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3226 = way0_hit ? _GEN_1048 : dirty_0_15; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3227 = way0_hit ? _GEN_1049 : dirty_0_16; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3228 = way0_hit ? _GEN_1050 : dirty_0_17; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3229 = way0_hit ? _GEN_1051 : dirty_0_18; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3230 = way0_hit ? _GEN_1052 : dirty_0_19; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3231 = way0_hit ? _GEN_1053 : dirty_0_20; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3232 = way0_hit ? _GEN_1054 : dirty_0_21; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3233 = way0_hit ? _GEN_1055 : dirty_0_22; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3234 = way0_hit ? _GEN_1056 : dirty_0_23; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3235 = way0_hit ? _GEN_1057 : dirty_0_24; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3236 = way0_hit ? _GEN_1058 : dirty_0_25; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3237 = way0_hit ? _GEN_1059 : dirty_0_26; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3238 = way0_hit ? _GEN_1060 : dirty_0_27; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3239 = way0_hit ? _GEN_1061 : dirty_0_28; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3240 = way0_hit ? _GEN_1062 : dirty_0_29; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3241 = way0_hit ? _GEN_1063 : dirty_0_30; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3242 = way0_hit ? _GEN_1064 : dirty_0_31; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3243 = way0_hit ? _GEN_1065 : dirty_0_32; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3244 = way0_hit ? _GEN_1066 : dirty_0_33; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3245 = way0_hit ? _GEN_1067 : dirty_0_34; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3246 = way0_hit ? _GEN_1068 : dirty_0_35; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3247 = way0_hit ? _GEN_1069 : dirty_0_36; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3248 = way0_hit ? _GEN_1070 : dirty_0_37; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3249 = way0_hit ? _GEN_1071 : dirty_0_38; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3250 = way0_hit ? _GEN_1072 : dirty_0_39; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3251 = way0_hit ? _GEN_1073 : dirty_0_40; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3252 = way0_hit ? _GEN_1074 : dirty_0_41; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3253 = way0_hit ? _GEN_1075 : dirty_0_42; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3254 = way0_hit ? _GEN_1076 : dirty_0_43; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3255 = way0_hit ? _GEN_1077 : dirty_0_44; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3256 = way0_hit ? _GEN_1078 : dirty_0_45; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3257 = way0_hit ? _GEN_1079 : dirty_0_46; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3258 = way0_hit ? _GEN_1080 : dirty_0_47; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3259 = way0_hit ? _GEN_1081 : dirty_0_48; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3260 = way0_hit ? _GEN_1082 : dirty_0_49; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3261 = way0_hit ? _GEN_1083 : dirty_0_50; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3262 = way0_hit ? _GEN_1084 : dirty_0_51; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3263 = way0_hit ? _GEN_1085 : dirty_0_52; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3264 = way0_hit ? _GEN_1086 : dirty_0_53; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3265 = way0_hit ? _GEN_1087 : dirty_0_54; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3266 = way0_hit ? _GEN_1088 : dirty_0_55; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3267 = way0_hit ? _GEN_1089 : dirty_0_56; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3268 = way0_hit ? _GEN_1090 : dirty_0_57; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3269 = way0_hit ? _GEN_1091 : dirty_0_58; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3270 = way0_hit ? _GEN_1092 : dirty_0_59; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3271 = way0_hit ? _GEN_1093 : dirty_0_60; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3272 = way0_hit ? _GEN_1094 : dirty_0_61; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3273 = way0_hit ? _GEN_1095 : dirty_0_62; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3274 = way0_hit ? _GEN_1096 : dirty_0_63; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3275 = way0_hit ? _GEN_1097 : dirty_0_64; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3276 = way0_hit ? _GEN_1098 : dirty_0_65; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3277 = way0_hit ? _GEN_1099 : dirty_0_66; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3278 = way0_hit ? _GEN_1100 : dirty_0_67; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3279 = way0_hit ? _GEN_1101 : dirty_0_68; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3280 = way0_hit ? _GEN_1102 : dirty_0_69; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3281 = way0_hit ? _GEN_1103 : dirty_0_70; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3282 = way0_hit ? _GEN_1104 : dirty_0_71; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3283 = way0_hit ? _GEN_1105 : dirty_0_72; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3284 = way0_hit ? _GEN_1106 : dirty_0_73; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3285 = way0_hit ? _GEN_1107 : dirty_0_74; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3286 = way0_hit ? _GEN_1108 : dirty_0_75; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3287 = way0_hit ? _GEN_1109 : dirty_0_76; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3288 = way0_hit ? _GEN_1110 : dirty_0_77; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3289 = way0_hit ? _GEN_1111 : dirty_0_78; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3290 = way0_hit ? _GEN_1112 : dirty_0_79; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3291 = way0_hit ? _GEN_1113 : dirty_0_80; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3292 = way0_hit ? _GEN_1114 : dirty_0_81; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3293 = way0_hit ? _GEN_1115 : dirty_0_82; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3294 = way0_hit ? _GEN_1116 : dirty_0_83; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3295 = way0_hit ? _GEN_1117 : dirty_0_84; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3296 = way0_hit ? _GEN_1118 : dirty_0_85; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3297 = way0_hit ? _GEN_1119 : dirty_0_86; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3298 = way0_hit ? _GEN_1120 : dirty_0_87; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3299 = way0_hit ? _GEN_1121 : dirty_0_88; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3300 = way0_hit ? _GEN_1122 : dirty_0_89; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3301 = way0_hit ? _GEN_1123 : dirty_0_90; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3302 = way0_hit ? _GEN_1124 : dirty_0_91; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3303 = way0_hit ? _GEN_1125 : dirty_0_92; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3304 = way0_hit ? _GEN_1126 : dirty_0_93; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3305 = way0_hit ? _GEN_1127 : dirty_0_94; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3306 = way0_hit ? _GEN_1128 : dirty_0_95; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3307 = way0_hit ? _GEN_1129 : dirty_0_96; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3308 = way0_hit ? _GEN_1130 : dirty_0_97; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3309 = way0_hit ? _GEN_1131 : dirty_0_98; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3310 = way0_hit ? _GEN_1132 : dirty_0_99; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3311 = way0_hit ? _GEN_1133 : dirty_0_100; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3312 = way0_hit ? _GEN_1134 : dirty_0_101; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3313 = way0_hit ? _GEN_1135 : dirty_0_102; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3314 = way0_hit ? _GEN_1136 : dirty_0_103; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3315 = way0_hit ? _GEN_1137 : dirty_0_104; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3316 = way0_hit ? _GEN_1138 : dirty_0_105; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3317 = way0_hit ? _GEN_1139 : dirty_0_106; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3318 = way0_hit ? _GEN_1140 : dirty_0_107; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3319 = way0_hit ? _GEN_1141 : dirty_0_108; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3320 = way0_hit ? _GEN_1142 : dirty_0_109; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3321 = way0_hit ? _GEN_1143 : dirty_0_110; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3322 = way0_hit ? _GEN_1144 : dirty_0_111; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3323 = way0_hit ? _GEN_1145 : dirty_0_112; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3324 = way0_hit ? _GEN_1146 : dirty_0_113; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3325 = way0_hit ? _GEN_1147 : dirty_0_114; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3326 = way0_hit ? _GEN_1148 : dirty_0_115; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3327 = way0_hit ? _GEN_1149 : dirty_0_116; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3328 = way0_hit ? _GEN_1150 : dirty_0_117; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3329 = way0_hit ? _GEN_1151 : dirty_0_118; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3330 = way0_hit ? _GEN_1152 : dirty_0_119; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3331 = way0_hit ? _GEN_1153 : dirty_0_120; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3332 = way0_hit ? _GEN_1154 : dirty_0_121; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3333 = way0_hit ? _GEN_1155 : dirty_0_122; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3334 = way0_hit ? _GEN_1156 : dirty_0_123; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3335 = way0_hit ? _GEN_1157 : dirty_0_124; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3336 = way0_hit ? _GEN_1158 : dirty_0_125; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3337 = way0_hit ? _GEN_1159 : dirty_0_126; // @[d_cache.scala 113:27 32:26]
  wire  _GEN_3338 = way0_hit ? _GEN_1160 : dirty_0_127; // @[d_cache.scala 113:27 32:26]
  wire [63:0] _GEN_3339 = way0_hit ? record_olddata_0 : _GEN_2186; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3340 = way0_hit ? record_olddata_1 : _GEN_2187; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3341 = way0_hit ? record_olddata_2 : _GEN_2188; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3342 = way0_hit ? record_olddata_3 : _GEN_2189; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3343 = way0_hit ? record_olddata_4 : _GEN_2190; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3344 = way0_hit ? record_olddata_5 : _GEN_2191; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3345 = way0_hit ? record_olddata_6 : _GEN_2192; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3346 = way0_hit ? record_olddata_7 : _GEN_2193; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3347 = way0_hit ? record_olddata_8 : _GEN_2194; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3348 = way0_hit ? record_olddata_9 : _GEN_2195; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3349 = way0_hit ? record_olddata_10 : _GEN_2196; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3350 = way0_hit ? record_olddata_11 : _GEN_2197; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3351 = way0_hit ? record_olddata_12 : _GEN_2198; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3352 = way0_hit ? record_olddata_13 : _GEN_2199; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3353 = way0_hit ? record_olddata_14 : _GEN_2200; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3354 = way0_hit ? record_olddata_15 : _GEN_2201; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3355 = way0_hit ? record_olddata_16 : _GEN_2202; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3356 = way0_hit ? record_olddata_17 : _GEN_2203; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3357 = way0_hit ? record_olddata_18 : _GEN_2204; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3358 = way0_hit ? record_olddata_19 : _GEN_2205; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3359 = way0_hit ? record_olddata_20 : _GEN_2206; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3360 = way0_hit ? record_olddata_21 : _GEN_2207; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3361 = way0_hit ? record_olddata_22 : _GEN_2208; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3362 = way0_hit ? record_olddata_23 : _GEN_2209; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3363 = way0_hit ? record_olddata_24 : _GEN_2210; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3364 = way0_hit ? record_olddata_25 : _GEN_2211; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3365 = way0_hit ? record_olddata_26 : _GEN_2212; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3366 = way0_hit ? record_olddata_27 : _GEN_2213; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3367 = way0_hit ? record_olddata_28 : _GEN_2214; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3368 = way0_hit ? record_olddata_29 : _GEN_2215; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3369 = way0_hit ? record_olddata_30 : _GEN_2216; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3370 = way0_hit ? record_olddata_31 : _GEN_2217; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3371 = way0_hit ? record_olddata_32 : _GEN_2218; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3372 = way0_hit ? record_olddata_33 : _GEN_2219; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3373 = way0_hit ? record_olddata_34 : _GEN_2220; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3374 = way0_hit ? record_olddata_35 : _GEN_2221; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3375 = way0_hit ? record_olddata_36 : _GEN_2222; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3376 = way0_hit ? record_olddata_37 : _GEN_2223; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3377 = way0_hit ? record_olddata_38 : _GEN_2224; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3378 = way0_hit ? record_olddata_39 : _GEN_2225; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3379 = way0_hit ? record_olddata_40 : _GEN_2226; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3380 = way0_hit ? record_olddata_41 : _GEN_2227; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3381 = way0_hit ? record_olddata_42 : _GEN_2228; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3382 = way0_hit ? record_olddata_43 : _GEN_2229; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3383 = way0_hit ? record_olddata_44 : _GEN_2230; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3384 = way0_hit ? record_olddata_45 : _GEN_2231; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3385 = way0_hit ? record_olddata_46 : _GEN_2232; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3386 = way0_hit ? record_olddata_47 : _GEN_2233; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3387 = way0_hit ? record_olddata_48 : _GEN_2234; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3388 = way0_hit ? record_olddata_49 : _GEN_2235; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3389 = way0_hit ? record_olddata_50 : _GEN_2236; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3390 = way0_hit ? record_olddata_51 : _GEN_2237; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3391 = way0_hit ? record_olddata_52 : _GEN_2238; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3392 = way0_hit ? record_olddata_53 : _GEN_2239; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3393 = way0_hit ? record_olddata_54 : _GEN_2240; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3394 = way0_hit ? record_olddata_55 : _GEN_2241; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3395 = way0_hit ? record_olddata_56 : _GEN_2242; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3396 = way0_hit ? record_olddata_57 : _GEN_2243; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3397 = way0_hit ? record_olddata_58 : _GEN_2244; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3398 = way0_hit ? record_olddata_59 : _GEN_2245; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3399 = way0_hit ? record_olddata_60 : _GEN_2246; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3400 = way0_hit ? record_olddata_61 : _GEN_2247; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3401 = way0_hit ? record_olddata_62 : _GEN_2248; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3402 = way0_hit ? record_olddata_63 : _GEN_2249; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3403 = way0_hit ? record_olddata_64 : _GEN_2250; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3404 = way0_hit ? record_olddata_65 : _GEN_2251; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3405 = way0_hit ? record_olddata_66 : _GEN_2252; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3406 = way0_hit ? record_olddata_67 : _GEN_2253; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3407 = way0_hit ? record_olddata_68 : _GEN_2254; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3408 = way0_hit ? record_olddata_69 : _GEN_2255; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3409 = way0_hit ? record_olddata_70 : _GEN_2256; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3410 = way0_hit ? record_olddata_71 : _GEN_2257; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3411 = way0_hit ? record_olddata_72 : _GEN_2258; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3412 = way0_hit ? record_olddata_73 : _GEN_2259; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3413 = way0_hit ? record_olddata_74 : _GEN_2260; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3414 = way0_hit ? record_olddata_75 : _GEN_2261; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3415 = way0_hit ? record_olddata_76 : _GEN_2262; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3416 = way0_hit ? record_olddata_77 : _GEN_2263; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3417 = way0_hit ? record_olddata_78 : _GEN_2264; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3418 = way0_hit ? record_olddata_79 : _GEN_2265; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3419 = way0_hit ? record_olddata_80 : _GEN_2266; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3420 = way0_hit ? record_olddata_81 : _GEN_2267; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3421 = way0_hit ? record_olddata_82 : _GEN_2268; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3422 = way0_hit ? record_olddata_83 : _GEN_2269; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3423 = way0_hit ? record_olddata_84 : _GEN_2270; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3424 = way0_hit ? record_olddata_85 : _GEN_2271; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3425 = way0_hit ? record_olddata_86 : _GEN_2272; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3426 = way0_hit ? record_olddata_87 : _GEN_2273; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3427 = way0_hit ? record_olddata_88 : _GEN_2274; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3428 = way0_hit ? record_olddata_89 : _GEN_2275; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3429 = way0_hit ? record_olddata_90 : _GEN_2276; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3430 = way0_hit ? record_olddata_91 : _GEN_2277; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3431 = way0_hit ? record_olddata_92 : _GEN_2278; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3432 = way0_hit ? record_olddata_93 : _GEN_2279; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3433 = way0_hit ? record_olddata_94 : _GEN_2280; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3434 = way0_hit ? record_olddata_95 : _GEN_2281; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3435 = way0_hit ? record_olddata_96 : _GEN_2282; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3436 = way0_hit ? record_olddata_97 : _GEN_2283; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3437 = way0_hit ? record_olddata_98 : _GEN_2284; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3438 = way0_hit ? record_olddata_99 : _GEN_2285; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3439 = way0_hit ? record_olddata_100 : _GEN_2286; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3440 = way0_hit ? record_olddata_101 : _GEN_2287; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3441 = way0_hit ? record_olddata_102 : _GEN_2288; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3442 = way0_hit ? record_olddata_103 : _GEN_2289; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3443 = way0_hit ? record_olddata_104 : _GEN_2290; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3444 = way0_hit ? record_olddata_105 : _GEN_2291; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3445 = way0_hit ? record_olddata_106 : _GEN_2292; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3446 = way0_hit ? record_olddata_107 : _GEN_2293; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3447 = way0_hit ? record_olddata_108 : _GEN_2294; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3448 = way0_hit ? record_olddata_109 : _GEN_2295; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3449 = way0_hit ? record_olddata_110 : _GEN_2296; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3450 = way0_hit ? record_olddata_111 : _GEN_2297; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3451 = way0_hit ? record_olddata_112 : _GEN_2298; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3452 = way0_hit ? record_olddata_113 : _GEN_2299; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3453 = way0_hit ? record_olddata_114 : _GEN_2300; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3454 = way0_hit ? record_olddata_115 : _GEN_2301; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3455 = way0_hit ? record_olddata_116 : _GEN_2302; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3456 = way0_hit ? record_olddata_117 : _GEN_2303; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3457 = way0_hit ? record_olddata_118 : _GEN_2304; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3458 = way0_hit ? record_olddata_119 : _GEN_2305; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3459 = way0_hit ? record_olddata_120 : _GEN_2306; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3460 = way0_hit ? record_olddata_121 : _GEN_2307; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3461 = way0_hit ? record_olddata_122 : _GEN_2308; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3462 = way0_hit ? record_olddata_123 : _GEN_2309; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3463 = way0_hit ? record_olddata_124 : _GEN_2310; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3464 = way0_hit ? record_olddata_125 : _GEN_2311; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3465 = way0_hit ? record_olddata_126 : _GEN_2312; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3466 = way0_hit ? record_olddata_127 : _GEN_2313; // @[d_cache.scala 113:27 25:33]
  wire [63:0] _GEN_3467 = way0_hit ? ram_1_0 : _GEN_2314; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3468 = way0_hit ? ram_1_1 : _GEN_2315; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3469 = way0_hit ? ram_1_2 : _GEN_2316; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3470 = way0_hit ? ram_1_3 : _GEN_2317; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3471 = way0_hit ? ram_1_4 : _GEN_2318; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3472 = way0_hit ? ram_1_5 : _GEN_2319; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3473 = way0_hit ? ram_1_6 : _GEN_2320; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3474 = way0_hit ? ram_1_7 : _GEN_2321; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3475 = way0_hit ? ram_1_8 : _GEN_2322; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3476 = way0_hit ? ram_1_9 : _GEN_2323; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3477 = way0_hit ? ram_1_10 : _GEN_2324; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3478 = way0_hit ? ram_1_11 : _GEN_2325; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3479 = way0_hit ? ram_1_12 : _GEN_2326; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3480 = way0_hit ? ram_1_13 : _GEN_2327; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3481 = way0_hit ? ram_1_14 : _GEN_2328; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3482 = way0_hit ? ram_1_15 : _GEN_2329; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3483 = way0_hit ? ram_1_16 : _GEN_2330; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3484 = way0_hit ? ram_1_17 : _GEN_2331; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3485 = way0_hit ? ram_1_18 : _GEN_2332; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3486 = way0_hit ? ram_1_19 : _GEN_2333; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3487 = way0_hit ? ram_1_20 : _GEN_2334; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3488 = way0_hit ? ram_1_21 : _GEN_2335; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3489 = way0_hit ? ram_1_22 : _GEN_2336; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3490 = way0_hit ? ram_1_23 : _GEN_2337; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3491 = way0_hit ? ram_1_24 : _GEN_2338; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3492 = way0_hit ? ram_1_25 : _GEN_2339; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3493 = way0_hit ? ram_1_26 : _GEN_2340; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3494 = way0_hit ? ram_1_27 : _GEN_2341; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3495 = way0_hit ? ram_1_28 : _GEN_2342; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3496 = way0_hit ? ram_1_29 : _GEN_2343; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3497 = way0_hit ? ram_1_30 : _GEN_2344; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3498 = way0_hit ? ram_1_31 : _GEN_2345; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3499 = way0_hit ? ram_1_32 : _GEN_2346; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3500 = way0_hit ? ram_1_33 : _GEN_2347; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3501 = way0_hit ? ram_1_34 : _GEN_2348; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3502 = way0_hit ? ram_1_35 : _GEN_2349; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3503 = way0_hit ? ram_1_36 : _GEN_2350; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3504 = way0_hit ? ram_1_37 : _GEN_2351; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3505 = way0_hit ? ram_1_38 : _GEN_2352; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3506 = way0_hit ? ram_1_39 : _GEN_2353; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3507 = way0_hit ? ram_1_40 : _GEN_2354; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3508 = way0_hit ? ram_1_41 : _GEN_2355; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3509 = way0_hit ? ram_1_42 : _GEN_2356; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3510 = way0_hit ? ram_1_43 : _GEN_2357; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3511 = way0_hit ? ram_1_44 : _GEN_2358; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3512 = way0_hit ? ram_1_45 : _GEN_2359; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3513 = way0_hit ? ram_1_46 : _GEN_2360; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3514 = way0_hit ? ram_1_47 : _GEN_2361; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3515 = way0_hit ? ram_1_48 : _GEN_2362; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3516 = way0_hit ? ram_1_49 : _GEN_2363; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3517 = way0_hit ? ram_1_50 : _GEN_2364; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3518 = way0_hit ? ram_1_51 : _GEN_2365; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3519 = way0_hit ? ram_1_52 : _GEN_2366; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3520 = way0_hit ? ram_1_53 : _GEN_2367; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3521 = way0_hit ? ram_1_54 : _GEN_2368; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3522 = way0_hit ? ram_1_55 : _GEN_2369; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3523 = way0_hit ? ram_1_56 : _GEN_2370; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3524 = way0_hit ? ram_1_57 : _GEN_2371; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3525 = way0_hit ? ram_1_58 : _GEN_2372; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3526 = way0_hit ? ram_1_59 : _GEN_2373; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3527 = way0_hit ? ram_1_60 : _GEN_2374; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3528 = way0_hit ? ram_1_61 : _GEN_2375; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3529 = way0_hit ? ram_1_62 : _GEN_2376; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3530 = way0_hit ? ram_1_63 : _GEN_2377; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3531 = way0_hit ? ram_1_64 : _GEN_2378; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3532 = way0_hit ? ram_1_65 : _GEN_2379; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3533 = way0_hit ? ram_1_66 : _GEN_2380; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3534 = way0_hit ? ram_1_67 : _GEN_2381; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3535 = way0_hit ? ram_1_68 : _GEN_2382; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3536 = way0_hit ? ram_1_69 : _GEN_2383; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3537 = way0_hit ? ram_1_70 : _GEN_2384; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3538 = way0_hit ? ram_1_71 : _GEN_2385; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3539 = way0_hit ? ram_1_72 : _GEN_2386; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3540 = way0_hit ? ram_1_73 : _GEN_2387; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3541 = way0_hit ? ram_1_74 : _GEN_2388; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3542 = way0_hit ? ram_1_75 : _GEN_2389; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3543 = way0_hit ? ram_1_76 : _GEN_2390; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3544 = way0_hit ? ram_1_77 : _GEN_2391; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3545 = way0_hit ? ram_1_78 : _GEN_2392; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3546 = way0_hit ? ram_1_79 : _GEN_2393; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3547 = way0_hit ? ram_1_80 : _GEN_2394; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3548 = way0_hit ? ram_1_81 : _GEN_2395; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3549 = way0_hit ? ram_1_82 : _GEN_2396; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3550 = way0_hit ? ram_1_83 : _GEN_2397; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3551 = way0_hit ? ram_1_84 : _GEN_2398; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3552 = way0_hit ? ram_1_85 : _GEN_2399; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3553 = way0_hit ? ram_1_86 : _GEN_2400; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3554 = way0_hit ? ram_1_87 : _GEN_2401; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3555 = way0_hit ? ram_1_88 : _GEN_2402; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3556 = way0_hit ? ram_1_89 : _GEN_2403; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3557 = way0_hit ? ram_1_90 : _GEN_2404; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3558 = way0_hit ? ram_1_91 : _GEN_2405; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3559 = way0_hit ? ram_1_92 : _GEN_2406; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3560 = way0_hit ? ram_1_93 : _GEN_2407; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3561 = way0_hit ? ram_1_94 : _GEN_2408; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3562 = way0_hit ? ram_1_95 : _GEN_2409; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3563 = way0_hit ? ram_1_96 : _GEN_2410; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3564 = way0_hit ? ram_1_97 : _GEN_2411; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3565 = way0_hit ? ram_1_98 : _GEN_2412; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3566 = way0_hit ? ram_1_99 : _GEN_2413; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3567 = way0_hit ? ram_1_100 : _GEN_2414; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3568 = way0_hit ? ram_1_101 : _GEN_2415; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3569 = way0_hit ? ram_1_102 : _GEN_2416; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3570 = way0_hit ? ram_1_103 : _GEN_2417; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3571 = way0_hit ? ram_1_104 : _GEN_2418; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3572 = way0_hit ? ram_1_105 : _GEN_2419; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3573 = way0_hit ? ram_1_106 : _GEN_2420; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3574 = way0_hit ? ram_1_107 : _GEN_2421; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3575 = way0_hit ? ram_1_108 : _GEN_2422; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3576 = way0_hit ? ram_1_109 : _GEN_2423; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3577 = way0_hit ? ram_1_110 : _GEN_2424; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3578 = way0_hit ? ram_1_111 : _GEN_2425; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3579 = way0_hit ? ram_1_112 : _GEN_2426; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3580 = way0_hit ? ram_1_113 : _GEN_2427; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3581 = way0_hit ? ram_1_114 : _GEN_2428; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3582 = way0_hit ? ram_1_115 : _GEN_2429; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3583 = way0_hit ? ram_1_116 : _GEN_2430; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3584 = way0_hit ? ram_1_117 : _GEN_2431; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3585 = way0_hit ? ram_1_118 : _GEN_2432; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3586 = way0_hit ? ram_1_119 : _GEN_2433; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3587 = way0_hit ? ram_1_120 : _GEN_2434; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3588 = way0_hit ? ram_1_121 : _GEN_2435; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3589 = way0_hit ? ram_1_122 : _GEN_2436; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3590 = way0_hit ? ram_1_123 : _GEN_2437; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3591 = way0_hit ? ram_1_124 : _GEN_2438; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3592 = way0_hit ? ram_1_125 : _GEN_2439; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3593 = way0_hit ? ram_1_126 : _GEN_2440; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3594 = way0_hit ? ram_1_127 : _GEN_2441; // @[d_cache.scala 113:27 20:24]
  wire [63:0] _GEN_3595 = way0_hit ? record_wdata1_0 : _GEN_2442; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3596 = way0_hit ? record_wdata1_1 : _GEN_2443; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3597 = way0_hit ? record_wdata1_2 : _GEN_2444; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3598 = way0_hit ? record_wdata1_3 : _GEN_2445; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3599 = way0_hit ? record_wdata1_4 : _GEN_2446; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3600 = way0_hit ? record_wdata1_5 : _GEN_2447; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3601 = way0_hit ? record_wdata1_6 : _GEN_2448; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3602 = way0_hit ? record_wdata1_7 : _GEN_2449; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3603 = way0_hit ? record_wdata1_8 : _GEN_2450; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3604 = way0_hit ? record_wdata1_9 : _GEN_2451; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3605 = way0_hit ? record_wdata1_10 : _GEN_2452; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3606 = way0_hit ? record_wdata1_11 : _GEN_2453; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3607 = way0_hit ? record_wdata1_12 : _GEN_2454; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3608 = way0_hit ? record_wdata1_13 : _GEN_2455; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3609 = way0_hit ? record_wdata1_14 : _GEN_2456; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3610 = way0_hit ? record_wdata1_15 : _GEN_2457; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3611 = way0_hit ? record_wdata1_16 : _GEN_2458; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3612 = way0_hit ? record_wdata1_17 : _GEN_2459; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3613 = way0_hit ? record_wdata1_18 : _GEN_2460; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3614 = way0_hit ? record_wdata1_19 : _GEN_2461; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3615 = way0_hit ? record_wdata1_20 : _GEN_2462; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3616 = way0_hit ? record_wdata1_21 : _GEN_2463; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3617 = way0_hit ? record_wdata1_22 : _GEN_2464; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3618 = way0_hit ? record_wdata1_23 : _GEN_2465; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3619 = way0_hit ? record_wdata1_24 : _GEN_2466; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3620 = way0_hit ? record_wdata1_25 : _GEN_2467; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3621 = way0_hit ? record_wdata1_26 : _GEN_2468; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3622 = way0_hit ? record_wdata1_27 : _GEN_2469; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3623 = way0_hit ? record_wdata1_28 : _GEN_2470; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3624 = way0_hit ? record_wdata1_29 : _GEN_2471; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3625 = way0_hit ? record_wdata1_30 : _GEN_2472; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3626 = way0_hit ? record_wdata1_31 : _GEN_2473; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3627 = way0_hit ? record_wdata1_32 : _GEN_2474; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3628 = way0_hit ? record_wdata1_33 : _GEN_2475; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3629 = way0_hit ? record_wdata1_34 : _GEN_2476; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3630 = way0_hit ? record_wdata1_35 : _GEN_2477; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3631 = way0_hit ? record_wdata1_36 : _GEN_2478; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3632 = way0_hit ? record_wdata1_37 : _GEN_2479; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3633 = way0_hit ? record_wdata1_38 : _GEN_2480; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3634 = way0_hit ? record_wdata1_39 : _GEN_2481; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3635 = way0_hit ? record_wdata1_40 : _GEN_2482; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3636 = way0_hit ? record_wdata1_41 : _GEN_2483; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3637 = way0_hit ? record_wdata1_42 : _GEN_2484; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3638 = way0_hit ? record_wdata1_43 : _GEN_2485; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3639 = way0_hit ? record_wdata1_44 : _GEN_2486; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3640 = way0_hit ? record_wdata1_45 : _GEN_2487; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3641 = way0_hit ? record_wdata1_46 : _GEN_2488; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3642 = way0_hit ? record_wdata1_47 : _GEN_2489; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3643 = way0_hit ? record_wdata1_48 : _GEN_2490; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3644 = way0_hit ? record_wdata1_49 : _GEN_2491; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3645 = way0_hit ? record_wdata1_50 : _GEN_2492; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3646 = way0_hit ? record_wdata1_51 : _GEN_2493; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3647 = way0_hit ? record_wdata1_52 : _GEN_2494; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3648 = way0_hit ? record_wdata1_53 : _GEN_2495; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3649 = way0_hit ? record_wdata1_54 : _GEN_2496; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3650 = way0_hit ? record_wdata1_55 : _GEN_2497; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3651 = way0_hit ? record_wdata1_56 : _GEN_2498; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3652 = way0_hit ? record_wdata1_57 : _GEN_2499; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3653 = way0_hit ? record_wdata1_58 : _GEN_2500; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3654 = way0_hit ? record_wdata1_59 : _GEN_2501; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3655 = way0_hit ? record_wdata1_60 : _GEN_2502; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3656 = way0_hit ? record_wdata1_61 : _GEN_2503; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3657 = way0_hit ? record_wdata1_62 : _GEN_2504; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3658 = way0_hit ? record_wdata1_63 : _GEN_2505; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3659 = way0_hit ? record_wdata1_64 : _GEN_2506; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3660 = way0_hit ? record_wdata1_65 : _GEN_2507; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3661 = way0_hit ? record_wdata1_66 : _GEN_2508; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3662 = way0_hit ? record_wdata1_67 : _GEN_2509; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3663 = way0_hit ? record_wdata1_68 : _GEN_2510; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3664 = way0_hit ? record_wdata1_69 : _GEN_2511; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3665 = way0_hit ? record_wdata1_70 : _GEN_2512; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3666 = way0_hit ? record_wdata1_71 : _GEN_2513; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3667 = way0_hit ? record_wdata1_72 : _GEN_2514; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3668 = way0_hit ? record_wdata1_73 : _GEN_2515; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3669 = way0_hit ? record_wdata1_74 : _GEN_2516; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3670 = way0_hit ? record_wdata1_75 : _GEN_2517; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3671 = way0_hit ? record_wdata1_76 : _GEN_2518; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3672 = way0_hit ? record_wdata1_77 : _GEN_2519; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3673 = way0_hit ? record_wdata1_78 : _GEN_2520; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3674 = way0_hit ? record_wdata1_79 : _GEN_2521; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3675 = way0_hit ? record_wdata1_80 : _GEN_2522; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3676 = way0_hit ? record_wdata1_81 : _GEN_2523; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3677 = way0_hit ? record_wdata1_82 : _GEN_2524; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3678 = way0_hit ? record_wdata1_83 : _GEN_2525; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3679 = way0_hit ? record_wdata1_84 : _GEN_2526; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3680 = way0_hit ? record_wdata1_85 : _GEN_2527; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3681 = way0_hit ? record_wdata1_86 : _GEN_2528; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3682 = way0_hit ? record_wdata1_87 : _GEN_2529; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3683 = way0_hit ? record_wdata1_88 : _GEN_2530; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3684 = way0_hit ? record_wdata1_89 : _GEN_2531; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3685 = way0_hit ? record_wdata1_90 : _GEN_2532; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3686 = way0_hit ? record_wdata1_91 : _GEN_2533; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3687 = way0_hit ? record_wdata1_92 : _GEN_2534; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3688 = way0_hit ? record_wdata1_93 : _GEN_2535; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3689 = way0_hit ? record_wdata1_94 : _GEN_2536; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3690 = way0_hit ? record_wdata1_95 : _GEN_2537; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3691 = way0_hit ? record_wdata1_96 : _GEN_2538; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3692 = way0_hit ? record_wdata1_97 : _GEN_2539; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3693 = way0_hit ? record_wdata1_98 : _GEN_2540; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3694 = way0_hit ? record_wdata1_99 : _GEN_2541; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3695 = way0_hit ? record_wdata1_100 : _GEN_2542; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3696 = way0_hit ? record_wdata1_101 : _GEN_2543; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3697 = way0_hit ? record_wdata1_102 : _GEN_2544; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3698 = way0_hit ? record_wdata1_103 : _GEN_2545; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3699 = way0_hit ? record_wdata1_104 : _GEN_2546; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3700 = way0_hit ? record_wdata1_105 : _GEN_2547; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3701 = way0_hit ? record_wdata1_106 : _GEN_2548; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3702 = way0_hit ? record_wdata1_107 : _GEN_2549; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3703 = way0_hit ? record_wdata1_108 : _GEN_2550; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3704 = way0_hit ? record_wdata1_109 : _GEN_2551; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3705 = way0_hit ? record_wdata1_110 : _GEN_2552; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3706 = way0_hit ? record_wdata1_111 : _GEN_2553; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3707 = way0_hit ? record_wdata1_112 : _GEN_2554; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3708 = way0_hit ? record_wdata1_113 : _GEN_2555; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3709 = way0_hit ? record_wdata1_114 : _GEN_2556; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3710 = way0_hit ? record_wdata1_115 : _GEN_2557; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3711 = way0_hit ? record_wdata1_116 : _GEN_2558; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3712 = way0_hit ? record_wdata1_117 : _GEN_2559; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3713 = way0_hit ? record_wdata1_118 : _GEN_2560; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3714 = way0_hit ? record_wdata1_119 : _GEN_2561; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3715 = way0_hit ? record_wdata1_120 : _GEN_2562; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3716 = way0_hit ? record_wdata1_121 : _GEN_2563; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3717 = way0_hit ? record_wdata1_122 : _GEN_2564; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3718 = way0_hit ? record_wdata1_123 : _GEN_2565; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3719 = way0_hit ? record_wdata1_124 : _GEN_2566; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3720 = way0_hit ? record_wdata1_125 : _GEN_2567; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3721 = way0_hit ? record_wdata1_126 : _GEN_2568; // @[d_cache.scala 113:27 21:32]
  wire [63:0] _GEN_3722 = way0_hit ? record_wdata1_127 : _GEN_2569; // @[d_cache.scala 113:27 21:32]
  wire [7:0] _GEN_3723 = way0_hit ? record_wstrb1_0 : _GEN_2570; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3724 = way0_hit ? record_wstrb1_1 : _GEN_2571; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3725 = way0_hit ? record_wstrb1_2 : _GEN_2572; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3726 = way0_hit ? record_wstrb1_3 : _GEN_2573; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3727 = way0_hit ? record_wstrb1_4 : _GEN_2574; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3728 = way0_hit ? record_wstrb1_5 : _GEN_2575; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3729 = way0_hit ? record_wstrb1_6 : _GEN_2576; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3730 = way0_hit ? record_wstrb1_7 : _GEN_2577; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3731 = way0_hit ? record_wstrb1_8 : _GEN_2578; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3732 = way0_hit ? record_wstrb1_9 : _GEN_2579; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3733 = way0_hit ? record_wstrb1_10 : _GEN_2580; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3734 = way0_hit ? record_wstrb1_11 : _GEN_2581; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3735 = way0_hit ? record_wstrb1_12 : _GEN_2582; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3736 = way0_hit ? record_wstrb1_13 : _GEN_2583; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3737 = way0_hit ? record_wstrb1_14 : _GEN_2584; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3738 = way0_hit ? record_wstrb1_15 : _GEN_2585; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3739 = way0_hit ? record_wstrb1_16 : _GEN_2586; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3740 = way0_hit ? record_wstrb1_17 : _GEN_2587; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3741 = way0_hit ? record_wstrb1_18 : _GEN_2588; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3742 = way0_hit ? record_wstrb1_19 : _GEN_2589; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3743 = way0_hit ? record_wstrb1_20 : _GEN_2590; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3744 = way0_hit ? record_wstrb1_21 : _GEN_2591; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3745 = way0_hit ? record_wstrb1_22 : _GEN_2592; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3746 = way0_hit ? record_wstrb1_23 : _GEN_2593; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3747 = way0_hit ? record_wstrb1_24 : _GEN_2594; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3748 = way0_hit ? record_wstrb1_25 : _GEN_2595; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3749 = way0_hit ? record_wstrb1_26 : _GEN_2596; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3750 = way0_hit ? record_wstrb1_27 : _GEN_2597; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3751 = way0_hit ? record_wstrb1_28 : _GEN_2598; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3752 = way0_hit ? record_wstrb1_29 : _GEN_2599; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3753 = way0_hit ? record_wstrb1_30 : _GEN_2600; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3754 = way0_hit ? record_wstrb1_31 : _GEN_2601; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3755 = way0_hit ? record_wstrb1_32 : _GEN_2602; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3756 = way0_hit ? record_wstrb1_33 : _GEN_2603; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3757 = way0_hit ? record_wstrb1_34 : _GEN_2604; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3758 = way0_hit ? record_wstrb1_35 : _GEN_2605; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3759 = way0_hit ? record_wstrb1_36 : _GEN_2606; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3760 = way0_hit ? record_wstrb1_37 : _GEN_2607; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3761 = way0_hit ? record_wstrb1_38 : _GEN_2608; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3762 = way0_hit ? record_wstrb1_39 : _GEN_2609; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3763 = way0_hit ? record_wstrb1_40 : _GEN_2610; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3764 = way0_hit ? record_wstrb1_41 : _GEN_2611; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3765 = way0_hit ? record_wstrb1_42 : _GEN_2612; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3766 = way0_hit ? record_wstrb1_43 : _GEN_2613; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3767 = way0_hit ? record_wstrb1_44 : _GEN_2614; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3768 = way0_hit ? record_wstrb1_45 : _GEN_2615; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3769 = way0_hit ? record_wstrb1_46 : _GEN_2616; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3770 = way0_hit ? record_wstrb1_47 : _GEN_2617; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3771 = way0_hit ? record_wstrb1_48 : _GEN_2618; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3772 = way0_hit ? record_wstrb1_49 : _GEN_2619; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3773 = way0_hit ? record_wstrb1_50 : _GEN_2620; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3774 = way0_hit ? record_wstrb1_51 : _GEN_2621; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3775 = way0_hit ? record_wstrb1_52 : _GEN_2622; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3776 = way0_hit ? record_wstrb1_53 : _GEN_2623; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3777 = way0_hit ? record_wstrb1_54 : _GEN_2624; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3778 = way0_hit ? record_wstrb1_55 : _GEN_2625; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3779 = way0_hit ? record_wstrb1_56 : _GEN_2626; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3780 = way0_hit ? record_wstrb1_57 : _GEN_2627; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3781 = way0_hit ? record_wstrb1_58 : _GEN_2628; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3782 = way0_hit ? record_wstrb1_59 : _GEN_2629; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3783 = way0_hit ? record_wstrb1_60 : _GEN_2630; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3784 = way0_hit ? record_wstrb1_61 : _GEN_2631; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3785 = way0_hit ? record_wstrb1_62 : _GEN_2632; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3786 = way0_hit ? record_wstrb1_63 : _GEN_2633; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3787 = way0_hit ? record_wstrb1_64 : _GEN_2634; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3788 = way0_hit ? record_wstrb1_65 : _GEN_2635; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3789 = way0_hit ? record_wstrb1_66 : _GEN_2636; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3790 = way0_hit ? record_wstrb1_67 : _GEN_2637; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3791 = way0_hit ? record_wstrb1_68 : _GEN_2638; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3792 = way0_hit ? record_wstrb1_69 : _GEN_2639; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3793 = way0_hit ? record_wstrb1_70 : _GEN_2640; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3794 = way0_hit ? record_wstrb1_71 : _GEN_2641; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3795 = way0_hit ? record_wstrb1_72 : _GEN_2642; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3796 = way0_hit ? record_wstrb1_73 : _GEN_2643; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3797 = way0_hit ? record_wstrb1_74 : _GEN_2644; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3798 = way0_hit ? record_wstrb1_75 : _GEN_2645; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3799 = way0_hit ? record_wstrb1_76 : _GEN_2646; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3800 = way0_hit ? record_wstrb1_77 : _GEN_2647; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3801 = way0_hit ? record_wstrb1_78 : _GEN_2648; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3802 = way0_hit ? record_wstrb1_79 : _GEN_2649; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3803 = way0_hit ? record_wstrb1_80 : _GEN_2650; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3804 = way0_hit ? record_wstrb1_81 : _GEN_2651; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3805 = way0_hit ? record_wstrb1_82 : _GEN_2652; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3806 = way0_hit ? record_wstrb1_83 : _GEN_2653; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3807 = way0_hit ? record_wstrb1_84 : _GEN_2654; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3808 = way0_hit ? record_wstrb1_85 : _GEN_2655; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3809 = way0_hit ? record_wstrb1_86 : _GEN_2656; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3810 = way0_hit ? record_wstrb1_87 : _GEN_2657; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3811 = way0_hit ? record_wstrb1_88 : _GEN_2658; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3812 = way0_hit ? record_wstrb1_89 : _GEN_2659; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3813 = way0_hit ? record_wstrb1_90 : _GEN_2660; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3814 = way0_hit ? record_wstrb1_91 : _GEN_2661; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3815 = way0_hit ? record_wstrb1_92 : _GEN_2662; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3816 = way0_hit ? record_wstrb1_93 : _GEN_2663; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3817 = way0_hit ? record_wstrb1_94 : _GEN_2664; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3818 = way0_hit ? record_wstrb1_95 : _GEN_2665; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3819 = way0_hit ? record_wstrb1_96 : _GEN_2666; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3820 = way0_hit ? record_wstrb1_97 : _GEN_2667; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3821 = way0_hit ? record_wstrb1_98 : _GEN_2668; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3822 = way0_hit ? record_wstrb1_99 : _GEN_2669; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3823 = way0_hit ? record_wstrb1_100 : _GEN_2670; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3824 = way0_hit ? record_wstrb1_101 : _GEN_2671; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3825 = way0_hit ? record_wstrb1_102 : _GEN_2672; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3826 = way0_hit ? record_wstrb1_103 : _GEN_2673; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3827 = way0_hit ? record_wstrb1_104 : _GEN_2674; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3828 = way0_hit ? record_wstrb1_105 : _GEN_2675; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3829 = way0_hit ? record_wstrb1_106 : _GEN_2676; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3830 = way0_hit ? record_wstrb1_107 : _GEN_2677; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3831 = way0_hit ? record_wstrb1_108 : _GEN_2678; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3832 = way0_hit ? record_wstrb1_109 : _GEN_2679; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3833 = way0_hit ? record_wstrb1_110 : _GEN_2680; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3834 = way0_hit ? record_wstrb1_111 : _GEN_2681; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3835 = way0_hit ? record_wstrb1_112 : _GEN_2682; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3836 = way0_hit ? record_wstrb1_113 : _GEN_2683; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3837 = way0_hit ? record_wstrb1_114 : _GEN_2684; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3838 = way0_hit ? record_wstrb1_115 : _GEN_2685; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3839 = way0_hit ? record_wstrb1_116 : _GEN_2686; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3840 = way0_hit ? record_wstrb1_117 : _GEN_2687; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3841 = way0_hit ? record_wstrb1_118 : _GEN_2688; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3842 = way0_hit ? record_wstrb1_119 : _GEN_2689; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3843 = way0_hit ? record_wstrb1_120 : _GEN_2690; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3844 = way0_hit ? record_wstrb1_121 : _GEN_2691; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3845 = way0_hit ? record_wstrb1_122 : _GEN_2692; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3846 = way0_hit ? record_wstrb1_123 : _GEN_2693; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3847 = way0_hit ? record_wstrb1_124 : _GEN_2694; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3848 = way0_hit ? record_wstrb1_125 : _GEN_2695; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3849 = way0_hit ? record_wstrb1_126 : _GEN_2696; // @[d_cache.scala 113:27 22:32]
  wire [7:0] _GEN_3850 = way0_hit ? record_wstrb1_127 : _GEN_2697; // @[d_cache.scala 113:27 22:32]
  wire [63:0] _GEN_3851 = way0_hit ? record_pc_0 : _GEN_2698; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3852 = way0_hit ? record_pc_1 : _GEN_2699; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3853 = way0_hit ? record_pc_2 : _GEN_2700; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3854 = way0_hit ? record_pc_3 : _GEN_2701; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3855 = way0_hit ? record_pc_4 : _GEN_2702; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3856 = way0_hit ? record_pc_5 : _GEN_2703; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3857 = way0_hit ? record_pc_6 : _GEN_2704; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3858 = way0_hit ? record_pc_7 : _GEN_2705; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3859 = way0_hit ? record_pc_8 : _GEN_2706; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3860 = way0_hit ? record_pc_9 : _GEN_2707; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3861 = way0_hit ? record_pc_10 : _GEN_2708; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3862 = way0_hit ? record_pc_11 : _GEN_2709; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3863 = way0_hit ? record_pc_12 : _GEN_2710; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3864 = way0_hit ? record_pc_13 : _GEN_2711; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3865 = way0_hit ? record_pc_14 : _GEN_2712; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3866 = way0_hit ? record_pc_15 : _GEN_2713; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3867 = way0_hit ? record_pc_16 : _GEN_2714; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3868 = way0_hit ? record_pc_17 : _GEN_2715; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3869 = way0_hit ? record_pc_18 : _GEN_2716; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3870 = way0_hit ? record_pc_19 : _GEN_2717; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3871 = way0_hit ? record_pc_20 : _GEN_2718; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3872 = way0_hit ? record_pc_21 : _GEN_2719; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3873 = way0_hit ? record_pc_22 : _GEN_2720; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3874 = way0_hit ? record_pc_23 : _GEN_2721; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3875 = way0_hit ? record_pc_24 : _GEN_2722; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3876 = way0_hit ? record_pc_25 : _GEN_2723; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3877 = way0_hit ? record_pc_26 : _GEN_2724; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3878 = way0_hit ? record_pc_27 : _GEN_2725; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3879 = way0_hit ? record_pc_28 : _GEN_2726; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3880 = way0_hit ? record_pc_29 : _GEN_2727; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3881 = way0_hit ? record_pc_30 : _GEN_2728; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3882 = way0_hit ? record_pc_31 : _GEN_2729; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3883 = way0_hit ? record_pc_32 : _GEN_2730; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3884 = way0_hit ? record_pc_33 : _GEN_2731; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3885 = way0_hit ? record_pc_34 : _GEN_2732; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3886 = way0_hit ? record_pc_35 : _GEN_2733; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3887 = way0_hit ? record_pc_36 : _GEN_2734; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3888 = way0_hit ? record_pc_37 : _GEN_2735; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3889 = way0_hit ? record_pc_38 : _GEN_2736; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3890 = way0_hit ? record_pc_39 : _GEN_2737; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3891 = way0_hit ? record_pc_40 : _GEN_2738; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3892 = way0_hit ? record_pc_41 : _GEN_2739; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3893 = way0_hit ? record_pc_42 : _GEN_2740; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3894 = way0_hit ? record_pc_43 : _GEN_2741; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3895 = way0_hit ? record_pc_44 : _GEN_2742; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3896 = way0_hit ? record_pc_45 : _GEN_2743; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3897 = way0_hit ? record_pc_46 : _GEN_2744; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3898 = way0_hit ? record_pc_47 : _GEN_2745; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3899 = way0_hit ? record_pc_48 : _GEN_2746; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3900 = way0_hit ? record_pc_49 : _GEN_2747; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3901 = way0_hit ? record_pc_50 : _GEN_2748; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3902 = way0_hit ? record_pc_51 : _GEN_2749; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3903 = way0_hit ? record_pc_52 : _GEN_2750; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3904 = way0_hit ? record_pc_53 : _GEN_2751; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3905 = way0_hit ? record_pc_54 : _GEN_2752; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3906 = way0_hit ? record_pc_55 : _GEN_2753; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3907 = way0_hit ? record_pc_56 : _GEN_2754; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3908 = way0_hit ? record_pc_57 : _GEN_2755; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3909 = way0_hit ? record_pc_58 : _GEN_2756; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3910 = way0_hit ? record_pc_59 : _GEN_2757; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3911 = way0_hit ? record_pc_60 : _GEN_2758; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3912 = way0_hit ? record_pc_61 : _GEN_2759; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3913 = way0_hit ? record_pc_62 : _GEN_2760; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3914 = way0_hit ? record_pc_63 : _GEN_2761; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3915 = way0_hit ? record_pc_64 : _GEN_2762; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3916 = way0_hit ? record_pc_65 : _GEN_2763; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3917 = way0_hit ? record_pc_66 : _GEN_2764; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3918 = way0_hit ? record_pc_67 : _GEN_2765; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3919 = way0_hit ? record_pc_68 : _GEN_2766; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3920 = way0_hit ? record_pc_69 : _GEN_2767; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3921 = way0_hit ? record_pc_70 : _GEN_2768; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3922 = way0_hit ? record_pc_71 : _GEN_2769; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3923 = way0_hit ? record_pc_72 : _GEN_2770; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3924 = way0_hit ? record_pc_73 : _GEN_2771; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3925 = way0_hit ? record_pc_74 : _GEN_2772; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3926 = way0_hit ? record_pc_75 : _GEN_2773; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3927 = way0_hit ? record_pc_76 : _GEN_2774; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3928 = way0_hit ? record_pc_77 : _GEN_2775; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3929 = way0_hit ? record_pc_78 : _GEN_2776; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3930 = way0_hit ? record_pc_79 : _GEN_2777; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3931 = way0_hit ? record_pc_80 : _GEN_2778; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3932 = way0_hit ? record_pc_81 : _GEN_2779; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3933 = way0_hit ? record_pc_82 : _GEN_2780; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3934 = way0_hit ? record_pc_83 : _GEN_2781; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3935 = way0_hit ? record_pc_84 : _GEN_2782; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3936 = way0_hit ? record_pc_85 : _GEN_2783; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3937 = way0_hit ? record_pc_86 : _GEN_2784; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3938 = way0_hit ? record_pc_87 : _GEN_2785; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3939 = way0_hit ? record_pc_88 : _GEN_2786; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3940 = way0_hit ? record_pc_89 : _GEN_2787; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3941 = way0_hit ? record_pc_90 : _GEN_2788; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3942 = way0_hit ? record_pc_91 : _GEN_2789; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3943 = way0_hit ? record_pc_92 : _GEN_2790; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3944 = way0_hit ? record_pc_93 : _GEN_2791; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3945 = way0_hit ? record_pc_94 : _GEN_2792; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3946 = way0_hit ? record_pc_95 : _GEN_2793; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3947 = way0_hit ? record_pc_96 : _GEN_2794; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3948 = way0_hit ? record_pc_97 : _GEN_2795; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3949 = way0_hit ? record_pc_98 : _GEN_2796; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3950 = way0_hit ? record_pc_99 : _GEN_2797; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3951 = way0_hit ? record_pc_100 : _GEN_2798; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3952 = way0_hit ? record_pc_101 : _GEN_2799; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3953 = way0_hit ? record_pc_102 : _GEN_2800; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3954 = way0_hit ? record_pc_103 : _GEN_2801; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3955 = way0_hit ? record_pc_104 : _GEN_2802; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3956 = way0_hit ? record_pc_105 : _GEN_2803; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3957 = way0_hit ? record_pc_106 : _GEN_2804; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3958 = way0_hit ? record_pc_107 : _GEN_2805; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3959 = way0_hit ? record_pc_108 : _GEN_2806; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3960 = way0_hit ? record_pc_109 : _GEN_2807; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3961 = way0_hit ? record_pc_110 : _GEN_2808; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3962 = way0_hit ? record_pc_111 : _GEN_2809; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3963 = way0_hit ? record_pc_112 : _GEN_2810; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3964 = way0_hit ? record_pc_113 : _GEN_2811; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3965 = way0_hit ? record_pc_114 : _GEN_2812; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3966 = way0_hit ? record_pc_115 : _GEN_2813; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3967 = way0_hit ? record_pc_116 : _GEN_2814; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3968 = way0_hit ? record_pc_117 : _GEN_2815; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3969 = way0_hit ? record_pc_118 : _GEN_2816; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3970 = way0_hit ? record_pc_119 : _GEN_2817; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3971 = way0_hit ? record_pc_120 : _GEN_2818; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3972 = way0_hit ? record_pc_121 : _GEN_2819; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3973 = way0_hit ? record_pc_122 : _GEN_2820; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3974 = way0_hit ? record_pc_123 : _GEN_2821; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3975 = way0_hit ? record_pc_124 : _GEN_2822; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3976 = way0_hit ? record_pc_125 : _GEN_2823; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3977 = way0_hit ? record_pc_126 : _GEN_2824; // @[d_cache.scala 113:27 23:28]
  wire [63:0] _GEN_3978 = way0_hit ? record_pc_127 : _GEN_2825; // @[d_cache.scala 113:27 23:28]
  wire [31:0] _GEN_3979 = way0_hit ? record_addr_0 : _GEN_2826; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3980 = way0_hit ? record_addr_1 : _GEN_2827; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3981 = way0_hit ? record_addr_2 : _GEN_2828; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3982 = way0_hit ? record_addr_3 : _GEN_2829; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3983 = way0_hit ? record_addr_4 : _GEN_2830; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3984 = way0_hit ? record_addr_5 : _GEN_2831; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3985 = way0_hit ? record_addr_6 : _GEN_2832; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3986 = way0_hit ? record_addr_7 : _GEN_2833; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3987 = way0_hit ? record_addr_8 : _GEN_2834; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3988 = way0_hit ? record_addr_9 : _GEN_2835; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3989 = way0_hit ? record_addr_10 : _GEN_2836; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3990 = way0_hit ? record_addr_11 : _GEN_2837; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3991 = way0_hit ? record_addr_12 : _GEN_2838; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3992 = way0_hit ? record_addr_13 : _GEN_2839; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3993 = way0_hit ? record_addr_14 : _GEN_2840; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3994 = way0_hit ? record_addr_15 : _GEN_2841; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3995 = way0_hit ? record_addr_16 : _GEN_2842; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3996 = way0_hit ? record_addr_17 : _GEN_2843; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3997 = way0_hit ? record_addr_18 : _GEN_2844; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3998 = way0_hit ? record_addr_19 : _GEN_2845; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_3999 = way0_hit ? record_addr_20 : _GEN_2846; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4000 = way0_hit ? record_addr_21 : _GEN_2847; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4001 = way0_hit ? record_addr_22 : _GEN_2848; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4002 = way0_hit ? record_addr_23 : _GEN_2849; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4003 = way0_hit ? record_addr_24 : _GEN_2850; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4004 = way0_hit ? record_addr_25 : _GEN_2851; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4005 = way0_hit ? record_addr_26 : _GEN_2852; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4006 = way0_hit ? record_addr_27 : _GEN_2853; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4007 = way0_hit ? record_addr_28 : _GEN_2854; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4008 = way0_hit ? record_addr_29 : _GEN_2855; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4009 = way0_hit ? record_addr_30 : _GEN_2856; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4010 = way0_hit ? record_addr_31 : _GEN_2857; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4011 = way0_hit ? record_addr_32 : _GEN_2858; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4012 = way0_hit ? record_addr_33 : _GEN_2859; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4013 = way0_hit ? record_addr_34 : _GEN_2860; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4014 = way0_hit ? record_addr_35 : _GEN_2861; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4015 = way0_hit ? record_addr_36 : _GEN_2862; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4016 = way0_hit ? record_addr_37 : _GEN_2863; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4017 = way0_hit ? record_addr_38 : _GEN_2864; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4018 = way0_hit ? record_addr_39 : _GEN_2865; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4019 = way0_hit ? record_addr_40 : _GEN_2866; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4020 = way0_hit ? record_addr_41 : _GEN_2867; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4021 = way0_hit ? record_addr_42 : _GEN_2868; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4022 = way0_hit ? record_addr_43 : _GEN_2869; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4023 = way0_hit ? record_addr_44 : _GEN_2870; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4024 = way0_hit ? record_addr_45 : _GEN_2871; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4025 = way0_hit ? record_addr_46 : _GEN_2872; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4026 = way0_hit ? record_addr_47 : _GEN_2873; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4027 = way0_hit ? record_addr_48 : _GEN_2874; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4028 = way0_hit ? record_addr_49 : _GEN_2875; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4029 = way0_hit ? record_addr_50 : _GEN_2876; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4030 = way0_hit ? record_addr_51 : _GEN_2877; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4031 = way0_hit ? record_addr_52 : _GEN_2878; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4032 = way0_hit ? record_addr_53 : _GEN_2879; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4033 = way0_hit ? record_addr_54 : _GEN_2880; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4034 = way0_hit ? record_addr_55 : _GEN_2881; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4035 = way0_hit ? record_addr_56 : _GEN_2882; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4036 = way0_hit ? record_addr_57 : _GEN_2883; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4037 = way0_hit ? record_addr_58 : _GEN_2884; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4038 = way0_hit ? record_addr_59 : _GEN_2885; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4039 = way0_hit ? record_addr_60 : _GEN_2886; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4040 = way0_hit ? record_addr_61 : _GEN_2887; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4041 = way0_hit ? record_addr_62 : _GEN_2888; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4042 = way0_hit ? record_addr_63 : _GEN_2889; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4043 = way0_hit ? record_addr_64 : _GEN_2890; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4044 = way0_hit ? record_addr_65 : _GEN_2891; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4045 = way0_hit ? record_addr_66 : _GEN_2892; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4046 = way0_hit ? record_addr_67 : _GEN_2893; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4047 = way0_hit ? record_addr_68 : _GEN_2894; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4048 = way0_hit ? record_addr_69 : _GEN_2895; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4049 = way0_hit ? record_addr_70 : _GEN_2896; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4050 = way0_hit ? record_addr_71 : _GEN_2897; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4051 = way0_hit ? record_addr_72 : _GEN_2898; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4052 = way0_hit ? record_addr_73 : _GEN_2899; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4053 = way0_hit ? record_addr_74 : _GEN_2900; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4054 = way0_hit ? record_addr_75 : _GEN_2901; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4055 = way0_hit ? record_addr_76 : _GEN_2902; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4056 = way0_hit ? record_addr_77 : _GEN_2903; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4057 = way0_hit ? record_addr_78 : _GEN_2904; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4058 = way0_hit ? record_addr_79 : _GEN_2905; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4059 = way0_hit ? record_addr_80 : _GEN_2906; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4060 = way0_hit ? record_addr_81 : _GEN_2907; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4061 = way0_hit ? record_addr_82 : _GEN_2908; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4062 = way0_hit ? record_addr_83 : _GEN_2909; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4063 = way0_hit ? record_addr_84 : _GEN_2910; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4064 = way0_hit ? record_addr_85 : _GEN_2911; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4065 = way0_hit ? record_addr_86 : _GEN_2912; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4066 = way0_hit ? record_addr_87 : _GEN_2913; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4067 = way0_hit ? record_addr_88 : _GEN_2914; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4068 = way0_hit ? record_addr_89 : _GEN_2915; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4069 = way0_hit ? record_addr_90 : _GEN_2916; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4070 = way0_hit ? record_addr_91 : _GEN_2917; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4071 = way0_hit ? record_addr_92 : _GEN_2918; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4072 = way0_hit ? record_addr_93 : _GEN_2919; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4073 = way0_hit ? record_addr_94 : _GEN_2920; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4074 = way0_hit ? record_addr_95 : _GEN_2921; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4075 = way0_hit ? record_addr_96 : _GEN_2922; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4076 = way0_hit ? record_addr_97 : _GEN_2923; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4077 = way0_hit ? record_addr_98 : _GEN_2924; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4078 = way0_hit ? record_addr_99 : _GEN_2925; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4079 = way0_hit ? record_addr_100 : _GEN_2926; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4080 = way0_hit ? record_addr_101 : _GEN_2927; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4081 = way0_hit ? record_addr_102 : _GEN_2928; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4082 = way0_hit ? record_addr_103 : _GEN_2929; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4083 = way0_hit ? record_addr_104 : _GEN_2930; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4084 = way0_hit ? record_addr_105 : _GEN_2931; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4085 = way0_hit ? record_addr_106 : _GEN_2932; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4086 = way0_hit ? record_addr_107 : _GEN_2933; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4087 = way0_hit ? record_addr_108 : _GEN_2934; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4088 = way0_hit ? record_addr_109 : _GEN_2935; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4089 = way0_hit ? record_addr_110 : _GEN_2936; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4090 = way0_hit ? record_addr_111 : _GEN_2937; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4091 = way0_hit ? record_addr_112 : _GEN_2938; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4092 = way0_hit ? record_addr_113 : _GEN_2939; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4093 = way0_hit ? record_addr_114 : _GEN_2940; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4094 = way0_hit ? record_addr_115 : _GEN_2941; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4095 = way0_hit ? record_addr_116 : _GEN_2942; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4096 = way0_hit ? record_addr_117 : _GEN_2943; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4097 = way0_hit ? record_addr_118 : _GEN_2944; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4098 = way0_hit ? record_addr_119 : _GEN_2945; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4099 = way0_hit ? record_addr_120 : _GEN_2946; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4100 = way0_hit ? record_addr_121 : _GEN_2947; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4101 = way0_hit ? record_addr_122 : _GEN_2948; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4102 = way0_hit ? record_addr_123 : _GEN_2949; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4103 = way0_hit ? record_addr_124 : _GEN_2950; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4104 = way0_hit ? record_addr_125 : _GEN_2951; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4105 = way0_hit ? record_addr_126 : _GEN_2952; // @[d_cache.scala 113:27 24:30]
  wire [31:0] _GEN_4106 = way0_hit ? record_addr_127 : _GEN_2953; // @[d_cache.scala 113:27 24:30]
  wire  _GEN_4107 = way0_hit ? dirty_1_0 : _GEN_2954; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4108 = way0_hit ? dirty_1_1 : _GEN_2955; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4109 = way0_hit ? dirty_1_2 : _GEN_2956; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4110 = way0_hit ? dirty_1_3 : _GEN_2957; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4111 = way0_hit ? dirty_1_4 : _GEN_2958; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4112 = way0_hit ? dirty_1_5 : _GEN_2959; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4113 = way0_hit ? dirty_1_6 : _GEN_2960; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4114 = way0_hit ? dirty_1_7 : _GEN_2961; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4115 = way0_hit ? dirty_1_8 : _GEN_2962; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4116 = way0_hit ? dirty_1_9 : _GEN_2963; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4117 = way0_hit ? dirty_1_10 : _GEN_2964; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4118 = way0_hit ? dirty_1_11 : _GEN_2965; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4119 = way0_hit ? dirty_1_12 : _GEN_2966; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4120 = way0_hit ? dirty_1_13 : _GEN_2967; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4121 = way0_hit ? dirty_1_14 : _GEN_2968; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4122 = way0_hit ? dirty_1_15 : _GEN_2969; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4123 = way0_hit ? dirty_1_16 : _GEN_2970; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4124 = way0_hit ? dirty_1_17 : _GEN_2971; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4125 = way0_hit ? dirty_1_18 : _GEN_2972; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4126 = way0_hit ? dirty_1_19 : _GEN_2973; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4127 = way0_hit ? dirty_1_20 : _GEN_2974; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4128 = way0_hit ? dirty_1_21 : _GEN_2975; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4129 = way0_hit ? dirty_1_22 : _GEN_2976; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4130 = way0_hit ? dirty_1_23 : _GEN_2977; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4131 = way0_hit ? dirty_1_24 : _GEN_2978; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4132 = way0_hit ? dirty_1_25 : _GEN_2979; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4133 = way0_hit ? dirty_1_26 : _GEN_2980; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4134 = way0_hit ? dirty_1_27 : _GEN_2981; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4135 = way0_hit ? dirty_1_28 : _GEN_2982; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4136 = way0_hit ? dirty_1_29 : _GEN_2983; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4137 = way0_hit ? dirty_1_30 : _GEN_2984; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4138 = way0_hit ? dirty_1_31 : _GEN_2985; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4139 = way0_hit ? dirty_1_32 : _GEN_2986; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4140 = way0_hit ? dirty_1_33 : _GEN_2987; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4141 = way0_hit ? dirty_1_34 : _GEN_2988; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4142 = way0_hit ? dirty_1_35 : _GEN_2989; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4143 = way0_hit ? dirty_1_36 : _GEN_2990; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4144 = way0_hit ? dirty_1_37 : _GEN_2991; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4145 = way0_hit ? dirty_1_38 : _GEN_2992; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4146 = way0_hit ? dirty_1_39 : _GEN_2993; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4147 = way0_hit ? dirty_1_40 : _GEN_2994; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4148 = way0_hit ? dirty_1_41 : _GEN_2995; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4149 = way0_hit ? dirty_1_42 : _GEN_2996; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4150 = way0_hit ? dirty_1_43 : _GEN_2997; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4151 = way0_hit ? dirty_1_44 : _GEN_2998; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4152 = way0_hit ? dirty_1_45 : _GEN_2999; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4153 = way0_hit ? dirty_1_46 : _GEN_3000; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4154 = way0_hit ? dirty_1_47 : _GEN_3001; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4155 = way0_hit ? dirty_1_48 : _GEN_3002; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4156 = way0_hit ? dirty_1_49 : _GEN_3003; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4157 = way0_hit ? dirty_1_50 : _GEN_3004; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4158 = way0_hit ? dirty_1_51 : _GEN_3005; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4159 = way0_hit ? dirty_1_52 : _GEN_3006; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4160 = way0_hit ? dirty_1_53 : _GEN_3007; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4161 = way0_hit ? dirty_1_54 : _GEN_3008; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4162 = way0_hit ? dirty_1_55 : _GEN_3009; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4163 = way0_hit ? dirty_1_56 : _GEN_3010; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4164 = way0_hit ? dirty_1_57 : _GEN_3011; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4165 = way0_hit ? dirty_1_58 : _GEN_3012; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4166 = way0_hit ? dirty_1_59 : _GEN_3013; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4167 = way0_hit ? dirty_1_60 : _GEN_3014; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4168 = way0_hit ? dirty_1_61 : _GEN_3015; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4169 = way0_hit ? dirty_1_62 : _GEN_3016; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4170 = way0_hit ? dirty_1_63 : _GEN_3017; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4171 = way0_hit ? dirty_1_64 : _GEN_3018; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4172 = way0_hit ? dirty_1_65 : _GEN_3019; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4173 = way0_hit ? dirty_1_66 : _GEN_3020; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4174 = way0_hit ? dirty_1_67 : _GEN_3021; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4175 = way0_hit ? dirty_1_68 : _GEN_3022; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4176 = way0_hit ? dirty_1_69 : _GEN_3023; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4177 = way0_hit ? dirty_1_70 : _GEN_3024; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4178 = way0_hit ? dirty_1_71 : _GEN_3025; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4179 = way0_hit ? dirty_1_72 : _GEN_3026; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4180 = way0_hit ? dirty_1_73 : _GEN_3027; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4181 = way0_hit ? dirty_1_74 : _GEN_3028; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4182 = way0_hit ? dirty_1_75 : _GEN_3029; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4183 = way0_hit ? dirty_1_76 : _GEN_3030; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4184 = way0_hit ? dirty_1_77 : _GEN_3031; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4185 = way0_hit ? dirty_1_78 : _GEN_3032; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4186 = way0_hit ? dirty_1_79 : _GEN_3033; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4187 = way0_hit ? dirty_1_80 : _GEN_3034; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4188 = way0_hit ? dirty_1_81 : _GEN_3035; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4189 = way0_hit ? dirty_1_82 : _GEN_3036; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4190 = way0_hit ? dirty_1_83 : _GEN_3037; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4191 = way0_hit ? dirty_1_84 : _GEN_3038; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4192 = way0_hit ? dirty_1_85 : _GEN_3039; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4193 = way0_hit ? dirty_1_86 : _GEN_3040; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4194 = way0_hit ? dirty_1_87 : _GEN_3041; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4195 = way0_hit ? dirty_1_88 : _GEN_3042; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4196 = way0_hit ? dirty_1_89 : _GEN_3043; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4197 = way0_hit ? dirty_1_90 : _GEN_3044; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4198 = way0_hit ? dirty_1_91 : _GEN_3045; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4199 = way0_hit ? dirty_1_92 : _GEN_3046; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4200 = way0_hit ? dirty_1_93 : _GEN_3047; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4201 = way0_hit ? dirty_1_94 : _GEN_3048; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4202 = way0_hit ? dirty_1_95 : _GEN_3049; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4203 = way0_hit ? dirty_1_96 : _GEN_3050; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4204 = way0_hit ? dirty_1_97 : _GEN_3051; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4205 = way0_hit ? dirty_1_98 : _GEN_3052; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4206 = way0_hit ? dirty_1_99 : _GEN_3053; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4207 = way0_hit ? dirty_1_100 : _GEN_3054; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4208 = way0_hit ? dirty_1_101 : _GEN_3055; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4209 = way0_hit ? dirty_1_102 : _GEN_3056; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4210 = way0_hit ? dirty_1_103 : _GEN_3057; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4211 = way0_hit ? dirty_1_104 : _GEN_3058; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4212 = way0_hit ? dirty_1_105 : _GEN_3059; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4213 = way0_hit ? dirty_1_106 : _GEN_3060; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4214 = way0_hit ? dirty_1_107 : _GEN_3061; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4215 = way0_hit ? dirty_1_108 : _GEN_3062; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4216 = way0_hit ? dirty_1_109 : _GEN_3063; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4217 = way0_hit ? dirty_1_110 : _GEN_3064; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4218 = way0_hit ? dirty_1_111 : _GEN_3065; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4219 = way0_hit ? dirty_1_112 : _GEN_3066; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4220 = way0_hit ? dirty_1_113 : _GEN_3067; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4221 = way0_hit ? dirty_1_114 : _GEN_3068; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4222 = way0_hit ? dirty_1_115 : _GEN_3069; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4223 = way0_hit ? dirty_1_116 : _GEN_3070; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4224 = way0_hit ? dirty_1_117 : _GEN_3071; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4225 = way0_hit ? dirty_1_118 : _GEN_3072; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4226 = way0_hit ? dirty_1_119 : _GEN_3073; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4227 = way0_hit ? dirty_1_120 : _GEN_3074; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4228 = way0_hit ? dirty_1_121 : _GEN_3075; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4229 = way0_hit ? dirty_1_122 : _GEN_3076; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4230 = way0_hit ? dirty_1_123 : _GEN_3077; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4231 = way0_hit ? dirty_1_124 : _GEN_3078; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4232 = way0_hit ? dirty_1_125 : _GEN_3079; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4233 = way0_hit ? dirty_1_126 : _GEN_3080; // @[d_cache.scala 113:27 33:26]
  wire  _GEN_4234 = way0_hit ? dirty_1_127 : _GEN_3081; // @[d_cache.scala 113:27 33:26]
  wire [2:0] _GEN_4235 = io_from_axi_rvalid ? 3'h5 : state; // @[d_cache.scala 137:37 138:23 82:24]
  wire [63:0] _GEN_4236 = io_from_axi_rvalid ? io_from_axi_rdata : receive_data; // @[d_cache.scala 140:37 141:30 42:31]
  wire [2:0] _GEN_4237 = io_from_axi_bvalid ? 3'h0 : state; // @[d_cache.scala 145:37 146:23 82:24]
  wire [63:0] _GEN_4238 = 7'h0 == index ? receive_data : ram_0_0; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4239 = 7'h1 == index ? receive_data : ram_0_1; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4240 = 7'h2 == index ? receive_data : ram_0_2; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4241 = 7'h3 == index ? receive_data : ram_0_3; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4242 = 7'h4 == index ? receive_data : ram_0_4; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4243 = 7'h5 == index ? receive_data : ram_0_5; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4244 = 7'h6 == index ? receive_data : ram_0_6; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4245 = 7'h7 == index ? receive_data : ram_0_7; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4246 = 7'h8 == index ? receive_data : ram_0_8; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4247 = 7'h9 == index ? receive_data : ram_0_9; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4248 = 7'ha == index ? receive_data : ram_0_10; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4249 = 7'hb == index ? receive_data : ram_0_11; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4250 = 7'hc == index ? receive_data : ram_0_12; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4251 = 7'hd == index ? receive_data : ram_0_13; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4252 = 7'he == index ? receive_data : ram_0_14; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4253 = 7'hf == index ? receive_data : ram_0_15; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4254 = 7'h10 == index ? receive_data : ram_0_16; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4255 = 7'h11 == index ? receive_data : ram_0_17; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4256 = 7'h12 == index ? receive_data : ram_0_18; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4257 = 7'h13 == index ? receive_data : ram_0_19; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4258 = 7'h14 == index ? receive_data : ram_0_20; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4259 = 7'h15 == index ? receive_data : ram_0_21; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4260 = 7'h16 == index ? receive_data : ram_0_22; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4261 = 7'h17 == index ? receive_data : ram_0_23; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4262 = 7'h18 == index ? receive_data : ram_0_24; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4263 = 7'h19 == index ? receive_data : ram_0_25; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4264 = 7'h1a == index ? receive_data : ram_0_26; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4265 = 7'h1b == index ? receive_data : ram_0_27; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4266 = 7'h1c == index ? receive_data : ram_0_28; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4267 = 7'h1d == index ? receive_data : ram_0_29; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4268 = 7'h1e == index ? receive_data : ram_0_30; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4269 = 7'h1f == index ? receive_data : ram_0_31; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4270 = 7'h20 == index ? receive_data : ram_0_32; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4271 = 7'h21 == index ? receive_data : ram_0_33; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4272 = 7'h22 == index ? receive_data : ram_0_34; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4273 = 7'h23 == index ? receive_data : ram_0_35; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4274 = 7'h24 == index ? receive_data : ram_0_36; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4275 = 7'h25 == index ? receive_data : ram_0_37; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4276 = 7'h26 == index ? receive_data : ram_0_38; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4277 = 7'h27 == index ? receive_data : ram_0_39; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4278 = 7'h28 == index ? receive_data : ram_0_40; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4279 = 7'h29 == index ? receive_data : ram_0_41; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4280 = 7'h2a == index ? receive_data : ram_0_42; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4281 = 7'h2b == index ? receive_data : ram_0_43; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4282 = 7'h2c == index ? receive_data : ram_0_44; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4283 = 7'h2d == index ? receive_data : ram_0_45; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4284 = 7'h2e == index ? receive_data : ram_0_46; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4285 = 7'h2f == index ? receive_data : ram_0_47; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4286 = 7'h30 == index ? receive_data : ram_0_48; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4287 = 7'h31 == index ? receive_data : ram_0_49; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4288 = 7'h32 == index ? receive_data : ram_0_50; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4289 = 7'h33 == index ? receive_data : ram_0_51; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4290 = 7'h34 == index ? receive_data : ram_0_52; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4291 = 7'h35 == index ? receive_data : ram_0_53; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4292 = 7'h36 == index ? receive_data : ram_0_54; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4293 = 7'h37 == index ? receive_data : ram_0_55; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4294 = 7'h38 == index ? receive_data : ram_0_56; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4295 = 7'h39 == index ? receive_data : ram_0_57; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4296 = 7'h3a == index ? receive_data : ram_0_58; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4297 = 7'h3b == index ? receive_data : ram_0_59; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4298 = 7'h3c == index ? receive_data : ram_0_60; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4299 = 7'h3d == index ? receive_data : ram_0_61; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4300 = 7'h3e == index ? receive_data : ram_0_62; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4301 = 7'h3f == index ? receive_data : ram_0_63; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4302 = 7'h40 == index ? receive_data : ram_0_64; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4303 = 7'h41 == index ? receive_data : ram_0_65; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4304 = 7'h42 == index ? receive_data : ram_0_66; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4305 = 7'h43 == index ? receive_data : ram_0_67; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4306 = 7'h44 == index ? receive_data : ram_0_68; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4307 = 7'h45 == index ? receive_data : ram_0_69; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4308 = 7'h46 == index ? receive_data : ram_0_70; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4309 = 7'h47 == index ? receive_data : ram_0_71; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4310 = 7'h48 == index ? receive_data : ram_0_72; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4311 = 7'h49 == index ? receive_data : ram_0_73; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4312 = 7'h4a == index ? receive_data : ram_0_74; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4313 = 7'h4b == index ? receive_data : ram_0_75; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4314 = 7'h4c == index ? receive_data : ram_0_76; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4315 = 7'h4d == index ? receive_data : ram_0_77; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4316 = 7'h4e == index ? receive_data : ram_0_78; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4317 = 7'h4f == index ? receive_data : ram_0_79; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4318 = 7'h50 == index ? receive_data : ram_0_80; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4319 = 7'h51 == index ? receive_data : ram_0_81; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4320 = 7'h52 == index ? receive_data : ram_0_82; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4321 = 7'h53 == index ? receive_data : ram_0_83; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4322 = 7'h54 == index ? receive_data : ram_0_84; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4323 = 7'h55 == index ? receive_data : ram_0_85; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4324 = 7'h56 == index ? receive_data : ram_0_86; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4325 = 7'h57 == index ? receive_data : ram_0_87; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4326 = 7'h58 == index ? receive_data : ram_0_88; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4327 = 7'h59 == index ? receive_data : ram_0_89; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4328 = 7'h5a == index ? receive_data : ram_0_90; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4329 = 7'h5b == index ? receive_data : ram_0_91; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4330 = 7'h5c == index ? receive_data : ram_0_92; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4331 = 7'h5d == index ? receive_data : ram_0_93; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4332 = 7'h5e == index ? receive_data : ram_0_94; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4333 = 7'h5f == index ? receive_data : ram_0_95; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4334 = 7'h60 == index ? receive_data : ram_0_96; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4335 = 7'h61 == index ? receive_data : ram_0_97; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4336 = 7'h62 == index ? receive_data : ram_0_98; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4337 = 7'h63 == index ? receive_data : ram_0_99; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4338 = 7'h64 == index ? receive_data : ram_0_100; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4339 = 7'h65 == index ? receive_data : ram_0_101; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4340 = 7'h66 == index ? receive_data : ram_0_102; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4341 = 7'h67 == index ? receive_data : ram_0_103; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4342 = 7'h68 == index ? receive_data : ram_0_104; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4343 = 7'h69 == index ? receive_data : ram_0_105; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4344 = 7'h6a == index ? receive_data : ram_0_106; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4345 = 7'h6b == index ? receive_data : ram_0_107; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4346 = 7'h6c == index ? receive_data : ram_0_108; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4347 = 7'h6d == index ? receive_data : ram_0_109; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4348 = 7'h6e == index ? receive_data : ram_0_110; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4349 = 7'h6f == index ? receive_data : ram_0_111; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4350 = 7'h70 == index ? receive_data : ram_0_112; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4351 = 7'h71 == index ? receive_data : ram_0_113; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4352 = 7'h72 == index ? receive_data : ram_0_114; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4353 = 7'h73 == index ? receive_data : ram_0_115; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4354 = 7'h74 == index ? receive_data : ram_0_116; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4355 = 7'h75 == index ? receive_data : ram_0_117; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4356 = 7'h76 == index ? receive_data : ram_0_118; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4357 = 7'h77 == index ? receive_data : ram_0_119; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4358 = 7'h78 == index ? receive_data : ram_0_120; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4359 = 7'h79 == index ? receive_data : ram_0_121; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4360 = 7'h7a == index ? receive_data : ram_0_122; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4361 = 7'h7b == index ? receive_data : ram_0_123; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4362 = 7'h7c == index ? receive_data : ram_0_124; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4363 = 7'h7d == index ? receive_data : ram_0_125; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4364 = 7'h7e == index ? receive_data : ram_0_126; // @[d_cache.scala 152:{30,30} 19:24]
  wire [63:0] _GEN_4365 = 7'h7f == index ? receive_data : ram_0_127; // @[d_cache.scala 152:{30,30} 19:24]
  wire [31:0] _GEN_4366 = 7'h0 == index ? _GEN_19745 : tag_0_0; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4367 = 7'h1 == index ? _GEN_19745 : tag_0_1; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4368 = 7'h2 == index ? _GEN_19745 : tag_0_2; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4369 = 7'h3 == index ? _GEN_19745 : tag_0_3; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4370 = 7'h4 == index ? _GEN_19745 : tag_0_4; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4371 = 7'h5 == index ? _GEN_19745 : tag_0_5; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4372 = 7'h6 == index ? _GEN_19745 : tag_0_6; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4373 = 7'h7 == index ? _GEN_19745 : tag_0_7; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4374 = 7'h8 == index ? _GEN_19745 : tag_0_8; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4375 = 7'h9 == index ? _GEN_19745 : tag_0_9; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4376 = 7'ha == index ? _GEN_19745 : tag_0_10; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4377 = 7'hb == index ? _GEN_19745 : tag_0_11; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4378 = 7'hc == index ? _GEN_19745 : tag_0_12; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4379 = 7'hd == index ? _GEN_19745 : tag_0_13; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4380 = 7'he == index ? _GEN_19745 : tag_0_14; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4381 = 7'hf == index ? _GEN_19745 : tag_0_15; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4382 = 7'h10 == index ? _GEN_19745 : tag_0_16; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4383 = 7'h11 == index ? _GEN_19745 : tag_0_17; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4384 = 7'h12 == index ? _GEN_19745 : tag_0_18; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4385 = 7'h13 == index ? _GEN_19745 : tag_0_19; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4386 = 7'h14 == index ? _GEN_19745 : tag_0_20; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4387 = 7'h15 == index ? _GEN_19745 : tag_0_21; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4388 = 7'h16 == index ? _GEN_19745 : tag_0_22; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4389 = 7'h17 == index ? _GEN_19745 : tag_0_23; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4390 = 7'h18 == index ? _GEN_19745 : tag_0_24; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4391 = 7'h19 == index ? _GEN_19745 : tag_0_25; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4392 = 7'h1a == index ? _GEN_19745 : tag_0_26; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4393 = 7'h1b == index ? _GEN_19745 : tag_0_27; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4394 = 7'h1c == index ? _GEN_19745 : tag_0_28; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4395 = 7'h1d == index ? _GEN_19745 : tag_0_29; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4396 = 7'h1e == index ? _GEN_19745 : tag_0_30; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4397 = 7'h1f == index ? _GEN_19745 : tag_0_31; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4398 = 7'h20 == index ? _GEN_19745 : tag_0_32; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4399 = 7'h21 == index ? _GEN_19745 : tag_0_33; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4400 = 7'h22 == index ? _GEN_19745 : tag_0_34; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4401 = 7'h23 == index ? _GEN_19745 : tag_0_35; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4402 = 7'h24 == index ? _GEN_19745 : tag_0_36; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4403 = 7'h25 == index ? _GEN_19745 : tag_0_37; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4404 = 7'h26 == index ? _GEN_19745 : tag_0_38; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4405 = 7'h27 == index ? _GEN_19745 : tag_0_39; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4406 = 7'h28 == index ? _GEN_19745 : tag_0_40; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4407 = 7'h29 == index ? _GEN_19745 : tag_0_41; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4408 = 7'h2a == index ? _GEN_19745 : tag_0_42; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4409 = 7'h2b == index ? _GEN_19745 : tag_0_43; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4410 = 7'h2c == index ? _GEN_19745 : tag_0_44; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4411 = 7'h2d == index ? _GEN_19745 : tag_0_45; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4412 = 7'h2e == index ? _GEN_19745 : tag_0_46; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4413 = 7'h2f == index ? _GEN_19745 : tag_0_47; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4414 = 7'h30 == index ? _GEN_19745 : tag_0_48; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4415 = 7'h31 == index ? _GEN_19745 : tag_0_49; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4416 = 7'h32 == index ? _GEN_19745 : tag_0_50; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4417 = 7'h33 == index ? _GEN_19745 : tag_0_51; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4418 = 7'h34 == index ? _GEN_19745 : tag_0_52; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4419 = 7'h35 == index ? _GEN_19745 : tag_0_53; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4420 = 7'h36 == index ? _GEN_19745 : tag_0_54; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4421 = 7'h37 == index ? _GEN_19745 : tag_0_55; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4422 = 7'h38 == index ? _GEN_19745 : tag_0_56; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4423 = 7'h39 == index ? _GEN_19745 : tag_0_57; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4424 = 7'h3a == index ? _GEN_19745 : tag_0_58; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4425 = 7'h3b == index ? _GEN_19745 : tag_0_59; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4426 = 7'h3c == index ? _GEN_19745 : tag_0_60; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4427 = 7'h3d == index ? _GEN_19745 : tag_0_61; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4428 = 7'h3e == index ? _GEN_19745 : tag_0_62; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4429 = 7'h3f == index ? _GEN_19745 : tag_0_63; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4430 = 7'h40 == index ? _GEN_19745 : tag_0_64; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4431 = 7'h41 == index ? _GEN_19745 : tag_0_65; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4432 = 7'h42 == index ? _GEN_19745 : tag_0_66; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4433 = 7'h43 == index ? _GEN_19745 : tag_0_67; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4434 = 7'h44 == index ? _GEN_19745 : tag_0_68; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4435 = 7'h45 == index ? _GEN_19745 : tag_0_69; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4436 = 7'h46 == index ? _GEN_19745 : tag_0_70; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4437 = 7'h47 == index ? _GEN_19745 : tag_0_71; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4438 = 7'h48 == index ? _GEN_19745 : tag_0_72; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4439 = 7'h49 == index ? _GEN_19745 : tag_0_73; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4440 = 7'h4a == index ? _GEN_19745 : tag_0_74; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4441 = 7'h4b == index ? _GEN_19745 : tag_0_75; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4442 = 7'h4c == index ? _GEN_19745 : tag_0_76; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4443 = 7'h4d == index ? _GEN_19745 : tag_0_77; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4444 = 7'h4e == index ? _GEN_19745 : tag_0_78; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4445 = 7'h4f == index ? _GEN_19745 : tag_0_79; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4446 = 7'h50 == index ? _GEN_19745 : tag_0_80; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4447 = 7'h51 == index ? _GEN_19745 : tag_0_81; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4448 = 7'h52 == index ? _GEN_19745 : tag_0_82; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4449 = 7'h53 == index ? _GEN_19745 : tag_0_83; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4450 = 7'h54 == index ? _GEN_19745 : tag_0_84; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4451 = 7'h55 == index ? _GEN_19745 : tag_0_85; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4452 = 7'h56 == index ? _GEN_19745 : tag_0_86; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4453 = 7'h57 == index ? _GEN_19745 : tag_0_87; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4454 = 7'h58 == index ? _GEN_19745 : tag_0_88; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4455 = 7'h59 == index ? _GEN_19745 : tag_0_89; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4456 = 7'h5a == index ? _GEN_19745 : tag_0_90; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4457 = 7'h5b == index ? _GEN_19745 : tag_0_91; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4458 = 7'h5c == index ? _GEN_19745 : tag_0_92; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4459 = 7'h5d == index ? _GEN_19745 : tag_0_93; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4460 = 7'h5e == index ? _GEN_19745 : tag_0_94; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4461 = 7'h5f == index ? _GEN_19745 : tag_0_95; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4462 = 7'h60 == index ? _GEN_19745 : tag_0_96; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4463 = 7'h61 == index ? _GEN_19745 : tag_0_97; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4464 = 7'h62 == index ? _GEN_19745 : tag_0_98; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4465 = 7'h63 == index ? _GEN_19745 : tag_0_99; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4466 = 7'h64 == index ? _GEN_19745 : tag_0_100; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4467 = 7'h65 == index ? _GEN_19745 : tag_0_101; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4468 = 7'h66 == index ? _GEN_19745 : tag_0_102; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4469 = 7'h67 == index ? _GEN_19745 : tag_0_103; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4470 = 7'h68 == index ? _GEN_19745 : tag_0_104; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4471 = 7'h69 == index ? _GEN_19745 : tag_0_105; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4472 = 7'h6a == index ? _GEN_19745 : tag_0_106; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4473 = 7'h6b == index ? _GEN_19745 : tag_0_107; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4474 = 7'h6c == index ? _GEN_19745 : tag_0_108; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4475 = 7'h6d == index ? _GEN_19745 : tag_0_109; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4476 = 7'h6e == index ? _GEN_19745 : tag_0_110; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4477 = 7'h6f == index ? _GEN_19745 : tag_0_111; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4478 = 7'h70 == index ? _GEN_19745 : tag_0_112; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4479 = 7'h71 == index ? _GEN_19745 : tag_0_113; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4480 = 7'h72 == index ? _GEN_19745 : tag_0_114; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4481 = 7'h73 == index ? _GEN_19745 : tag_0_115; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4482 = 7'h74 == index ? _GEN_19745 : tag_0_116; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4483 = 7'h75 == index ? _GEN_19745 : tag_0_117; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4484 = 7'h76 == index ? _GEN_19745 : tag_0_118; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4485 = 7'h77 == index ? _GEN_19745 : tag_0_119; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4486 = 7'h78 == index ? _GEN_19745 : tag_0_120; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4487 = 7'h79 == index ? _GEN_19745 : tag_0_121; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4488 = 7'h7a == index ? _GEN_19745 : tag_0_122; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4489 = 7'h7b == index ? _GEN_19745 : tag_0_123; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4490 = 7'h7c == index ? _GEN_19745 : tag_0_124; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4491 = 7'h7d == index ? _GEN_19745 : tag_0_125; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4492 = 7'h7e == index ? _GEN_19745 : tag_0_126; // @[d_cache.scala 153:{30,30} 28:24]
  wire [31:0] _GEN_4493 = 7'h7f == index ? _GEN_19745 : tag_0_127; // @[d_cache.scala 153:{30,30} 28:24]
  wire  _GEN_4494 = _GEN_19748 | valid_0_0; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4495 = _GEN_19749 | valid_0_1; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4496 = _GEN_19750 | valid_0_2; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4497 = _GEN_19751 | valid_0_3; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4498 = _GEN_19752 | valid_0_4; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4499 = _GEN_19753 | valid_0_5; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4500 = _GEN_19754 | valid_0_6; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4501 = _GEN_19755 | valid_0_7; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4502 = _GEN_19756 | valid_0_8; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4503 = _GEN_19757 | valid_0_9; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4504 = _GEN_19758 | valid_0_10; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4505 = _GEN_19759 | valid_0_11; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4506 = _GEN_19760 | valid_0_12; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4507 = _GEN_19761 | valid_0_13; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4508 = _GEN_19762 | valid_0_14; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4509 = _GEN_19763 | valid_0_15; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4510 = _GEN_19764 | valid_0_16; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4511 = _GEN_19765 | valid_0_17; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4512 = _GEN_19766 | valid_0_18; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4513 = _GEN_19767 | valid_0_19; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4514 = _GEN_19768 | valid_0_20; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4515 = _GEN_19769 | valid_0_21; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4516 = _GEN_19770 | valid_0_22; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4517 = _GEN_19771 | valid_0_23; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4518 = _GEN_19772 | valid_0_24; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4519 = _GEN_19773 | valid_0_25; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4520 = _GEN_19774 | valid_0_26; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4521 = _GEN_19775 | valid_0_27; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4522 = _GEN_19776 | valid_0_28; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4523 = _GEN_19777 | valid_0_29; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4524 = _GEN_19778 | valid_0_30; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4525 = _GEN_19779 | valid_0_31; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4526 = _GEN_19780 | valid_0_32; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4527 = _GEN_19781 | valid_0_33; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4528 = _GEN_19782 | valid_0_34; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4529 = _GEN_19783 | valid_0_35; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4530 = _GEN_19784 | valid_0_36; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4531 = _GEN_19785 | valid_0_37; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4532 = _GEN_19786 | valid_0_38; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4533 = _GEN_19787 | valid_0_39; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4534 = _GEN_19788 | valid_0_40; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4535 = _GEN_19789 | valid_0_41; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4536 = _GEN_19790 | valid_0_42; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4537 = _GEN_19791 | valid_0_43; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4538 = _GEN_19792 | valid_0_44; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4539 = _GEN_19793 | valid_0_45; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4540 = _GEN_19794 | valid_0_46; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4541 = _GEN_19795 | valid_0_47; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4542 = _GEN_19796 | valid_0_48; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4543 = _GEN_19797 | valid_0_49; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4544 = _GEN_19798 | valid_0_50; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4545 = _GEN_19799 | valid_0_51; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4546 = _GEN_19800 | valid_0_52; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4547 = _GEN_19801 | valid_0_53; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4548 = _GEN_19802 | valid_0_54; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4549 = _GEN_19803 | valid_0_55; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4550 = _GEN_19804 | valid_0_56; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4551 = _GEN_19805 | valid_0_57; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4552 = _GEN_19806 | valid_0_58; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4553 = _GEN_19807 | valid_0_59; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4554 = _GEN_19808 | valid_0_60; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4555 = _GEN_19809 | valid_0_61; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4556 = _GEN_19810 | valid_0_62; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4557 = _GEN_19811 | valid_0_63; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4558 = _GEN_19812 | valid_0_64; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4559 = _GEN_19813 | valid_0_65; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4560 = _GEN_19814 | valid_0_66; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4561 = _GEN_19815 | valid_0_67; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4562 = _GEN_19816 | valid_0_68; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4563 = _GEN_19817 | valid_0_69; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4564 = _GEN_19818 | valid_0_70; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4565 = _GEN_19819 | valid_0_71; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4566 = _GEN_19820 | valid_0_72; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4567 = _GEN_19821 | valid_0_73; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4568 = _GEN_19822 | valid_0_74; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4569 = _GEN_19823 | valid_0_75; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4570 = _GEN_19824 | valid_0_76; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4571 = _GEN_19825 | valid_0_77; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4572 = _GEN_19826 | valid_0_78; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4573 = _GEN_19827 | valid_0_79; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4574 = _GEN_19828 | valid_0_80; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4575 = _GEN_19829 | valid_0_81; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4576 = _GEN_19830 | valid_0_82; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4577 = _GEN_19831 | valid_0_83; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4578 = _GEN_19832 | valid_0_84; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4579 = _GEN_19833 | valid_0_85; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4580 = _GEN_19834 | valid_0_86; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4581 = _GEN_19835 | valid_0_87; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4582 = _GEN_19836 | valid_0_88; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4583 = _GEN_19837 | valid_0_89; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4584 = _GEN_19838 | valid_0_90; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4585 = _GEN_19839 | valid_0_91; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4586 = _GEN_19840 | valid_0_92; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4587 = _GEN_19841 | valid_0_93; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4588 = _GEN_19842 | valid_0_94; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4589 = _GEN_19843 | valid_0_95; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4590 = _GEN_19844 | valid_0_96; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4591 = _GEN_19845 | valid_0_97; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4592 = _GEN_19846 | valid_0_98; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4593 = _GEN_19847 | valid_0_99; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4594 = _GEN_19848 | valid_0_100; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4595 = _GEN_19849 | valid_0_101; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4596 = _GEN_19850 | valid_0_102; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4597 = _GEN_19851 | valid_0_103; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4598 = _GEN_19852 | valid_0_104; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4599 = _GEN_19853 | valid_0_105; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4600 = _GEN_19854 | valid_0_106; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4601 = _GEN_19855 | valid_0_107; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4602 = _GEN_19856 | valid_0_108; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4603 = _GEN_19857 | valid_0_109; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4604 = _GEN_19858 | valid_0_110; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4605 = _GEN_19859 | valid_0_111; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4606 = _GEN_19860 | valid_0_112; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4607 = _GEN_19861 | valid_0_113; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4608 = _GEN_19862 | valid_0_114; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4609 = _GEN_19863 | valid_0_115; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4610 = _GEN_19864 | valid_0_116; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4611 = _GEN_19865 | valid_0_117; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4612 = _GEN_19866 | valid_0_118; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4613 = _GEN_19867 | valid_0_119; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4614 = _GEN_19868 | valid_0_120; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4615 = _GEN_19869 | valid_0_121; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4616 = _GEN_19870 | valid_0_122; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4617 = _GEN_19871 | valid_0_123; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4618 = _GEN_19872 | valid_0_124; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4619 = _GEN_19873 | valid_0_125; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4620 = _GEN_19874 | valid_0_126; // @[d_cache.scala 154:{32,32} 30:26]
  wire  _GEN_4621 = _GEN_19875 | valid_0_127; // @[d_cache.scala 154:{32,32} 30:26]
  wire [63:0] _GEN_4622 = 7'h0 == index ? receive_data : ram_1_0; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4623 = 7'h1 == index ? receive_data : ram_1_1; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4624 = 7'h2 == index ? receive_data : ram_1_2; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4625 = 7'h3 == index ? receive_data : ram_1_3; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4626 = 7'h4 == index ? receive_data : ram_1_4; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4627 = 7'h5 == index ? receive_data : ram_1_5; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4628 = 7'h6 == index ? receive_data : ram_1_6; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4629 = 7'h7 == index ? receive_data : ram_1_7; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4630 = 7'h8 == index ? receive_data : ram_1_8; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4631 = 7'h9 == index ? receive_data : ram_1_9; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4632 = 7'ha == index ? receive_data : ram_1_10; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4633 = 7'hb == index ? receive_data : ram_1_11; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4634 = 7'hc == index ? receive_data : ram_1_12; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4635 = 7'hd == index ? receive_data : ram_1_13; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4636 = 7'he == index ? receive_data : ram_1_14; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4637 = 7'hf == index ? receive_data : ram_1_15; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4638 = 7'h10 == index ? receive_data : ram_1_16; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4639 = 7'h11 == index ? receive_data : ram_1_17; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4640 = 7'h12 == index ? receive_data : ram_1_18; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4641 = 7'h13 == index ? receive_data : ram_1_19; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4642 = 7'h14 == index ? receive_data : ram_1_20; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4643 = 7'h15 == index ? receive_data : ram_1_21; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4644 = 7'h16 == index ? receive_data : ram_1_22; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4645 = 7'h17 == index ? receive_data : ram_1_23; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4646 = 7'h18 == index ? receive_data : ram_1_24; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4647 = 7'h19 == index ? receive_data : ram_1_25; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4648 = 7'h1a == index ? receive_data : ram_1_26; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4649 = 7'h1b == index ? receive_data : ram_1_27; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4650 = 7'h1c == index ? receive_data : ram_1_28; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4651 = 7'h1d == index ? receive_data : ram_1_29; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4652 = 7'h1e == index ? receive_data : ram_1_30; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4653 = 7'h1f == index ? receive_data : ram_1_31; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4654 = 7'h20 == index ? receive_data : ram_1_32; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4655 = 7'h21 == index ? receive_data : ram_1_33; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4656 = 7'h22 == index ? receive_data : ram_1_34; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4657 = 7'h23 == index ? receive_data : ram_1_35; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4658 = 7'h24 == index ? receive_data : ram_1_36; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4659 = 7'h25 == index ? receive_data : ram_1_37; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4660 = 7'h26 == index ? receive_data : ram_1_38; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4661 = 7'h27 == index ? receive_data : ram_1_39; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4662 = 7'h28 == index ? receive_data : ram_1_40; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4663 = 7'h29 == index ? receive_data : ram_1_41; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4664 = 7'h2a == index ? receive_data : ram_1_42; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4665 = 7'h2b == index ? receive_data : ram_1_43; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4666 = 7'h2c == index ? receive_data : ram_1_44; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4667 = 7'h2d == index ? receive_data : ram_1_45; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4668 = 7'h2e == index ? receive_data : ram_1_46; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4669 = 7'h2f == index ? receive_data : ram_1_47; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4670 = 7'h30 == index ? receive_data : ram_1_48; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4671 = 7'h31 == index ? receive_data : ram_1_49; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4672 = 7'h32 == index ? receive_data : ram_1_50; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4673 = 7'h33 == index ? receive_data : ram_1_51; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4674 = 7'h34 == index ? receive_data : ram_1_52; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4675 = 7'h35 == index ? receive_data : ram_1_53; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4676 = 7'h36 == index ? receive_data : ram_1_54; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4677 = 7'h37 == index ? receive_data : ram_1_55; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4678 = 7'h38 == index ? receive_data : ram_1_56; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4679 = 7'h39 == index ? receive_data : ram_1_57; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4680 = 7'h3a == index ? receive_data : ram_1_58; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4681 = 7'h3b == index ? receive_data : ram_1_59; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4682 = 7'h3c == index ? receive_data : ram_1_60; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4683 = 7'h3d == index ? receive_data : ram_1_61; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4684 = 7'h3e == index ? receive_data : ram_1_62; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4685 = 7'h3f == index ? receive_data : ram_1_63; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4686 = 7'h40 == index ? receive_data : ram_1_64; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4687 = 7'h41 == index ? receive_data : ram_1_65; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4688 = 7'h42 == index ? receive_data : ram_1_66; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4689 = 7'h43 == index ? receive_data : ram_1_67; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4690 = 7'h44 == index ? receive_data : ram_1_68; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4691 = 7'h45 == index ? receive_data : ram_1_69; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4692 = 7'h46 == index ? receive_data : ram_1_70; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4693 = 7'h47 == index ? receive_data : ram_1_71; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4694 = 7'h48 == index ? receive_data : ram_1_72; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4695 = 7'h49 == index ? receive_data : ram_1_73; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4696 = 7'h4a == index ? receive_data : ram_1_74; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4697 = 7'h4b == index ? receive_data : ram_1_75; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4698 = 7'h4c == index ? receive_data : ram_1_76; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4699 = 7'h4d == index ? receive_data : ram_1_77; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4700 = 7'h4e == index ? receive_data : ram_1_78; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4701 = 7'h4f == index ? receive_data : ram_1_79; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4702 = 7'h50 == index ? receive_data : ram_1_80; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4703 = 7'h51 == index ? receive_data : ram_1_81; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4704 = 7'h52 == index ? receive_data : ram_1_82; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4705 = 7'h53 == index ? receive_data : ram_1_83; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4706 = 7'h54 == index ? receive_data : ram_1_84; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4707 = 7'h55 == index ? receive_data : ram_1_85; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4708 = 7'h56 == index ? receive_data : ram_1_86; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4709 = 7'h57 == index ? receive_data : ram_1_87; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4710 = 7'h58 == index ? receive_data : ram_1_88; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4711 = 7'h59 == index ? receive_data : ram_1_89; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4712 = 7'h5a == index ? receive_data : ram_1_90; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4713 = 7'h5b == index ? receive_data : ram_1_91; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4714 = 7'h5c == index ? receive_data : ram_1_92; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4715 = 7'h5d == index ? receive_data : ram_1_93; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4716 = 7'h5e == index ? receive_data : ram_1_94; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4717 = 7'h5f == index ? receive_data : ram_1_95; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4718 = 7'h60 == index ? receive_data : ram_1_96; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4719 = 7'h61 == index ? receive_data : ram_1_97; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4720 = 7'h62 == index ? receive_data : ram_1_98; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4721 = 7'h63 == index ? receive_data : ram_1_99; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4722 = 7'h64 == index ? receive_data : ram_1_100; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4723 = 7'h65 == index ? receive_data : ram_1_101; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4724 = 7'h66 == index ? receive_data : ram_1_102; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4725 = 7'h67 == index ? receive_data : ram_1_103; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4726 = 7'h68 == index ? receive_data : ram_1_104; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4727 = 7'h69 == index ? receive_data : ram_1_105; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4728 = 7'h6a == index ? receive_data : ram_1_106; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4729 = 7'h6b == index ? receive_data : ram_1_107; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4730 = 7'h6c == index ? receive_data : ram_1_108; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4731 = 7'h6d == index ? receive_data : ram_1_109; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4732 = 7'h6e == index ? receive_data : ram_1_110; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4733 = 7'h6f == index ? receive_data : ram_1_111; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4734 = 7'h70 == index ? receive_data : ram_1_112; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4735 = 7'h71 == index ? receive_data : ram_1_113; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4736 = 7'h72 == index ? receive_data : ram_1_114; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4737 = 7'h73 == index ? receive_data : ram_1_115; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4738 = 7'h74 == index ? receive_data : ram_1_116; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4739 = 7'h75 == index ? receive_data : ram_1_117; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4740 = 7'h76 == index ? receive_data : ram_1_118; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4741 = 7'h77 == index ? receive_data : ram_1_119; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4742 = 7'h78 == index ? receive_data : ram_1_120; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4743 = 7'h79 == index ? receive_data : ram_1_121; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4744 = 7'h7a == index ? receive_data : ram_1_122; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4745 = 7'h7b == index ? receive_data : ram_1_123; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4746 = 7'h7c == index ? receive_data : ram_1_124; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4747 = 7'h7d == index ? receive_data : ram_1_125; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4748 = 7'h7e == index ? receive_data : ram_1_126; // @[d_cache.scala 158:{30,30} 20:24]
  wire [63:0] _GEN_4749 = 7'h7f == index ? receive_data : ram_1_127; // @[d_cache.scala 158:{30,30} 20:24]
  wire [31:0] _GEN_4750 = 7'h0 == index ? _GEN_19745 : tag_1_0; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4751 = 7'h1 == index ? _GEN_19745 : tag_1_1; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4752 = 7'h2 == index ? _GEN_19745 : tag_1_2; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4753 = 7'h3 == index ? _GEN_19745 : tag_1_3; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4754 = 7'h4 == index ? _GEN_19745 : tag_1_4; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4755 = 7'h5 == index ? _GEN_19745 : tag_1_5; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4756 = 7'h6 == index ? _GEN_19745 : tag_1_6; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4757 = 7'h7 == index ? _GEN_19745 : tag_1_7; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4758 = 7'h8 == index ? _GEN_19745 : tag_1_8; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4759 = 7'h9 == index ? _GEN_19745 : tag_1_9; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4760 = 7'ha == index ? _GEN_19745 : tag_1_10; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4761 = 7'hb == index ? _GEN_19745 : tag_1_11; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4762 = 7'hc == index ? _GEN_19745 : tag_1_12; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4763 = 7'hd == index ? _GEN_19745 : tag_1_13; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4764 = 7'he == index ? _GEN_19745 : tag_1_14; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4765 = 7'hf == index ? _GEN_19745 : tag_1_15; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4766 = 7'h10 == index ? _GEN_19745 : tag_1_16; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4767 = 7'h11 == index ? _GEN_19745 : tag_1_17; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4768 = 7'h12 == index ? _GEN_19745 : tag_1_18; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4769 = 7'h13 == index ? _GEN_19745 : tag_1_19; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4770 = 7'h14 == index ? _GEN_19745 : tag_1_20; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4771 = 7'h15 == index ? _GEN_19745 : tag_1_21; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4772 = 7'h16 == index ? _GEN_19745 : tag_1_22; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4773 = 7'h17 == index ? _GEN_19745 : tag_1_23; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4774 = 7'h18 == index ? _GEN_19745 : tag_1_24; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4775 = 7'h19 == index ? _GEN_19745 : tag_1_25; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4776 = 7'h1a == index ? _GEN_19745 : tag_1_26; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4777 = 7'h1b == index ? _GEN_19745 : tag_1_27; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4778 = 7'h1c == index ? _GEN_19745 : tag_1_28; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4779 = 7'h1d == index ? _GEN_19745 : tag_1_29; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4780 = 7'h1e == index ? _GEN_19745 : tag_1_30; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4781 = 7'h1f == index ? _GEN_19745 : tag_1_31; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4782 = 7'h20 == index ? _GEN_19745 : tag_1_32; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4783 = 7'h21 == index ? _GEN_19745 : tag_1_33; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4784 = 7'h22 == index ? _GEN_19745 : tag_1_34; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4785 = 7'h23 == index ? _GEN_19745 : tag_1_35; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4786 = 7'h24 == index ? _GEN_19745 : tag_1_36; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4787 = 7'h25 == index ? _GEN_19745 : tag_1_37; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4788 = 7'h26 == index ? _GEN_19745 : tag_1_38; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4789 = 7'h27 == index ? _GEN_19745 : tag_1_39; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4790 = 7'h28 == index ? _GEN_19745 : tag_1_40; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4791 = 7'h29 == index ? _GEN_19745 : tag_1_41; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4792 = 7'h2a == index ? _GEN_19745 : tag_1_42; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4793 = 7'h2b == index ? _GEN_19745 : tag_1_43; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4794 = 7'h2c == index ? _GEN_19745 : tag_1_44; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4795 = 7'h2d == index ? _GEN_19745 : tag_1_45; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4796 = 7'h2e == index ? _GEN_19745 : tag_1_46; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4797 = 7'h2f == index ? _GEN_19745 : tag_1_47; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4798 = 7'h30 == index ? _GEN_19745 : tag_1_48; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4799 = 7'h31 == index ? _GEN_19745 : tag_1_49; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4800 = 7'h32 == index ? _GEN_19745 : tag_1_50; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4801 = 7'h33 == index ? _GEN_19745 : tag_1_51; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4802 = 7'h34 == index ? _GEN_19745 : tag_1_52; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4803 = 7'h35 == index ? _GEN_19745 : tag_1_53; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4804 = 7'h36 == index ? _GEN_19745 : tag_1_54; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4805 = 7'h37 == index ? _GEN_19745 : tag_1_55; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4806 = 7'h38 == index ? _GEN_19745 : tag_1_56; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4807 = 7'h39 == index ? _GEN_19745 : tag_1_57; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4808 = 7'h3a == index ? _GEN_19745 : tag_1_58; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4809 = 7'h3b == index ? _GEN_19745 : tag_1_59; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4810 = 7'h3c == index ? _GEN_19745 : tag_1_60; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4811 = 7'h3d == index ? _GEN_19745 : tag_1_61; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4812 = 7'h3e == index ? _GEN_19745 : tag_1_62; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4813 = 7'h3f == index ? _GEN_19745 : tag_1_63; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4814 = 7'h40 == index ? _GEN_19745 : tag_1_64; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4815 = 7'h41 == index ? _GEN_19745 : tag_1_65; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4816 = 7'h42 == index ? _GEN_19745 : tag_1_66; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4817 = 7'h43 == index ? _GEN_19745 : tag_1_67; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4818 = 7'h44 == index ? _GEN_19745 : tag_1_68; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4819 = 7'h45 == index ? _GEN_19745 : tag_1_69; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4820 = 7'h46 == index ? _GEN_19745 : tag_1_70; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4821 = 7'h47 == index ? _GEN_19745 : tag_1_71; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4822 = 7'h48 == index ? _GEN_19745 : tag_1_72; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4823 = 7'h49 == index ? _GEN_19745 : tag_1_73; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4824 = 7'h4a == index ? _GEN_19745 : tag_1_74; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4825 = 7'h4b == index ? _GEN_19745 : tag_1_75; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4826 = 7'h4c == index ? _GEN_19745 : tag_1_76; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4827 = 7'h4d == index ? _GEN_19745 : tag_1_77; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4828 = 7'h4e == index ? _GEN_19745 : tag_1_78; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4829 = 7'h4f == index ? _GEN_19745 : tag_1_79; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4830 = 7'h50 == index ? _GEN_19745 : tag_1_80; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4831 = 7'h51 == index ? _GEN_19745 : tag_1_81; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4832 = 7'h52 == index ? _GEN_19745 : tag_1_82; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4833 = 7'h53 == index ? _GEN_19745 : tag_1_83; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4834 = 7'h54 == index ? _GEN_19745 : tag_1_84; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4835 = 7'h55 == index ? _GEN_19745 : tag_1_85; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4836 = 7'h56 == index ? _GEN_19745 : tag_1_86; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4837 = 7'h57 == index ? _GEN_19745 : tag_1_87; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4838 = 7'h58 == index ? _GEN_19745 : tag_1_88; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4839 = 7'h59 == index ? _GEN_19745 : tag_1_89; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4840 = 7'h5a == index ? _GEN_19745 : tag_1_90; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4841 = 7'h5b == index ? _GEN_19745 : tag_1_91; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4842 = 7'h5c == index ? _GEN_19745 : tag_1_92; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4843 = 7'h5d == index ? _GEN_19745 : tag_1_93; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4844 = 7'h5e == index ? _GEN_19745 : tag_1_94; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4845 = 7'h5f == index ? _GEN_19745 : tag_1_95; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4846 = 7'h60 == index ? _GEN_19745 : tag_1_96; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4847 = 7'h61 == index ? _GEN_19745 : tag_1_97; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4848 = 7'h62 == index ? _GEN_19745 : tag_1_98; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4849 = 7'h63 == index ? _GEN_19745 : tag_1_99; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4850 = 7'h64 == index ? _GEN_19745 : tag_1_100; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4851 = 7'h65 == index ? _GEN_19745 : tag_1_101; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4852 = 7'h66 == index ? _GEN_19745 : tag_1_102; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4853 = 7'h67 == index ? _GEN_19745 : tag_1_103; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4854 = 7'h68 == index ? _GEN_19745 : tag_1_104; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4855 = 7'h69 == index ? _GEN_19745 : tag_1_105; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4856 = 7'h6a == index ? _GEN_19745 : tag_1_106; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4857 = 7'h6b == index ? _GEN_19745 : tag_1_107; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4858 = 7'h6c == index ? _GEN_19745 : tag_1_108; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4859 = 7'h6d == index ? _GEN_19745 : tag_1_109; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4860 = 7'h6e == index ? _GEN_19745 : tag_1_110; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4861 = 7'h6f == index ? _GEN_19745 : tag_1_111; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4862 = 7'h70 == index ? _GEN_19745 : tag_1_112; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4863 = 7'h71 == index ? _GEN_19745 : tag_1_113; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4864 = 7'h72 == index ? _GEN_19745 : tag_1_114; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4865 = 7'h73 == index ? _GEN_19745 : tag_1_115; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4866 = 7'h74 == index ? _GEN_19745 : tag_1_116; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4867 = 7'h75 == index ? _GEN_19745 : tag_1_117; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4868 = 7'h76 == index ? _GEN_19745 : tag_1_118; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4869 = 7'h77 == index ? _GEN_19745 : tag_1_119; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4870 = 7'h78 == index ? _GEN_19745 : tag_1_120; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4871 = 7'h79 == index ? _GEN_19745 : tag_1_121; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4872 = 7'h7a == index ? _GEN_19745 : tag_1_122; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4873 = 7'h7b == index ? _GEN_19745 : tag_1_123; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4874 = 7'h7c == index ? _GEN_19745 : tag_1_124; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4875 = 7'h7d == index ? _GEN_19745 : tag_1_125; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4876 = 7'h7e == index ? _GEN_19745 : tag_1_126; // @[d_cache.scala 159:{30,30} 29:24]
  wire [31:0] _GEN_4877 = 7'h7f == index ? _GEN_19745 : tag_1_127; // @[d_cache.scala 159:{30,30} 29:24]
  wire  _GEN_4878 = _GEN_19748 | valid_1_0; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4879 = _GEN_19749 | valid_1_1; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4880 = _GEN_19750 | valid_1_2; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4881 = _GEN_19751 | valid_1_3; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4882 = _GEN_19752 | valid_1_4; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4883 = _GEN_19753 | valid_1_5; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4884 = _GEN_19754 | valid_1_6; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4885 = _GEN_19755 | valid_1_7; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4886 = _GEN_19756 | valid_1_8; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4887 = _GEN_19757 | valid_1_9; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4888 = _GEN_19758 | valid_1_10; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4889 = _GEN_19759 | valid_1_11; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4890 = _GEN_19760 | valid_1_12; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4891 = _GEN_19761 | valid_1_13; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4892 = _GEN_19762 | valid_1_14; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4893 = _GEN_19763 | valid_1_15; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4894 = _GEN_19764 | valid_1_16; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4895 = _GEN_19765 | valid_1_17; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4896 = _GEN_19766 | valid_1_18; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4897 = _GEN_19767 | valid_1_19; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4898 = _GEN_19768 | valid_1_20; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4899 = _GEN_19769 | valid_1_21; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4900 = _GEN_19770 | valid_1_22; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4901 = _GEN_19771 | valid_1_23; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4902 = _GEN_19772 | valid_1_24; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4903 = _GEN_19773 | valid_1_25; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4904 = _GEN_19774 | valid_1_26; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4905 = _GEN_19775 | valid_1_27; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4906 = _GEN_19776 | valid_1_28; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4907 = _GEN_19777 | valid_1_29; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4908 = _GEN_19778 | valid_1_30; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4909 = _GEN_19779 | valid_1_31; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4910 = _GEN_19780 | valid_1_32; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4911 = _GEN_19781 | valid_1_33; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4912 = _GEN_19782 | valid_1_34; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4913 = _GEN_19783 | valid_1_35; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4914 = _GEN_19784 | valid_1_36; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4915 = _GEN_19785 | valid_1_37; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4916 = _GEN_19786 | valid_1_38; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4917 = _GEN_19787 | valid_1_39; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4918 = _GEN_19788 | valid_1_40; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4919 = _GEN_19789 | valid_1_41; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4920 = _GEN_19790 | valid_1_42; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4921 = _GEN_19791 | valid_1_43; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4922 = _GEN_19792 | valid_1_44; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4923 = _GEN_19793 | valid_1_45; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4924 = _GEN_19794 | valid_1_46; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4925 = _GEN_19795 | valid_1_47; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4926 = _GEN_19796 | valid_1_48; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4927 = _GEN_19797 | valid_1_49; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4928 = _GEN_19798 | valid_1_50; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4929 = _GEN_19799 | valid_1_51; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4930 = _GEN_19800 | valid_1_52; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4931 = _GEN_19801 | valid_1_53; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4932 = _GEN_19802 | valid_1_54; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4933 = _GEN_19803 | valid_1_55; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4934 = _GEN_19804 | valid_1_56; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4935 = _GEN_19805 | valid_1_57; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4936 = _GEN_19806 | valid_1_58; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4937 = _GEN_19807 | valid_1_59; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4938 = _GEN_19808 | valid_1_60; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4939 = _GEN_19809 | valid_1_61; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4940 = _GEN_19810 | valid_1_62; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4941 = _GEN_19811 | valid_1_63; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4942 = _GEN_19812 | valid_1_64; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4943 = _GEN_19813 | valid_1_65; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4944 = _GEN_19814 | valid_1_66; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4945 = _GEN_19815 | valid_1_67; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4946 = _GEN_19816 | valid_1_68; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4947 = _GEN_19817 | valid_1_69; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4948 = _GEN_19818 | valid_1_70; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4949 = _GEN_19819 | valid_1_71; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4950 = _GEN_19820 | valid_1_72; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4951 = _GEN_19821 | valid_1_73; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4952 = _GEN_19822 | valid_1_74; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4953 = _GEN_19823 | valid_1_75; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4954 = _GEN_19824 | valid_1_76; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4955 = _GEN_19825 | valid_1_77; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4956 = _GEN_19826 | valid_1_78; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4957 = _GEN_19827 | valid_1_79; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4958 = _GEN_19828 | valid_1_80; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4959 = _GEN_19829 | valid_1_81; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4960 = _GEN_19830 | valid_1_82; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4961 = _GEN_19831 | valid_1_83; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4962 = _GEN_19832 | valid_1_84; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4963 = _GEN_19833 | valid_1_85; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4964 = _GEN_19834 | valid_1_86; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4965 = _GEN_19835 | valid_1_87; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4966 = _GEN_19836 | valid_1_88; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4967 = _GEN_19837 | valid_1_89; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4968 = _GEN_19838 | valid_1_90; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4969 = _GEN_19839 | valid_1_91; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4970 = _GEN_19840 | valid_1_92; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4971 = _GEN_19841 | valid_1_93; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4972 = _GEN_19842 | valid_1_94; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4973 = _GEN_19843 | valid_1_95; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4974 = _GEN_19844 | valid_1_96; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4975 = _GEN_19845 | valid_1_97; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4976 = _GEN_19846 | valid_1_98; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4977 = _GEN_19847 | valid_1_99; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4978 = _GEN_19848 | valid_1_100; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4979 = _GEN_19849 | valid_1_101; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4980 = _GEN_19850 | valid_1_102; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4981 = _GEN_19851 | valid_1_103; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4982 = _GEN_19852 | valid_1_104; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4983 = _GEN_19853 | valid_1_105; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4984 = _GEN_19854 | valid_1_106; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4985 = _GEN_19855 | valid_1_107; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4986 = _GEN_19856 | valid_1_108; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4987 = _GEN_19857 | valid_1_109; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4988 = _GEN_19858 | valid_1_110; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4989 = _GEN_19859 | valid_1_111; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4990 = _GEN_19860 | valid_1_112; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4991 = _GEN_19861 | valid_1_113; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4992 = _GEN_19862 | valid_1_114; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4993 = _GEN_19863 | valid_1_115; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4994 = _GEN_19864 | valid_1_116; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4995 = _GEN_19865 | valid_1_117; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4996 = _GEN_19866 | valid_1_118; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4997 = _GEN_19867 | valid_1_119; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4998 = _GEN_19868 | valid_1_120; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_4999 = _GEN_19869 | valid_1_121; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_5000 = _GEN_19870 | valid_1_122; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_5001 = _GEN_19871 | valid_1_123; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_5002 = _GEN_19872 | valid_1_124; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_5003 = _GEN_19873 | valid_1_125; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_5004 = _GEN_19874 | valid_1_126; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _GEN_5005 = _GEN_19875 | valid_1_127; // @[d_cache.scala 160:{32,32} 31:26]
  wire  _T_26 = ~quene; // @[d_cache.scala 163:27]
  wire [41:0] _write_back_addr_T_1 = {_GEN_127,index,3'h0}; // @[Cat.scala 31:58]
  wire  _GEN_5262 = 7'h0 == index ? 1'h0 : dirty_0_0; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5263 = 7'h1 == index ? 1'h0 : dirty_0_1; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5264 = 7'h2 == index ? 1'h0 : dirty_0_2; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5265 = 7'h3 == index ? 1'h0 : dirty_0_3; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5266 = 7'h4 == index ? 1'h0 : dirty_0_4; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5267 = 7'h5 == index ? 1'h0 : dirty_0_5; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5268 = 7'h6 == index ? 1'h0 : dirty_0_6; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5269 = 7'h7 == index ? 1'h0 : dirty_0_7; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5270 = 7'h8 == index ? 1'h0 : dirty_0_8; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5271 = 7'h9 == index ? 1'h0 : dirty_0_9; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5272 = 7'ha == index ? 1'h0 : dirty_0_10; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5273 = 7'hb == index ? 1'h0 : dirty_0_11; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5274 = 7'hc == index ? 1'h0 : dirty_0_12; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5275 = 7'hd == index ? 1'h0 : dirty_0_13; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5276 = 7'he == index ? 1'h0 : dirty_0_14; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5277 = 7'hf == index ? 1'h0 : dirty_0_15; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5278 = 7'h10 == index ? 1'h0 : dirty_0_16; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5279 = 7'h11 == index ? 1'h0 : dirty_0_17; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5280 = 7'h12 == index ? 1'h0 : dirty_0_18; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5281 = 7'h13 == index ? 1'h0 : dirty_0_19; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5282 = 7'h14 == index ? 1'h0 : dirty_0_20; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5283 = 7'h15 == index ? 1'h0 : dirty_0_21; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5284 = 7'h16 == index ? 1'h0 : dirty_0_22; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5285 = 7'h17 == index ? 1'h0 : dirty_0_23; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5286 = 7'h18 == index ? 1'h0 : dirty_0_24; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5287 = 7'h19 == index ? 1'h0 : dirty_0_25; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5288 = 7'h1a == index ? 1'h0 : dirty_0_26; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5289 = 7'h1b == index ? 1'h0 : dirty_0_27; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5290 = 7'h1c == index ? 1'h0 : dirty_0_28; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5291 = 7'h1d == index ? 1'h0 : dirty_0_29; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5292 = 7'h1e == index ? 1'h0 : dirty_0_30; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5293 = 7'h1f == index ? 1'h0 : dirty_0_31; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5294 = 7'h20 == index ? 1'h0 : dirty_0_32; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5295 = 7'h21 == index ? 1'h0 : dirty_0_33; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5296 = 7'h22 == index ? 1'h0 : dirty_0_34; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5297 = 7'h23 == index ? 1'h0 : dirty_0_35; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5298 = 7'h24 == index ? 1'h0 : dirty_0_36; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5299 = 7'h25 == index ? 1'h0 : dirty_0_37; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5300 = 7'h26 == index ? 1'h0 : dirty_0_38; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5301 = 7'h27 == index ? 1'h0 : dirty_0_39; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5302 = 7'h28 == index ? 1'h0 : dirty_0_40; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5303 = 7'h29 == index ? 1'h0 : dirty_0_41; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5304 = 7'h2a == index ? 1'h0 : dirty_0_42; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5305 = 7'h2b == index ? 1'h0 : dirty_0_43; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5306 = 7'h2c == index ? 1'h0 : dirty_0_44; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5307 = 7'h2d == index ? 1'h0 : dirty_0_45; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5308 = 7'h2e == index ? 1'h0 : dirty_0_46; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5309 = 7'h2f == index ? 1'h0 : dirty_0_47; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5310 = 7'h30 == index ? 1'h0 : dirty_0_48; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5311 = 7'h31 == index ? 1'h0 : dirty_0_49; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5312 = 7'h32 == index ? 1'h0 : dirty_0_50; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5313 = 7'h33 == index ? 1'h0 : dirty_0_51; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5314 = 7'h34 == index ? 1'h0 : dirty_0_52; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5315 = 7'h35 == index ? 1'h0 : dirty_0_53; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5316 = 7'h36 == index ? 1'h0 : dirty_0_54; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5317 = 7'h37 == index ? 1'h0 : dirty_0_55; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5318 = 7'h38 == index ? 1'h0 : dirty_0_56; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5319 = 7'h39 == index ? 1'h0 : dirty_0_57; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5320 = 7'h3a == index ? 1'h0 : dirty_0_58; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5321 = 7'h3b == index ? 1'h0 : dirty_0_59; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5322 = 7'h3c == index ? 1'h0 : dirty_0_60; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5323 = 7'h3d == index ? 1'h0 : dirty_0_61; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5324 = 7'h3e == index ? 1'h0 : dirty_0_62; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5325 = 7'h3f == index ? 1'h0 : dirty_0_63; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5326 = 7'h40 == index ? 1'h0 : dirty_0_64; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5327 = 7'h41 == index ? 1'h0 : dirty_0_65; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5328 = 7'h42 == index ? 1'h0 : dirty_0_66; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5329 = 7'h43 == index ? 1'h0 : dirty_0_67; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5330 = 7'h44 == index ? 1'h0 : dirty_0_68; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5331 = 7'h45 == index ? 1'h0 : dirty_0_69; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5332 = 7'h46 == index ? 1'h0 : dirty_0_70; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5333 = 7'h47 == index ? 1'h0 : dirty_0_71; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5334 = 7'h48 == index ? 1'h0 : dirty_0_72; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5335 = 7'h49 == index ? 1'h0 : dirty_0_73; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5336 = 7'h4a == index ? 1'h0 : dirty_0_74; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5337 = 7'h4b == index ? 1'h0 : dirty_0_75; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5338 = 7'h4c == index ? 1'h0 : dirty_0_76; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5339 = 7'h4d == index ? 1'h0 : dirty_0_77; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5340 = 7'h4e == index ? 1'h0 : dirty_0_78; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5341 = 7'h4f == index ? 1'h0 : dirty_0_79; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5342 = 7'h50 == index ? 1'h0 : dirty_0_80; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5343 = 7'h51 == index ? 1'h0 : dirty_0_81; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5344 = 7'h52 == index ? 1'h0 : dirty_0_82; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5345 = 7'h53 == index ? 1'h0 : dirty_0_83; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5346 = 7'h54 == index ? 1'h0 : dirty_0_84; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5347 = 7'h55 == index ? 1'h0 : dirty_0_85; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5348 = 7'h56 == index ? 1'h0 : dirty_0_86; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5349 = 7'h57 == index ? 1'h0 : dirty_0_87; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5350 = 7'h58 == index ? 1'h0 : dirty_0_88; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5351 = 7'h59 == index ? 1'h0 : dirty_0_89; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5352 = 7'h5a == index ? 1'h0 : dirty_0_90; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5353 = 7'h5b == index ? 1'h0 : dirty_0_91; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5354 = 7'h5c == index ? 1'h0 : dirty_0_92; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5355 = 7'h5d == index ? 1'h0 : dirty_0_93; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5356 = 7'h5e == index ? 1'h0 : dirty_0_94; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5357 = 7'h5f == index ? 1'h0 : dirty_0_95; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5358 = 7'h60 == index ? 1'h0 : dirty_0_96; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5359 = 7'h61 == index ? 1'h0 : dirty_0_97; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5360 = 7'h62 == index ? 1'h0 : dirty_0_98; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5361 = 7'h63 == index ? 1'h0 : dirty_0_99; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5362 = 7'h64 == index ? 1'h0 : dirty_0_100; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5363 = 7'h65 == index ? 1'h0 : dirty_0_101; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5364 = 7'h66 == index ? 1'h0 : dirty_0_102; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5365 = 7'h67 == index ? 1'h0 : dirty_0_103; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5366 = 7'h68 == index ? 1'h0 : dirty_0_104; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5367 = 7'h69 == index ? 1'h0 : dirty_0_105; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5368 = 7'h6a == index ? 1'h0 : dirty_0_106; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5369 = 7'h6b == index ? 1'h0 : dirty_0_107; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5370 = 7'h6c == index ? 1'h0 : dirty_0_108; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5371 = 7'h6d == index ? 1'h0 : dirty_0_109; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5372 = 7'h6e == index ? 1'h0 : dirty_0_110; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5373 = 7'h6f == index ? 1'h0 : dirty_0_111; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5374 = 7'h70 == index ? 1'h0 : dirty_0_112; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5375 = 7'h71 == index ? 1'h0 : dirty_0_113; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5376 = 7'h72 == index ? 1'h0 : dirty_0_114; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5377 = 7'h73 == index ? 1'h0 : dirty_0_115; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5378 = 7'h74 == index ? 1'h0 : dirty_0_116; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5379 = 7'h75 == index ? 1'h0 : dirty_0_117; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5380 = 7'h76 == index ? 1'h0 : dirty_0_118; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5381 = 7'h77 == index ? 1'h0 : dirty_0_119; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5382 = 7'h78 == index ? 1'h0 : dirty_0_120; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5383 = 7'h79 == index ? 1'h0 : dirty_0_121; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5384 = 7'h7a == index ? 1'h0 : dirty_0_122; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5385 = 7'h7b == index ? 1'h0 : dirty_0_123; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5386 = 7'h7c == index ? 1'h0 : dirty_0_124; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5387 = 7'h7d == index ? 1'h0 : dirty_0_125; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5388 = 7'h7e == index ? 1'h0 : dirty_0_126; // @[d_cache.scala 170:{40,40} 32:26]
  wire  _GEN_5389 = 7'h7f == index ? 1'h0 : dirty_0_127; // @[d_cache.scala 170:{40,40} 32:26]
  wire [63:0] _GEN_5902 = _GEN_645 ? _GEN_904 : write_back_data; // @[d_cache.scala 165:47 166:41 37:34]
  wire [41:0] _GEN_5903 = _GEN_645 ? _write_back_addr_T_1 : {{10'd0}, write_back_addr}; // @[d_cache.scala 165:47 167:41 38:34]
  wire [63:0] _GEN_5904 = _GEN_645 ? _GEN_4238 : _GEN_4238; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5905 = _GEN_645 ? _GEN_4239 : _GEN_4239; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5906 = _GEN_645 ? _GEN_4240 : _GEN_4240; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5907 = _GEN_645 ? _GEN_4241 : _GEN_4241; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5908 = _GEN_645 ? _GEN_4242 : _GEN_4242; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5909 = _GEN_645 ? _GEN_4243 : _GEN_4243; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5910 = _GEN_645 ? _GEN_4244 : _GEN_4244; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5911 = _GEN_645 ? _GEN_4245 : _GEN_4245; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5912 = _GEN_645 ? _GEN_4246 : _GEN_4246; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5913 = _GEN_645 ? _GEN_4247 : _GEN_4247; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5914 = _GEN_645 ? _GEN_4248 : _GEN_4248; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5915 = _GEN_645 ? _GEN_4249 : _GEN_4249; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5916 = _GEN_645 ? _GEN_4250 : _GEN_4250; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5917 = _GEN_645 ? _GEN_4251 : _GEN_4251; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5918 = _GEN_645 ? _GEN_4252 : _GEN_4252; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5919 = _GEN_645 ? _GEN_4253 : _GEN_4253; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5920 = _GEN_645 ? _GEN_4254 : _GEN_4254; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5921 = _GEN_645 ? _GEN_4255 : _GEN_4255; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5922 = _GEN_645 ? _GEN_4256 : _GEN_4256; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5923 = _GEN_645 ? _GEN_4257 : _GEN_4257; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5924 = _GEN_645 ? _GEN_4258 : _GEN_4258; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5925 = _GEN_645 ? _GEN_4259 : _GEN_4259; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5926 = _GEN_645 ? _GEN_4260 : _GEN_4260; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5927 = _GEN_645 ? _GEN_4261 : _GEN_4261; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5928 = _GEN_645 ? _GEN_4262 : _GEN_4262; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5929 = _GEN_645 ? _GEN_4263 : _GEN_4263; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5930 = _GEN_645 ? _GEN_4264 : _GEN_4264; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5931 = _GEN_645 ? _GEN_4265 : _GEN_4265; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5932 = _GEN_645 ? _GEN_4266 : _GEN_4266; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5933 = _GEN_645 ? _GEN_4267 : _GEN_4267; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5934 = _GEN_645 ? _GEN_4268 : _GEN_4268; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5935 = _GEN_645 ? _GEN_4269 : _GEN_4269; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5936 = _GEN_645 ? _GEN_4270 : _GEN_4270; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5937 = _GEN_645 ? _GEN_4271 : _GEN_4271; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5938 = _GEN_645 ? _GEN_4272 : _GEN_4272; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5939 = _GEN_645 ? _GEN_4273 : _GEN_4273; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5940 = _GEN_645 ? _GEN_4274 : _GEN_4274; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5941 = _GEN_645 ? _GEN_4275 : _GEN_4275; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5942 = _GEN_645 ? _GEN_4276 : _GEN_4276; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5943 = _GEN_645 ? _GEN_4277 : _GEN_4277; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5944 = _GEN_645 ? _GEN_4278 : _GEN_4278; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5945 = _GEN_645 ? _GEN_4279 : _GEN_4279; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5946 = _GEN_645 ? _GEN_4280 : _GEN_4280; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5947 = _GEN_645 ? _GEN_4281 : _GEN_4281; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5948 = _GEN_645 ? _GEN_4282 : _GEN_4282; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5949 = _GEN_645 ? _GEN_4283 : _GEN_4283; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5950 = _GEN_645 ? _GEN_4284 : _GEN_4284; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5951 = _GEN_645 ? _GEN_4285 : _GEN_4285; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5952 = _GEN_645 ? _GEN_4286 : _GEN_4286; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5953 = _GEN_645 ? _GEN_4287 : _GEN_4287; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5954 = _GEN_645 ? _GEN_4288 : _GEN_4288; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5955 = _GEN_645 ? _GEN_4289 : _GEN_4289; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5956 = _GEN_645 ? _GEN_4290 : _GEN_4290; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5957 = _GEN_645 ? _GEN_4291 : _GEN_4291; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5958 = _GEN_645 ? _GEN_4292 : _GEN_4292; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5959 = _GEN_645 ? _GEN_4293 : _GEN_4293; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5960 = _GEN_645 ? _GEN_4294 : _GEN_4294; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5961 = _GEN_645 ? _GEN_4295 : _GEN_4295; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5962 = _GEN_645 ? _GEN_4296 : _GEN_4296; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5963 = _GEN_645 ? _GEN_4297 : _GEN_4297; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5964 = _GEN_645 ? _GEN_4298 : _GEN_4298; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5965 = _GEN_645 ? _GEN_4299 : _GEN_4299; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5966 = _GEN_645 ? _GEN_4300 : _GEN_4300; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5967 = _GEN_645 ? _GEN_4301 : _GEN_4301; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5968 = _GEN_645 ? _GEN_4302 : _GEN_4302; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5969 = _GEN_645 ? _GEN_4303 : _GEN_4303; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5970 = _GEN_645 ? _GEN_4304 : _GEN_4304; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5971 = _GEN_645 ? _GEN_4305 : _GEN_4305; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5972 = _GEN_645 ? _GEN_4306 : _GEN_4306; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5973 = _GEN_645 ? _GEN_4307 : _GEN_4307; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5974 = _GEN_645 ? _GEN_4308 : _GEN_4308; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5975 = _GEN_645 ? _GEN_4309 : _GEN_4309; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5976 = _GEN_645 ? _GEN_4310 : _GEN_4310; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5977 = _GEN_645 ? _GEN_4311 : _GEN_4311; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5978 = _GEN_645 ? _GEN_4312 : _GEN_4312; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5979 = _GEN_645 ? _GEN_4313 : _GEN_4313; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5980 = _GEN_645 ? _GEN_4314 : _GEN_4314; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5981 = _GEN_645 ? _GEN_4315 : _GEN_4315; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5982 = _GEN_645 ? _GEN_4316 : _GEN_4316; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5983 = _GEN_645 ? _GEN_4317 : _GEN_4317; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5984 = _GEN_645 ? _GEN_4318 : _GEN_4318; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5985 = _GEN_645 ? _GEN_4319 : _GEN_4319; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5986 = _GEN_645 ? _GEN_4320 : _GEN_4320; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5987 = _GEN_645 ? _GEN_4321 : _GEN_4321; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5988 = _GEN_645 ? _GEN_4322 : _GEN_4322; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5989 = _GEN_645 ? _GEN_4323 : _GEN_4323; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5990 = _GEN_645 ? _GEN_4324 : _GEN_4324; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5991 = _GEN_645 ? _GEN_4325 : _GEN_4325; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5992 = _GEN_645 ? _GEN_4326 : _GEN_4326; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5993 = _GEN_645 ? _GEN_4327 : _GEN_4327; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5994 = _GEN_645 ? _GEN_4328 : _GEN_4328; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5995 = _GEN_645 ? _GEN_4329 : _GEN_4329; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5996 = _GEN_645 ? _GEN_4330 : _GEN_4330; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5997 = _GEN_645 ? _GEN_4331 : _GEN_4331; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5998 = _GEN_645 ? _GEN_4332 : _GEN_4332; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_5999 = _GEN_645 ? _GEN_4333 : _GEN_4333; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6000 = _GEN_645 ? _GEN_4334 : _GEN_4334; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6001 = _GEN_645 ? _GEN_4335 : _GEN_4335; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6002 = _GEN_645 ? _GEN_4336 : _GEN_4336; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6003 = _GEN_645 ? _GEN_4337 : _GEN_4337; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6004 = _GEN_645 ? _GEN_4338 : _GEN_4338; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6005 = _GEN_645 ? _GEN_4339 : _GEN_4339; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6006 = _GEN_645 ? _GEN_4340 : _GEN_4340; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6007 = _GEN_645 ? _GEN_4341 : _GEN_4341; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6008 = _GEN_645 ? _GEN_4342 : _GEN_4342; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6009 = _GEN_645 ? _GEN_4343 : _GEN_4343; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6010 = _GEN_645 ? _GEN_4344 : _GEN_4344; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6011 = _GEN_645 ? _GEN_4345 : _GEN_4345; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6012 = _GEN_645 ? _GEN_4346 : _GEN_4346; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6013 = _GEN_645 ? _GEN_4347 : _GEN_4347; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6014 = _GEN_645 ? _GEN_4348 : _GEN_4348; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6015 = _GEN_645 ? _GEN_4349 : _GEN_4349; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6016 = _GEN_645 ? _GEN_4350 : _GEN_4350; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6017 = _GEN_645 ? _GEN_4351 : _GEN_4351; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6018 = _GEN_645 ? _GEN_4352 : _GEN_4352; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6019 = _GEN_645 ? _GEN_4353 : _GEN_4353; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6020 = _GEN_645 ? _GEN_4354 : _GEN_4354; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6021 = _GEN_645 ? _GEN_4355 : _GEN_4355; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6022 = _GEN_645 ? _GEN_4356 : _GEN_4356; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6023 = _GEN_645 ? _GEN_4357 : _GEN_4357; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6024 = _GEN_645 ? _GEN_4358 : _GEN_4358; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6025 = _GEN_645 ? _GEN_4359 : _GEN_4359; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6026 = _GEN_645 ? _GEN_4360 : _GEN_4360; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6027 = _GEN_645 ? _GEN_4361 : _GEN_4361; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6028 = _GEN_645 ? _GEN_4362 : _GEN_4362; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6029 = _GEN_645 ? _GEN_4363 : _GEN_4363; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6030 = _GEN_645 ? _GEN_4364 : _GEN_4364; // @[d_cache.scala 165:47]
  wire [63:0] _GEN_6031 = _GEN_645 ? _GEN_4365 : _GEN_4365; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6032 = _GEN_645 ? _GEN_4366 : _GEN_4366; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6033 = _GEN_645 ? _GEN_4367 : _GEN_4367; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6034 = _GEN_645 ? _GEN_4368 : _GEN_4368; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6035 = _GEN_645 ? _GEN_4369 : _GEN_4369; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6036 = _GEN_645 ? _GEN_4370 : _GEN_4370; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6037 = _GEN_645 ? _GEN_4371 : _GEN_4371; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6038 = _GEN_645 ? _GEN_4372 : _GEN_4372; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6039 = _GEN_645 ? _GEN_4373 : _GEN_4373; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6040 = _GEN_645 ? _GEN_4374 : _GEN_4374; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6041 = _GEN_645 ? _GEN_4375 : _GEN_4375; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6042 = _GEN_645 ? _GEN_4376 : _GEN_4376; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6043 = _GEN_645 ? _GEN_4377 : _GEN_4377; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6044 = _GEN_645 ? _GEN_4378 : _GEN_4378; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6045 = _GEN_645 ? _GEN_4379 : _GEN_4379; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6046 = _GEN_645 ? _GEN_4380 : _GEN_4380; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6047 = _GEN_645 ? _GEN_4381 : _GEN_4381; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6048 = _GEN_645 ? _GEN_4382 : _GEN_4382; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6049 = _GEN_645 ? _GEN_4383 : _GEN_4383; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6050 = _GEN_645 ? _GEN_4384 : _GEN_4384; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6051 = _GEN_645 ? _GEN_4385 : _GEN_4385; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6052 = _GEN_645 ? _GEN_4386 : _GEN_4386; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6053 = _GEN_645 ? _GEN_4387 : _GEN_4387; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6054 = _GEN_645 ? _GEN_4388 : _GEN_4388; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6055 = _GEN_645 ? _GEN_4389 : _GEN_4389; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6056 = _GEN_645 ? _GEN_4390 : _GEN_4390; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6057 = _GEN_645 ? _GEN_4391 : _GEN_4391; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6058 = _GEN_645 ? _GEN_4392 : _GEN_4392; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6059 = _GEN_645 ? _GEN_4393 : _GEN_4393; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6060 = _GEN_645 ? _GEN_4394 : _GEN_4394; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6061 = _GEN_645 ? _GEN_4395 : _GEN_4395; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6062 = _GEN_645 ? _GEN_4396 : _GEN_4396; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6063 = _GEN_645 ? _GEN_4397 : _GEN_4397; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6064 = _GEN_645 ? _GEN_4398 : _GEN_4398; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6065 = _GEN_645 ? _GEN_4399 : _GEN_4399; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6066 = _GEN_645 ? _GEN_4400 : _GEN_4400; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6067 = _GEN_645 ? _GEN_4401 : _GEN_4401; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6068 = _GEN_645 ? _GEN_4402 : _GEN_4402; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6069 = _GEN_645 ? _GEN_4403 : _GEN_4403; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6070 = _GEN_645 ? _GEN_4404 : _GEN_4404; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6071 = _GEN_645 ? _GEN_4405 : _GEN_4405; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6072 = _GEN_645 ? _GEN_4406 : _GEN_4406; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6073 = _GEN_645 ? _GEN_4407 : _GEN_4407; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6074 = _GEN_645 ? _GEN_4408 : _GEN_4408; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6075 = _GEN_645 ? _GEN_4409 : _GEN_4409; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6076 = _GEN_645 ? _GEN_4410 : _GEN_4410; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6077 = _GEN_645 ? _GEN_4411 : _GEN_4411; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6078 = _GEN_645 ? _GEN_4412 : _GEN_4412; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6079 = _GEN_645 ? _GEN_4413 : _GEN_4413; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6080 = _GEN_645 ? _GEN_4414 : _GEN_4414; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6081 = _GEN_645 ? _GEN_4415 : _GEN_4415; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6082 = _GEN_645 ? _GEN_4416 : _GEN_4416; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6083 = _GEN_645 ? _GEN_4417 : _GEN_4417; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6084 = _GEN_645 ? _GEN_4418 : _GEN_4418; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6085 = _GEN_645 ? _GEN_4419 : _GEN_4419; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6086 = _GEN_645 ? _GEN_4420 : _GEN_4420; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6087 = _GEN_645 ? _GEN_4421 : _GEN_4421; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6088 = _GEN_645 ? _GEN_4422 : _GEN_4422; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6089 = _GEN_645 ? _GEN_4423 : _GEN_4423; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6090 = _GEN_645 ? _GEN_4424 : _GEN_4424; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6091 = _GEN_645 ? _GEN_4425 : _GEN_4425; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6092 = _GEN_645 ? _GEN_4426 : _GEN_4426; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6093 = _GEN_645 ? _GEN_4427 : _GEN_4427; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6094 = _GEN_645 ? _GEN_4428 : _GEN_4428; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6095 = _GEN_645 ? _GEN_4429 : _GEN_4429; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6096 = _GEN_645 ? _GEN_4430 : _GEN_4430; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6097 = _GEN_645 ? _GEN_4431 : _GEN_4431; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6098 = _GEN_645 ? _GEN_4432 : _GEN_4432; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6099 = _GEN_645 ? _GEN_4433 : _GEN_4433; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6100 = _GEN_645 ? _GEN_4434 : _GEN_4434; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6101 = _GEN_645 ? _GEN_4435 : _GEN_4435; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6102 = _GEN_645 ? _GEN_4436 : _GEN_4436; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6103 = _GEN_645 ? _GEN_4437 : _GEN_4437; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6104 = _GEN_645 ? _GEN_4438 : _GEN_4438; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6105 = _GEN_645 ? _GEN_4439 : _GEN_4439; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6106 = _GEN_645 ? _GEN_4440 : _GEN_4440; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6107 = _GEN_645 ? _GEN_4441 : _GEN_4441; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6108 = _GEN_645 ? _GEN_4442 : _GEN_4442; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6109 = _GEN_645 ? _GEN_4443 : _GEN_4443; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6110 = _GEN_645 ? _GEN_4444 : _GEN_4444; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6111 = _GEN_645 ? _GEN_4445 : _GEN_4445; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6112 = _GEN_645 ? _GEN_4446 : _GEN_4446; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6113 = _GEN_645 ? _GEN_4447 : _GEN_4447; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6114 = _GEN_645 ? _GEN_4448 : _GEN_4448; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6115 = _GEN_645 ? _GEN_4449 : _GEN_4449; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6116 = _GEN_645 ? _GEN_4450 : _GEN_4450; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6117 = _GEN_645 ? _GEN_4451 : _GEN_4451; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6118 = _GEN_645 ? _GEN_4452 : _GEN_4452; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6119 = _GEN_645 ? _GEN_4453 : _GEN_4453; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6120 = _GEN_645 ? _GEN_4454 : _GEN_4454; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6121 = _GEN_645 ? _GEN_4455 : _GEN_4455; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6122 = _GEN_645 ? _GEN_4456 : _GEN_4456; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6123 = _GEN_645 ? _GEN_4457 : _GEN_4457; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6124 = _GEN_645 ? _GEN_4458 : _GEN_4458; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6125 = _GEN_645 ? _GEN_4459 : _GEN_4459; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6126 = _GEN_645 ? _GEN_4460 : _GEN_4460; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6127 = _GEN_645 ? _GEN_4461 : _GEN_4461; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6128 = _GEN_645 ? _GEN_4462 : _GEN_4462; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6129 = _GEN_645 ? _GEN_4463 : _GEN_4463; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6130 = _GEN_645 ? _GEN_4464 : _GEN_4464; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6131 = _GEN_645 ? _GEN_4465 : _GEN_4465; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6132 = _GEN_645 ? _GEN_4466 : _GEN_4466; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6133 = _GEN_645 ? _GEN_4467 : _GEN_4467; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6134 = _GEN_645 ? _GEN_4468 : _GEN_4468; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6135 = _GEN_645 ? _GEN_4469 : _GEN_4469; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6136 = _GEN_645 ? _GEN_4470 : _GEN_4470; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6137 = _GEN_645 ? _GEN_4471 : _GEN_4471; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6138 = _GEN_645 ? _GEN_4472 : _GEN_4472; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6139 = _GEN_645 ? _GEN_4473 : _GEN_4473; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6140 = _GEN_645 ? _GEN_4474 : _GEN_4474; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6141 = _GEN_645 ? _GEN_4475 : _GEN_4475; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6142 = _GEN_645 ? _GEN_4476 : _GEN_4476; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6143 = _GEN_645 ? _GEN_4477 : _GEN_4477; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6144 = _GEN_645 ? _GEN_4478 : _GEN_4478; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6145 = _GEN_645 ? _GEN_4479 : _GEN_4479; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6146 = _GEN_645 ? _GEN_4480 : _GEN_4480; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6147 = _GEN_645 ? _GEN_4481 : _GEN_4481; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6148 = _GEN_645 ? _GEN_4482 : _GEN_4482; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6149 = _GEN_645 ? _GEN_4483 : _GEN_4483; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6150 = _GEN_645 ? _GEN_4484 : _GEN_4484; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6151 = _GEN_645 ? _GEN_4485 : _GEN_4485; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6152 = _GEN_645 ? _GEN_4486 : _GEN_4486; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6153 = _GEN_645 ? _GEN_4487 : _GEN_4487; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6154 = _GEN_645 ? _GEN_4488 : _GEN_4488; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6155 = _GEN_645 ? _GEN_4489 : _GEN_4489; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6156 = _GEN_645 ? _GEN_4490 : _GEN_4490; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6157 = _GEN_645 ? _GEN_4491 : _GEN_4491; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6158 = _GEN_645 ? _GEN_4492 : _GEN_4492; // @[d_cache.scala 165:47]
  wire [31:0] _GEN_6159 = _GEN_645 ? _GEN_4493 : _GEN_4493; // @[d_cache.scala 165:47]
  wire  _GEN_6160 = _GEN_645 ? _GEN_5262 : dirty_0_0; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6161 = _GEN_645 ? _GEN_5263 : dirty_0_1; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6162 = _GEN_645 ? _GEN_5264 : dirty_0_2; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6163 = _GEN_645 ? _GEN_5265 : dirty_0_3; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6164 = _GEN_645 ? _GEN_5266 : dirty_0_4; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6165 = _GEN_645 ? _GEN_5267 : dirty_0_5; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6166 = _GEN_645 ? _GEN_5268 : dirty_0_6; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6167 = _GEN_645 ? _GEN_5269 : dirty_0_7; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6168 = _GEN_645 ? _GEN_5270 : dirty_0_8; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6169 = _GEN_645 ? _GEN_5271 : dirty_0_9; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6170 = _GEN_645 ? _GEN_5272 : dirty_0_10; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6171 = _GEN_645 ? _GEN_5273 : dirty_0_11; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6172 = _GEN_645 ? _GEN_5274 : dirty_0_12; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6173 = _GEN_645 ? _GEN_5275 : dirty_0_13; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6174 = _GEN_645 ? _GEN_5276 : dirty_0_14; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6175 = _GEN_645 ? _GEN_5277 : dirty_0_15; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6176 = _GEN_645 ? _GEN_5278 : dirty_0_16; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6177 = _GEN_645 ? _GEN_5279 : dirty_0_17; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6178 = _GEN_645 ? _GEN_5280 : dirty_0_18; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6179 = _GEN_645 ? _GEN_5281 : dirty_0_19; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6180 = _GEN_645 ? _GEN_5282 : dirty_0_20; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6181 = _GEN_645 ? _GEN_5283 : dirty_0_21; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6182 = _GEN_645 ? _GEN_5284 : dirty_0_22; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6183 = _GEN_645 ? _GEN_5285 : dirty_0_23; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6184 = _GEN_645 ? _GEN_5286 : dirty_0_24; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6185 = _GEN_645 ? _GEN_5287 : dirty_0_25; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6186 = _GEN_645 ? _GEN_5288 : dirty_0_26; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6187 = _GEN_645 ? _GEN_5289 : dirty_0_27; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6188 = _GEN_645 ? _GEN_5290 : dirty_0_28; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6189 = _GEN_645 ? _GEN_5291 : dirty_0_29; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6190 = _GEN_645 ? _GEN_5292 : dirty_0_30; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6191 = _GEN_645 ? _GEN_5293 : dirty_0_31; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6192 = _GEN_645 ? _GEN_5294 : dirty_0_32; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6193 = _GEN_645 ? _GEN_5295 : dirty_0_33; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6194 = _GEN_645 ? _GEN_5296 : dirty_0_34; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6195 = _GEN_645 ? _GEN_5297 : dirty_0_35; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6196 = _GEN_645 ? _GEN_5298 : dirty_0_36; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6197 = _GEN_645 ? _GEN_5299 : dirty_0_37; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6198 = _GEN_645 ? _GEN_5300 : dirty_0_38; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6199 = _GEN_645 ? _GEN_5301 : dirty_0_39; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6200 = _GEN_645 ? _GEN_5302 : dirty_0_40; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6201 = _GEN_645 ? _GEN_5303 : dirty_0_41; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6202 = _GEN_645 ? _GEN_5304 : dirty_0_42; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6203 = _GEN_645 ? _GEN_5305 : dirty_0_43; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6204 = _GEN_645 ? _GEN_5306 : dirty_0_44; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6205 = _GEN_645 ? _GEN_5307 : dirty_0_45; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6206 = _GEN_645 ? _GEN_5308 : dirty_0_46; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6207 = _GEN_645 ? _GEN_5309 : dirty_0_47; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6208 = _GEN_645 ? _GEN_5310 : dirty_0_48; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6209 = _GEN_645 ? _GEN_5311 : dirty_0_49; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6210 = _GEN_645 ? _GEN_5312 : dirty_0_50; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6211 = _GEN_645 ? _GEN_5313 : dirty_0_51; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6212 = _GEN_645 ? _GEN_5314 : dirty_0_52; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6213 = _GEN_645 ? _GEN_5315 : dirty_0_53; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6214 = _GEN_645 ? _GEN_5316 : dirty_0_54; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6215 = _GEN_645 ? _GEN_5317 : dirty_0_55; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6216 = _GEN_645 ? _GEN_5318 : dirty_0_56; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6217 = _GEN_645 ? _GEN_5319 : dirty_0_57; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6218 = _GEN_645 ? _GEN_5320 : dirty_0_58; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6219 = _GEN_645 ? _GEN_5321 : dirty_0_59; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6220 = _GEN_645 ? _GEN_5322 : dirty_0_60; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6221 = _GEN_645 ? _GEN_5323 : dirty_0_61; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6222 = _GEN_645 ? _GEN_5324 : dirty_0_62; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6223 = _GEN_645 ? _GEN_5325 : dirty_0_63; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6224 = _GEN_645 ? _GEN_5326 : dirty_0_64; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6225 = _GEN_645 ? _GEN_5327 : dirty_0_65; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6226 = _GEN_645 ? _GEN_5328 : dirty_0_66; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6227 = _GEN_645 ? _GEN_5329 : dirty_0_67; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6228 = _GEN_645 ? _GEN_5330 : dirty_0_68; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6229 = _GEN_645 ? _GEN_5331 : dirty_0_69; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6230 = _GEN_645 ? _GEN_5332 : dirty_0_70; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6231 = _GEN_645 ? _GEN_5333 : dirty_0_71; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6232 = _GEN_645 ? _GEN_5334 : dirty_0_72; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6233 = _GEN_645 ? _GEN_5335 : dirty_0_73; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6234 = _GEN_645 ? _GEN_5336 : dirty_0_74; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6235 = _GEN_645 ? _GEN_5337 : dirty_0_75; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6236 = _GEN_645 ? _GEN_5338 : dirty_0_76; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6237 = _GEN_645 ? _GEN_5339 : dirty_0_77; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6238 = _GEN_645 ? _GEN_5340 : dirty_0_78; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6239 = _GEN_645 ? _GEN_5341 : dirty_0_79; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6240 = _GEN_645 ? _GEN_5342 : dirty_0_80; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6241 = _GEN_645 ? _GEN_5343 : dirty_0_81; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6242 = _GEN_645 ? _GEN_5344 : dirty_0_82; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6243 = _GEN_645 ? _GEN_5345 : dirty_0_83; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6244 = _GEN_645 ? _GEN_5346 : dirty_0_84; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6245 = _GEN_645 ? _GEN_5347 : dirty_0_85; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6246 = _GEN_645 ? _GEN_5348 : dirty_0_86; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6247 = _GEN_645 ? _GEN_5349 : dirty_0_87; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6248 = _GEN_645 ? _GEN_5350 : dirty_0_88; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6249 = _GEN_645 ? _GEN_5351 : dirty_0_89; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6250 = _GEN_645 ? _GEN_5352 : dirty_0_90; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6251 = _GEN_645 ? _GEN_5353 : dirty_0_91; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6252 = _GEN_645 ? _GEN_5354 : dirty_0_92; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6253 = _GEN_645 ? _GEN_5355 : dirty_0_93; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6254 = _GEN_645 ? _GEN_5356 : dirty_0_94; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6255 = _GEN_645 ? _GEN_5357 : dirty_0_95; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6256 = _GEN_645 ? _GEN_5358 : dirty_0_96; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6257 = _GEN_645 ? _GEN_5359 : dirty_0_97; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6258 = _GEN_645 ? _GEN_5360 : dirty_0_98; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6259 = _GEN_645 ? _GEN_5361 : dirty_0_99; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6260 = _GEN_645 ? _GEN_5362 : dirty_0_100; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6261 = _GEN_645 ? _GEN_5363 : dirty_0_101; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6262 = _GEN_645 ? _GEN_5364 : dirty_0_102; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6263 = _GEN_645 ? _GEN_5365 : dirty_0_103; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6264 = _GEN_645 ? _GEN_5366 : dirty_0_104; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6265 = _GEN_645 ? _GEN_5367 : dirty_0_105; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6266 = _GEN_645 ? _GEN_5368 : dirty_0_106; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6267 = _GEN_645 ? _GEN_5369 : dirty_0_107; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6268 = _GEN_645 ? _GEN_5370 : dirty_0_108; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6269 = _GEN_645 ? _GEN_5371 : dirty_0_109; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6270 = _GEN_645 ? _GEN_5372 : dirty_0_110; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6271 = _GEN_645 ? _GEN_5373 : dirty_0_111; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6272 = _GEN_645 ? _GEN_5374 : dirty_0_112; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6273 = _GEN_645 ? _GEN_5375 : dirty_0_113; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6274 = _GEN_645 ? _GEN_5376 : dirty_0_114; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6275 = _GEN_645 ? _GEN_5377 : dirty_0_115; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6276 = _GEN_645 ? _GEN_5378 : dirty_0_116; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6277 = _GEN_645 ? _GEN_5379 : dirty_0_117; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6278 = _GEN_645 ? _GEN_5380 : dirty_0_118; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6279 = _GEN_645 ? _GEN_5381 : dirty_0_119; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6280 = _GEN_645 ? _GEN_5382 : dirty_0_120; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6281 = _GEN_645 ? _GEN_5383 : dirty_0_121; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6282 = _GEN_645 ? _GEN_5384 : dirty_0_122; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6283 = _GEN_645 ? _GEN_5385 : dirty_0_123; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6284 = _GEN_645 ? _GEN_5386 : dirty_0_124; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6285 = _GEN_645 ? _GEN_5387 : dirty_0_125; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6286 = _GEN_645 ? _GEN_5388 : dirty_0_126; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6287 = _GEN_645 ? _GEN_5389 : dirty_0_127; // @[d_cache.scala 165:47 32:26]
  wire  _GEN_6288 = _GEN_645 ? _GEN_4494 : _GEN_4494; // @[d_cache.scala 165:47]
  wire  _GEN_6289 = _GEN_645 ? _GEN_4495 : _GEN_4495; // @[d_cache.scala 165:47]
  wire  _GEN_6290 = _GEN_645 ? _GEN_4496 : _GEN_4496; // @[d_cache.scala 165:47]
  wire  _GEN_6291 = _GEN_645 ? _GEN_4497 : _GEN_4497; // @[d_cache.scala 165:47]
  wire  _GEN_6292 = _GEN_645 ? _GEN_4498 : _GEN_4498; // @[d_cache.scala 165:47]
  wire  _GEN_6293 = _GEN_645 ? _GEN_4499 : _GEN_4499; // @[d_cache.scala 165:47]
  wire  _GEN_6294 = _GEN_645 ? _GEN_4500 : _GEN_4500; // @[d_cache.scala 165:47]
  wire  _GEN_6295 = _GEN_645 ? _GEN_4501 : _GEN_4501; // @[d_cache.scala 165:47]
  wire  _GEN_6296 = _GEN_645 ? _GEN_4502 : _GEN_4502; // @[d_cache.scala 165:47]
  wire  _GEN_6297 = _GEN_645 ? _GEN_4503 : _GEN_4503; // @[d_cache.scala 165:47]
  wire  _GEN_6298 = _GEN_645 ? _GEN_4504 : _GEN_4504; // @[d_cache.scala 165:47]
  wire  _GEN_6299 = _GEN_645 ? _GEN_4505 : _GEN_4505; // @[d_cache.scala 165:47]
  wire  _GEN_6300 = _GEN_645 ? _GEN_4506 : _GEN_4506; // @[d_cache.scala 165:47]
  wire  _GEN_6301 = _GEN_645 ? _GEN_4507 : _GEN_4507; // @[d_cache.scala 165:47]
  wire  _GEN_6302 = _GEN_645 ? _GEN_4508 : _GEN_4508; // @[d_cache.scala 165:47]
  wire  _GEN_6303 = _GEN_645 ? _GEN_4509 : _GEN_4509; // @[d_cache.scala 165:47]
  wire  _GEN_6304 = _GEN_645 ? _GEN_4510 : _GEN_4510; // @[d_cache.scala 165:47]
  wire  _GEN_6305 = _GEN_645 ? _GEN_4511 : _GEN_4511; // @[d_cache.scala 165:47]
  wire  _GEN_6306 = _GEN_645 ? _GEN_4512 : _GEN_4512; // @[d_cache.scala 165:47]
  wire  _GEN_6307 = _GEN_645 ? _GEN_4513 : _GEN_4513; // @[d_cache.scala 165:47]
  wire  _GEN_6308 = _GEN_645 ? _GEN_4514 : _GEN_4514; // @[d_cache.scala 165:47]
  wire  _GEN_6309 = _GEN_645 ? _GEN_4515 : _GEN_4515; // @[d_cache.scala 165:47]
  wire  _GEN_6310 = _GEN_645 ? _GEN_4516 : _GEN_4516; // @[d_cache.scala 165:47]
  wire  _GEN_6311 = _GEN_645 ? _GEN_4517 : _GEN_4517; // @[d_cache.scala 165:47]
  wire  _GEN_6312 = _GEN_645 ? _GEN_4518 : _GEN_4518; // @[d_cache.scala 165:47]
  wire  _GEN_6313 = _GEN_645 ? _GEN_4519 : _GEN_4519; // @[d_cache.scala 165:47]
  wire  _GEN_6314 = _GEN_645 ? _GEN_4520 : _GEN_4520; // @[d_cache.scala 165:47]
  wire  _GEN_6315 = _GEN_645 ? _GEN_4521 : _GEN_4521; // @[d_cache.scala 165:47]
  wire  _GEN_6316 = _GEN_645 ? _GEN_4522 : _GEN_4522; // @[d_cache.scala 165:47]
  wire  _GEN_6317 = _GEN_645 ? _GEN_4523 : _GEN_4523; // @[d_cache.scala 165:47]
  wire  _GEN_6318 = _GEN_645 ? _GEN_4524 : _GEN_4524; // @[d_cache.scala 165:47]
  wire  _GEN_6319 = _GEN_645 ? _GEN_4525 : _GEN_4525; // @[d_cache.scala 165:47]
  wire  _GEN_6320 = _GEN_645 ? _GEN_4526 : _GEN_4526; // @[d_cache.scala 165:47]
  wire  _GEN_6321 = _GEN_645 ? _GEN_4527 : _GEN_4527; // @[d_cache.scala 165:47]
  wire  _GEN_6322 = _GEN_645 ? _GEN_4528 : _GEN_4528; // @[d_cache.scala 165:47]
  wire  _GEN_6323 = _GEN_645 ? _GEN_4529 : _GEN_4529; // @[d_cache.scala 165:47]
  wire  _GEN_6324 = _GEN_645 ? _GEN_4530 : _GEN_4530; // @[d_cache.scala 165:47]
  wire  _GEN_6325 = _GEN_645 ? _GEN_4531 : _GEN_4531; // @[d_cache.scala 165:47]
  wire  _GEN_6326 = _GEN_645 ? _GEN_4532 : _GEN_4532; // @[d_cache.scala 165:47]
  wire  _GEN_6327 = _GEN_645 ? _GEN_4533 : _GEN_4533; // @[d_cache.scala 165:47]
  wire  _GEN_6328 = _GEN_645 ? _GEN_4534 : _GEN_4534; // @[d_cache.scala 165:47]
  wire  _GEN_6329 = _GEN_645 ? _GEN_4535 : _GEN_4535; // @[d_cache.scala 165:47]
  wire  _GEN_6330 = _GEN_645 ? _GEN_4536 : _GEN_4536; // @[d_cache.scala 165:47]
  wire  _GEN_6331 = _GEN_645 ? _GEN_4537 : _GEN_4537; // @[d_cache.scala 165:47]
  wire  _GEN_6332 = _GEN_645 ? _GEN_4538 : _GEN_4538; // @[d_cache.scala 165:47]
  wire  _GEN_6333 = _GEN_645 ? _GEN_4539 : _GEN_4539; // @[d_cache.scala 165:47]
  wire  _GEN_6334 = _GEN_645 ? _GEN_4540 : _GEN_4540; // @[d_cache.scala 165:47]
  wire  _GEN_6335 = _GEN_645 ? _GEN_4541 : _GEN_4541; // @[d_cache.scala 165:47]
  wire  _GEN_6336 = _GEN_645 ? _GEN_4542 : _GEN_4542; // @[d_cache.scala 165:47]
  wire  _GEN_6337 = _GEN_645 ? _GEN_4543 : _GEN_4543; // @[d_cache.scala 165:47]
  wire  _GEN_6338 = _GEN_645 ? _GEN_4544 : _GEN_4544; // @[d_cache.scala 165:47]
  wire  _GEN_6339 = _GEN_645 ? _GEN_4545 : _GEN_4545; // @[d_cache.scala 165:47]
  wire  _GEN_6340 = _GEN_645 ? _GEN_4546 : _GEN_4546; // @[d_cache.scala 165:47]
  wire  _GEN_6341 = _GEN_645 ? _GEN_4547 : _GEN_4547; // @[d_cache.scala 165:47]
  wire  _GEN_6342 = _GEN_645 ? _GEN_4548 : _GEN_4548; // @[d_cache.scala 165:47]
  wire  _GEN_6343 = _GEN_645 ? _GEN_4549 : _GEN_4549; // @[d_cache.scala 165:47]
  wire  _GEN_6344 = _GEN_645 ? _GEN_4550 : _GEN_4550; // @[d_cache.scala 165:47]
  wire  _GEN_6345 = _GEN_645 ? _GEN_4551 : _GEN_4551; // @[d_cache.scala 165:47]
  wire  _GEN_6346 = _GEN_645 ? _GEN_4552 : _GEN_4552; // @[d_cache.scala 165:47]
  wire  _GEN_6347 = _GEN_645 ? _GEN_4553 : _GEN_4553; // @[d_cache.scala 165:47]
  wire  _GEN_6348 = _GEN_645 ? _GEN_4554 : _GEN_4554; // @[d_cache.scala 165:47]
  wire  _GEN_6349 = _GEN_645 ? _GEN_4555 : _GEN_4555; // @[d_cache.scala 165:47]
  wire  _GEN_6350 = _GEN_645 ? _GEN_4556 : _GEN_4556; // @[d_cache.scala 165:47]
  wire  _GEN_6351 = _GEN_645 ? _GEN_4557 : _GEN_4557; // @[d_cache.scala 165:47]
  wire  _GEN_6352 = _GEN_645 ? _GEN_4558 : _GEN_4558; // @[d_cache.scala 165:47]
  wire  _GEN_6353 = _GEN_645 ? _GEN_4559 : _GEN_4559; // @[d_cache.scala 165:47]
  wire  _GEN_6354 = _GEN_645 ? _GEN_4560 : _GEN_4560; // @[d_cache.scala 165:47]
  wire  _GEN_6355 = _GEN_645 ? _GEN_4561 : _GEN_4561; // @[d_cache.scala 165:47]
  wire  _GEN_6356 = _GEN_645 ? _GEN_4562 : _GEN_4562; // @[d_cache.scala 165:47]
  wire  _GEN_6357 = _GEN_645 ? _GEN_4563 : _GEN_4563; // @[d_cache.scala 165:47]
  wire  _GEN_6358 = _GEN_645 ? _GEN_4564 : _GEN_4564; // @[d_cache.scala 165:47]
  wire  _GEN_6359 = _GEN_645 ? _GEN_4565 : _GEN_4565; // @[d_cache.scala 165:47]
  wire  _GEN_6360 = _GEN_645 ? _GEN_4566 : _GEN_4566; // @[d_cache.scala 165:47]
  wire  _GEN_6361 = _GEN_645 ? _GEN_4567 : _GEN_4567; // @[d_cache.scala 165:47]
  wire  _GEN_6362 = _GEN_645 ? _GEN_4568 : _GEN_4568; // @[d_cache.scala 165:47]
  wire  _GEN_6363 = _GEN_645 ? _GEN_4569 : _GEN_4569; // @[d_cache.scala 165:47]
  wire  _GEN_6364 = _GEN_645 ? _GEN_4570 : _GEN_4570; // @[d_cache.scala 165:47]
  wire  _GEN_6365 = _GEN_645 ? _GEN_4571 : _GEN_4571; // @[d_cache.scala 165:47]
  wire  _GEN_6366 = _GEN_645 ? _GEN_4572 : _GEN_4572; // @[d_cache.scala 165:47]
  wire  _GEN_6367 = _GEN_645 ? _GEN_4573 : _GEN_4573; // @[d_cache.scala 165:47]
  wire  _GEN_6368 = _GEN_645 ? _GEN_4574 : _GEN_4574; // @[d_cache.scala 165:47]
  wire  _GEN_6369 = _GEN_645 ? _GEN_4575 : _GEN_4575; // @[d_cache.scala 165:47]
  wire  _GEN_6370 = _GEN_645 ? _GEN_4576 : _GEN_4576; // @[d_cache.scala 165:47]
  wire  _GEN_6371 = _GEN_645 ? _GEN_4577 : _GEN_4577; // @[d_cache.scala 165:47]
  wire  _GEN_6372 = _GEN_645 ? _GEN_4578 : _GEN_4578; // @[d_cache.scala 165:47]
  wire  _GEN_6373 = _GEN_645 ? _GEN_4579 : _GEN_4579; // @[d_cache.scala 165:47]
  wire  _GEN_6374 = _GEN_645 ? _GEN_4580 : _GEN_4580; // @[d_cache.scala 165:47]
  wire  _GEN_6375 = _GEN_645 ? _GEN_4581 : _GEN_4581; // @[d_cache.scala 165:47]
  wire  _GEN_6376 = _GEN_645 ? _GEN_4582 : _GEN_4582; // @[d_cache.scala 165:47]
  wire  _GEN_6377 = _GEN_645 ? _GEN_4583 : _GEN_4583; // @[d_cache.scala 165:47]
  wire  _GEN_6378 = _GEN_645 ? _GEN_4584 : _GEN_4584; // @[d_cache.scala 165:47]
  wire  _GEN_6379 = _GEN_645 ? _GEN_4585 : _GEN_4585; // @[d_cache.scala 165:47]
  wire  _GEN_6380 = _GEN_645 ? _GEN_4586 : _GEN_4586; // @[d_cache.scala 165:47]
  wire  _GEN_6381 = _GEN_645 ? _GEN_4587 : _GEN_4587; // @[d_cache.scala 165:47]
  wire  _GEN_6382 = _GEN_645 ? _GEN_4588 : _GEN_4588; // @[d_cache.scala 165:47]
  wire  _GEN_6383 = _GEN_645 ? _GEN_4589 : _GEN_4589; // @[d_cache.scala 165:47]
  wire  _GEN_6384 = _GEN_645 ? _GEN_4590 : _GEN_4590; // @[d_cache.scala 165:47]
  wire  _GEN_6385 = _GEN_645 ? _GEN_4591 : _GEN_4591; // @[d_cache.scala 165:47]
  wire  _GEN_6386 = _GEN_645 ? _GEN_4592 : _GEN_4592; // @[d_cache.scala 165:47]
  wire  _GEN_6387 = _GEN_645 ? _GEN_4593 : _GEN_4593; // @[d_cache.scala 165:47]
  wire  _GEN_6388 = _GEN_645 ? _GEN_4594 : _GEN_4594; // @[d_cache.scala 165:47]
  wire  _GEN_6389 = _GEN_645 ? _GEN_4595 : _GEN_4595; // @[d_cache.scala 165:47]
  wire  _GEN_6390 = _GEN_645 ? _GEN_4596 : _GEN_4596; // @[d_cache.scala 165:47]
  wire  _GEN_6391 = _GEN_645 ? _GEN_4597 : _GEN_4597; // @[d_cache.scala 165:47]
  wire  _GEN_6392 = _GEN_645 ? _GEN_4598 : _GEN_4598; // @[d_cache.scala 165:47]
  wire  _GEN_6393 = _GEN_645 ? _GEN_4599 : _GEN_4599; // @[d_cache.scala 165:47]
  wire  _GEN_6394 = _GEN_645 ? _GEN_4600 : _GEN_4600; // @[d_cache.scala 165:47]
  wire  _GEN_6395 = _GEN_645 ? _GEN_4601 : _GEN_4601; // @[d_cache.scala 165:47]
  wire  _GEN_6396 = _GEN_645 ? _GEN_4602 : _GEN_4602; // @[d_cache.scala 165:47]
  wire  _GEN_6397 = _GEN_645 ? _GEN_4603 : _GEN_4603; // @[d_cache.scala 165:47]
  wire  _GEN_6398 = _GEN_645 ? _GEN_4604 : _GEN_4604; // @[d_cache.scala 165:47]
  wire  _GEN_6399 = _GEN_645 ? _GEN_4605 : _GEN_4605; // @[d_cache.scala 165:47]
  wire  _GEN_6400 = _GEN_645 ? _GEN_4606 : _GEN_4606; // @[d_cache.scala 165:47]
  wire  _GEN_6401 = _GEN_645 ? _GEN_4607 : _GEN_4607; // @[d_cache.scala 165:47]
  wire  _GEN_6402 = _GEN_645 ? _GEN_4608 : _GEN_4608; // @[d_cache.scala 165:47]
  wire  _GEN_6403 = _GEN_645 ? _GEN_4609 : _GEN_4609; // @[d_cache.scala 165:47]
  wire  _GEN_6404 = _GEN_645 ? _GEN_4610 : _GEN_4610; // @[d_cache.scala 165:47]
  wire  _GEN_6405 = _GEN_645 ? _GEN_4611 : _GEN_4611; // @[d_cache.scala 165:47]
  wire  _GEN_6406 = _GEN_645 ? _GEN_4612 : _GEN_4612; // @[d_cache.scala 165:47]
  wire  _GEN_6407 = _GEN_645 ? _GEN_4613 : _GEN_4613; // @[d_cache.scala 165:47]
  wire  _GEN_6408 = _GEN_645 ? _GEN_4614 : _GEN_4614; // @[d_cache.scala 165:47]
  wire  _GEN_6409 = _GEN_645 ? _GEN_4615 : _GEN_4615; // @[d_cache.scala 165:47]
  wire  _GEN_6410 = _GEN_645 ? _GEN_4616 : _GEN_4616; // @[d_cache.scala 165:47]
  wire  _GEN_6411 = _GEN_645 ? _GEN_4617 : _GEN_4617; // @[d_cache.scala 165:47]
  wire  _GEN_6412 = _GEN_645 ? _GEN_4618 : _GEN_4618; // @[d_cache.scala 165:47]
  wire  _GEN_6413 = _GEN_645 ? _GEN_4619 : _GEN_4619; // @[d_cache.scala 165:47]
  wire  _GEN_6414 = _GEN_645 ? _GEN_4620 : _GEN_4620; // @[d_cache.scala 165:47]
  wire  _GEN_6415 = _GEN_645 ? _GEN_4621 : _GEN_4621; // @[d_cache.scala 165:47]
  wire [2:0] _GEN_6416 = _GEN_645 ? 3'h6 : 3'h7; // @[d_cache.scala 165:47 172:31 175:31]
  wire [41:0] _write_back_addr_T_3 = {_GEN_384,index,3'h0}; // @[Cat.scala 31:58]
  wire  _GEN_6674 = 7'h0 == index ? 1'h0 : dirty_1_0; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6675 = 7'h1 == index ? 1'h0 : dirty_1_1; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6676 = 7'h2 == index ? 1'h0 : dirty_1_2; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6677 = 7'h3 == index ? 1'h0 : dirty_1_3; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6678 = 7'h4 == index ? 1'h0 : dirty_1_4; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6679 = 7'h5 == index ? 1'h0 : dirty_1_5; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6680 = 7'h6 == index ? 1'h0 : dirty_1_6; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6681 = 7'h7 == index ? 1'h0 : dirty_1_7; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6682 = 7'h8 == index ? 1'h0 : dirty_1_8; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6683 = 7'h9 == index ? 1'h0 : dirty_1_9; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6684 = 7'ha == index ? 1'h0 : dirty_1_10; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6685 = 7'hb == index ? 1'h0 : dirty_1_11; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6686 = 7'hc == index ? 1'h0 : dirty_1_12; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6687 = 7'hd == index ? 1'h0 : dirty_1_13; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6688 = 7'he == index ? 1'h0 : dirty_1_14; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6689 = 7'hf == index ? 1'h0 : dirty_1_15; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6690 = 7'h10 == index ? 1'h0 : dirty_1_16; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6691 = 7'h11 == index ? 1'h0 : dirty_1_17; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6692 = 7'h12 == index ? 1'h0 : dirty_1_18; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6693 = 7'h13 == index ? 1'h0 : dirty_1_19; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6694 = 7'h14 == index ? 1'h0 : dirty_1_20; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6695 = 7'h15 == index ? 1'h0 : dirty_1_21; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6696 = 7'h16 == index ? 1'h0 : dirty_1_22; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6697 = 7'h17 == index ? 1'h0 : dirty_1_23; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6698 = 7'h18 == index ? 1'h0 : dirty_1_24; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6699 = 7'h19 == index ? 1'h0 : dirty_1_25; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6700 = 7'h1a == index ? 1'h0 : dirty_1_26; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6701 = 7'h1b == index ? 1'h0 : dirty_1_27; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6702 = 7'h1c == index ? 1'h0 : dirty_1_28; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6703 = 7'h1d == index ? 1'h0 : dirty_1_29; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6704 = 7'h1e == index ? 1'h0 : dirty_1_30; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6705 = 7'h1f == index ? 1'h0 : dirty_1_31; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6706 = 7'h20 == index ? 1'h0 : dirty_1_32; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6707 = 7'h21 == index ? 1'h0 : dirty_1_33; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6708 = 7'h22 == index ? 1'h0 : dirty_1_34; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6709 = 7'h23 == index ? 1'h0 : dirty_1_35; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6710 = 7'h24 == index ? 1'h0 : dirty_1_36; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6711 = 7'h25 == index ? 1'h0 : dirty_1_37; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6712 = 7'h26 == index ? 1'h0 : dirty_1_38; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6713 = 7'h27 == index ? 1'h0 : dirty_1_39; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6714 = 7'h28 == index ? 1'h0 : dirty_1_40; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6715 = 7'h29 == index ? 1'h0 : dirty_1_41; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6716 = 7'h2a == index ? 1'h0 : dirty_1_42; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6717 = 7'h2b == index ? 1'h0 : dirty_1_43; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6718 = 7'h2c == index ? 1'h0 : dirty_1_44; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6719 = 7'h2d == index ? 1'h0 : dirty_1_45; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6720 = 7'h2e == index ? 1'h0 : dirty_1_46; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6721 = 7'h2f == index ? 1'h0 : dirty_1_47; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6722 = 7'h30 == index ? 1'h0 : dirty_1_48; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6723 = 7'h31 == index ? 1'h0 : dirty_1_49; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6724 = 7'h32 == index ? 1'h0 : dirty_1_50; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6725 = 7'h33 == index ? 1'h0 : dirty_1_51; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6726 = 7'h34 == index ? 1'h0 : dirty_1_52; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6727 = 7'h35 == index ? 1'h0 : dirty_1_53; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6728 = 7'h36 == index ? 1'h0 : dirty_1_54; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6729 = 7'h37 == index ? 1'h0 : dirty_1_55; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6730 = 7'h38 == index ? 1'h0 : dirty_1_56; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6731 = 7'h39 == index ? 1'h0 : dirty_1_57; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6732 = 7'h3a == index ? 1'h0 : dirty_1_58; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6733 = 7'h3b == index ? 1'h0 : dirty_1_59; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6734 = 7'h3c == index ? 1'h0 : dirty_1_60; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6735 = 7'h3d == index ? 1'h0 : dirty_1_61; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6736 = 7'h3e == index ? 1'h0 : dirty_1_62; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6737 = 7'h3f == index ? 1'h0 : dirty_1_63; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6738 = 7'h40 == index ? 1'h0 : dirty_1_64; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6739 = 7'h41 == index ? 1'h0 : dirty_1_65; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6740 = 7'h42 == index ? 1'h0 : dirty_1_66; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6741 = 7'h43 == index ? 1'h0 : dirty_1_67; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6742 = 7'h44 == index ? 1'h0 : dirty_1_68; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6743 = 7'h45 == index ? 1'h0 : dirty_1_69; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6744 = 7'h46 == index ? 1'h0 : dirty_1_70; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6745 = 7'h47 == index ? 1'h0 : dirty_1_71; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6746 = 7'h48 == index ? 1'h0 : dirty_1_72; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6747 = 7'h49 == index ? 1'h0 : dirty_1_73; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6748 = 7'h4a == index ? 1'h0 : dirty_1_74; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6749 = 7'h4b == index ? 1'h0 : dirty_1_75; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6750 = 7'h4c == index ? 1'h0 : dirty_1_76; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6751 = 7'h4d == index ? 1'h0 : dirty_1_77; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6752 = 7'h4e == index ? 1'h0 : dirty_1_78; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6753 = 7'h4f == index ? 1'h0 : dirty_1_79; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6754 = 7'h50 == index ? 1'h0 : dirty_1_80; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6755 = 7'h51 == index ? 1'h0 : dirty_1_81; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6756 = 7'h52 == index ? 1'h0 : dirty_1_82; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6757 = 7'h53 == index ? 1'h0 : dirty_1_83; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6758 = 7'h54 == index ? 1'h0 : dirty_1_84; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6759 = 7'h55 == index ? 1'h0 : dirty_1_85; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6760 = 7'h56 == index ? 1'h0 : dirty_1_86; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6761 = 7'h57 == index ? 1'h0 : dirty_1_87; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6762 = 7'h58 == index ? 1'h0 : dirty_1_88; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6763 = 7'h59 == index ? 1'h0 : dirty_1_89; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6764 = 7'h5a == index ? 1'h0 : dirty_1_90; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6765 = 7'h5b == index ? 1'h0 : dirty_1_91; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6766 = 7'h5c == index ? 1'h0 : dirty_1_92; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6767 = 7'h5d == index ? 1'h0 : dirty_1_93; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6768 = 7'h5e == index ? 1'h0 : dirty_1_94; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6769 = 7'h5f == index ? 1'h0 : dirty_1_95; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6770 = 7'h60 == index ? 1'h0 : dirty_1_96; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6771 = 7'h61 == index ? 1'h0 : dirty_1_97; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6772 = 7'h62 == index ? 1'h0 : dirty_1_98; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6773 = 7'h63 == index ? 1'h0 : dirty_1_99; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6774 = 7'h64 == index ? 1'h0 : dirty_1_100; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6775 = 7'h65 == index ? 1'h0 : dirty_1_101; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6776 = 7'h66 == index ? 1'h0 : dirty_1_102; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6777 = 7'h67 == index ? 1'h0 : dirty_1_103; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6778 = 7'h68 == index ? 1'h0 : dirty_1_104; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6779 = 7'h69 == index ? 1'h0 : dirty_1_105; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6780 = 7'h6a == index ? 1'h0 : dirty_1_106; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6781 = 7'h6b == index ? 1'h0 : dirty_1_107; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6782 = 7'h6c == index ? 1'h0 : dirty_1_108; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6783 = 7'h6d == index ? 1'h0 : dirty_1_109; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6784 = 7'h6e == index ? 1'h0 : dirty_1_110; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6785 = 7'h6f == index ? 1'h0 : dirty_1_111; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6786 = 7'h70 == index ? 1'h0 : dirty_1_112; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6787 = 7'h71 == index ? 1'h0 : dirty_1_113; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6788 = 7'h72 == index ? 1'h0 : dirty_1_114; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6789 = 7'h73 == index ? 1'h0 : dirty_1_115; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6790 = 7'h74 == index ? 1'h0 : dirty_1_116; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6791 = 7'h75 == index ? 1'h0 : dirty_1_117; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6792 = 7'h76 == index ? 1'h0 : dirty_1_118; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6793 = 7'h77 == index ? 1'h0 : dirty_1_119; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6794 = 7'h78 == index ? 1'h0 : dirty_1_120; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6795 = 7'h79 == index ? 1'h0 : dirty_1_121; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6796 = 7'h7a == index ? 1'h0 : dirty_1_122; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6797 = 7'h7b == index ? 1'h0 : dirty_1_123; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6798 = 7'h7c == index ? 1'h0 : dirty_1_124; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6799 = 7'h7d == index ? 1'h0 : dirty_1_125; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6800 = 7'h7e == index ? 1'h0 : dirty_1_126; // @[d_cache.scala 187:{40,40} 33:26]
  wire  _GEN_6801 = 7'h7f == index ? 1'h0 : dirty_1_127; // @[d_cache.scala 187:{40,40} 33:26]
  wire [63:0] _GEN_7314 = _GEN_774 ? _GEN_1416 : write_back_data; // @[d_cache.scala 182:47 183:41 37:34]
  wire [41:0] _GEN_7315 = _GEN_774 ? _write_back_addr_T_3 : {{10'd0}, write_back_addr}; // @[d_cache.scala 182:47 184:41 38:34]
  wire [63:0] _GEN_7316 = _GEN_774 ? _GEN_4622 : _GEN_4622; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7317 = _GEN_774 ? _GEN_4623 : _GEN_4623; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7318 = _GEN_774 ? _GEN_4624 : _GEN_4624; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7319 = _GEN_774 ? _GEN_4625 : _GEN_4625; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7320 = _GEN_774 ? _GEN_4626 : _GEN_4626; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7321 = _GEN_774 ? _GEN_4627 : _GEN_4627; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7322 = _GEN_774 ? _GEN_4628 : _GEN_4628; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7323 = _GEN_774 ? _GEN_4629 : _GEN_4629; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7324 = _GEN_774 ? _GEN_4630 : _GEN_4630; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7325 = _GEN_774 ? _GEN_4631 : _GEN_4631; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7326 = _GEN_774 ? _GEN_4632 : _GEN_4632; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7327 = _GEN_774 ? _GEN_4633 : _GEN_4633; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7328 = _GEN_774 ? _GEN_4634 : _GEN_4634; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7329 = _GEN_774 ? _GEN_4635 : _GEN_4635; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7330 = _GEN_774 ? _GEN_4636 : _GEN_4636; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7331 = _GEN_774 ? _GEN_4637 : _GEN_4637; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7332 = _GEN_774 ? _GEN_4638 : _GEN_4638; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7333 = _GEN_774 ? _GEN_4639 : _GEN_4639; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7334 = _GEN_774 ? _GEN_4640 : _GEN_4640; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7335 = _GEN_774 ? _GEN_4641 : _GEN_4641; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7336 = _GEN_774 ? _GEN_4642 : _GEN_4642; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7337 = _GEN_774 ? _GEN_4643 : _GEN_4643; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7338 = _GEN_774 ? _GEN_4644 : _GEN_4644; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7339 = _GEN_774 ? _GEN_4645 : _GEN_4645; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7340 = _GEN_774 ? _GEN_4646 : _GEN_4646; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7341 = _GEN_774 ? _GEN_4647 : _GEN_4647; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7342 = _GEN_774 ? _GEN_4648 : _GEN_4648; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7343 = _GEN_774 ? _GEN_4649 : _GEN_4649; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7344 = _GEN_774 ? _GEN_4650 : _GEN_4650; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7345 = _GEN_774 ? _GEN_4651 : _GEN_4651; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7346 = _GEN_774 ? _GEN_4652 : _GEN_4652; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7347 = _GEN_774 ? _GEN_4653 : _GEN_4653; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7348 = _GEN_774 ? _GEN_4654 : _GEN_4654; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7349 = _GEN_774 ? _GEN_4655 : _GEN_4655; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7350 = _GEN_774 ? _GEN_4656 : _GEN_4656; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7351 = _GEN_774 ? _GEN_4657 : _GEN_4657; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7352 = _GEN_774 ? _GEN_4658 : _GEN_4658; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7353 = _GEN_774 ? _GEN_4659 : _GEN_4659; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7354 = _GEN_774 ? _GEN_4660 : _GEN_4660; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7355 = _GEN_774 ? _GEN_4661 : _GEN_4661; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7356 = _GEN_774 ? _GEN_4662 : _GEN_4662; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7357 = _GEN_774 ? _GEN_4663 : _GEN_4663; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7358 = _GEN_774 ? _GEN_4664 : _GEN_4664; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7359 = _GEN_774 ? _GEN_4665 : _GEN_4665; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7360 = _GEN_774 ? _GEN_4666 : _GEN_4666; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7361 = _GEN_774 ? _GEN_4667 : _GEN_4667; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7362 = _GEN_774 ? _GEN_4668 : _GEN_4668; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7363 = _GEN_774 ? _GEN_4669 : _GEN_4669; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7364 = _GEN_774 ? _GEN_4670 : _GEN_4670; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7365 = _GEN_774 ? _GEN_4671 : _GEN_4671; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7366 = _GEN_774 ? _GEN_4672 : _GEN_4672; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7367 = _GEN_774 ? _GEN_4673 : _GEN_4673; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7368 = _GEN_774 ? _GEN_4674 : _GEN_4674; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7369 = _GEN_774 ? _GEN_4675 : _GEN_4675; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7370 = _GEN_774 ? _GEN_4676 : _GEN_4676; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7371 = _GEN_774 ? _GEN_4677 : _GEN_4677; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7372 = _GEN_774 ? _GEN_4678 : _GEN_4678; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7373 = _GEN_774 ? _GEN_4679 : _GEN_4679; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7374 = _GEN_774 ? _GEN_4680 : _GEN_4680; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7375 = _GEN_774 ? _GEN_4681 : _GEN_4681; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7376 = _GEN_774 ? _GEN_4682 : _GEN_4682; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7377 = _GEN_774 ? _GEN_4683 : _GEN_4683; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7378 = _GEN_774 ? _GEN_4684 : _GEN_4684; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7379 = _GEN_774 ? _GEN_4685 : _GEN_4685; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7380 = _GEN_774 ? _GEN_4686 : _GEN_4686; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7381 = _GEN_774 ? _GEN_4687 : _GEN_4687; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7382 = _GEN_774 ? _GEN_4688 : _GEN_4688; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7383 = _GEN_774 ? _GEN_4689 : _GEN_4689; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7384 = _GEN_774 ? _GEN_4690 : _GEN_4690; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7385 = _GEN_774 ? _GEN_4691 : _GEN_4691; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7386 = _GEN_774 ? _GEN_4692 : _GEN_4692; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7387 = _GEN_774 ? _GEN_4693 : _GEN_4693; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7388 = _GEN_774 ? _GEN_4694 : _GEN_4694; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7389 = _GEN_774 ? _GEN_4695 : _GEN_4695; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7390 = _GEN_774 ? _GEN_4696 : _GEN_4696; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7391 = _GEN_774 ? _GEN_4697 : _GEN_4697; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7392 = _GEN_774 ? _GEN_4698 : _GEN_4698; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7393 = _GEN_774 ? _GEN_4699 : _GEN_4699; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7394 = _GEN_774 ? _GEN_4700 : _GEN_4700; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7395 = _GEN_774 ? _GEN_4701 : _GEN_4701; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7396 = _GEN_774 ? _GEN_4702 : _GEN_4702; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7397 = _GEN_774 ? _GEN_4703 : _GEN_4703; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7398 = _GEN_774 ? _GEN_4704 : _GEN_4704; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7399 = _GEN_774 ? _GEN_4705 : _GEN_4705; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7400 = _GEN_774 ? _GEN_4706 : _GEN_4706; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7401 = _GEN_774 ? _GEN_4707 : _GEN_4707; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7402 = _GEN_774 ? _GEN_4708 : _GEN_4708; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7403 = _GEN_774 ? _GEN_4709 : _GEN_4709; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7404 = _GEN_774 ? _GEN_4710 : _GEN_4710; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7405 = _GEN_774 ? _GEN_4711 : _GEN_4711; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7406 = _GEN_774 ? _GEN_4712 : _GEN_4712; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7407 = _GEN_774 ? _GEN_4713 : _GEN_4713; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7408 = _GEN_774 ? _GEN_4714 : _GEN_4714; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7409 = _GEN_774 ? _GEN_4715 : _GEN_4715; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7410 = _GEN_774 ? _GEN_4716 : _GEN_4716; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7411 = _GEN_774 ? _GEN_4717 : _GEN_4717; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7412 = _GEN_774 ? _GEN_4718 : _GEN_4718; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7413 = _GEN_774 ? _GEN_4719 : _GEN_4719; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7414 = _GEN_774 ? _GEN_4720 : _GEN_4720; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7415 = _GEN_774 ? _GEN_4721 : _GEN_4721; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7416 = _GEN_774 ? _GEN_4722 : _GEN_4722; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7417 = _GEN_774 ? _GEN_4723 : _GEN_4723; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7418 = _GEN_774 ? _GEN_4724 : _GEN_4724; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7419 = _GEN_774 ? _GEN_4725 : _GEN_4725; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7420 = _GEN_774 ? _GEN_4726 : _GEN_4726; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7421 = _GEN_774 ? _GEN_4727 : _GEN_4727; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7422 = _GEN_774 ? _GEN_4728 : _GEN_4728; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7423 = _GEN_774 ? _GEN_4729 : _GEN_4729; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7424 = _GEN_774 ? _GEN_4730 : _GEN_4730; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7425 = _GEN_774 ? _GEN_4731 : _GEN_4731; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7426 = _GEN_774 ? _GEN_4732 : _GEN_4732; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7427 = _GEN_774 ? _GEN_4733 : _GEN_4733; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7428 = _GEN_774 ? _GEN_4734 : _GEN_4734; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7429 = _GEN_774 ? _GEN_4735 : _GEN_4735; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7430 = _GEN_774 ? _GEN_4736 : _GEN_4736; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7431 = _GEN_774 ? _GEN_4737 : _GEN_4737; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7432 = _GEN_774 ? _GEN_4738 : _GEN_4738; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7433 = _GEN_774 ? _GEN_4739 : _GEN_4739; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7434 = _GEN_774 ? _GEN_4740 : _GEN_4740; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7435 = _GEN_774 ? _GEN_4741 : _GEN_4741; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7436 = _GEN_774 ? _GEN_4742 : _GEN_4742; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7437 = _GEN_774 ? _GEN_4743 : _GEN_4743; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7438 = _GEN_774 ? _GEN_4744 : _GEN_4744; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7439 = _GEN_774 ? _GEN_4745 : _GEN_4745; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7440 = _GEN_774 ? _GEN_4746 : _GEN_4746; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7441 = _GEN_774 ? _GEN_4747 : _GEN_4747; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7442 = _GEN_774 ? _GEN_4748 : _GEN_4748; // @[d_cache.scala 182:47]
  wire [63:0] _GEN_7443 = _GEN_774 ? _GEN_4749 : _GEN_4749; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7444 = _GEN_774 ? _GEN_4750 : _GEN_4750; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7445 = _GEN_774 ? _GEN_4751 : _GEN_4751; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7446 = _GEN_774 ? _GEN_4752 : _GEN_4752; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7447 = _GEN_774 ? _GEN_4753 : _GEN_4753; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7448 = _GEN_774 ? _GEN_4754 : _GEN_4754; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7449 = _GEN_774 ? _GEN_4755 : _GEN_4755; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7450 = _GEN_774 ? _GEN_4756 : _GEN_4756; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7451 = _GEN_774 ? _GEN_4757 : _GEN_4757; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7452 = _GEN_774 ? _GEN_4758 : _GEN_4758; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7453 = _GEN_774 ? _GEN_4759 : _GEN_4759; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7454 = _GEN_774 ? _GEN_4760 : _GEN_4760; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7455 = _GEN_774 ? _GEN_4761 : _GEN_4761; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7456 = _GEN_774 ? _GEN_4762 : _GEN_4762; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7457 = _GEN_774 ? _GEN_4763 : _GEN_4763; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7458 = _GEN_774 ? _GEN_4764 : _GEN_4764; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7459 = _GEN_774 ? _GEN_4765 : _GEN_4765; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7460 = _GEN_774 ? _GEN_4766 : _GEN_4766; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7461 = _GEN_774 ? _GEN_4767 : _GEN_4767; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7462 = _GEN_774 ? _GEN_4768 : _GEN_4768; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7463 = _GEN_774 ? _GEN_4769 : _GEN_4769; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7464 = _GEN_774 ? _GEN_4770 : _GEN_4770; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7465 = _GEN_774 ? _GEN_4771 : _GEN_4771; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7466 = _GEN_774 ? _GEN_4772 : _GEN_4772; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7467 = _GEN_774 ? _GEN_4773 : _GEN_4773; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7468 = _GEN_774 ? _GEN_4774 : _GEN_4774; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7469 = _GEN_774 ? _GEN_4775 : _GEN_4775; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7470 = _GEN_774 ? _GEN_4776 : _GEN_4776; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7471 = _GEN_774 ? _GEN_4777 : _GEN_4777; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7472 = _GEN_774 ? _GEN_4778 : _GEN_4778; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7473 = _GEN_774 ? _GEN_4779 : _GEN_4779; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7474 = _GEN_774 ? _GEN_4780 : _GEN_4780; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7475 = _GEN_774 ? _GEN_4781 : _GEN_4781; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7476 = _GEN_774 ? _GEN_4782 : _GEN_4782; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7477 = _GEN_774 ? _GEN_4783 : _GEN_4783; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7478 = _GEN_774 ? _GEN_4784 : _GEN_4784; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7479 = _GEN_774 ? _GEN_4785 : _GEN_4785; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7480 = _GEN_774 ? _GEN_4786 : _GEN_4786; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7481 = _GEN_774 ? _GEN_4787 : _GEN_4787; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7482 = _GEN_774 ? _GEN_4788 : _GEN_4788; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7483 = _GEN_774 ? _GEN_4789 : _GEN_4789; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7484 = _GEN_774 ? _GEN_4790 : _GEN_4790; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7485 = _GEN_774 ? _GEN_4791 : _GEN_4791; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7486 = _GEN_774 ? _GEN_4792 : _GEN_4792; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7487 = _GEN_774 ? _GEN_4793 : _GEN_4793; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7488 = _GEN_774 ? _GEN_4794 : _GEN_4794; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7489 = _GEN_774 ? _GEN_4795 : _GEN_4795; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7490 = _GEN_774 ? _GEN_4796 : _GEN_4796; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7491 = _GEN_774 ? _GEN_4797 : _GEN_4797; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7492 = _GEN_774 ? _GEN_4798 : _GEN_4798; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7493 = _GEN_774 ? _GEN_4799 : _GEN_4799; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7494 = _GEN_774 ? _GEN_4800 : _GEN_4800; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7495 = _GEN_774 ? _GEN_4801 : _GEN_4801; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7496 = _GEN_774 ? _GEN_4802 : _GEN_4802; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7497 = _GEN_774 ? _GEN_4803 : _GEN_4803; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7498 = _GEN_774 ? _GEN_4804 : _GEN_4804; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7499 = _GEN_774 ? _GEN_4805 : _GEN_4805; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7500 = _GEN_774 ? _GEN_4806 : _GEN_4806; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7501 = _GEN_774 ? _GEN_4807 : _GEN_4807; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7502 = _GEN_774 ? _GEN_4808 : _GEN_4808; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7503 = _GEN_774 ? _GEN_4809 : _GEN_4809; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7504 = _GEN_774 ? _GEN_4810 : _GEN_4810; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7505 = _GEN_774 ? _GEN_4811 : _GEN_4811; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7506 = _GEN_774 ? _GEN_4812 : _GEN_4812; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7507 = _GEN_774 ? _GEN_4813 : _GEN_4813; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7508 = _GEN_774 ? _GEN_4814 : _GEN_4814; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7509 = _GEN_774 ? _GEN_4815 : _GEN_4815; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7510 = _GEN_774 ? _GEN_4816 : _GEN_4816; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7511 = _GEN_774 ? _GEN_4817 : _GEN_4817; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7512 = _GEN_774 ? _GEN_4818 : _GEN_4818; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7513 = _GEN_774 ? _GEN_4819 : _GEN_4819; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7514 = _GEN_774 ? _GEN_4820 : _GEN_4820; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7515 = _GEN_774 ? _GEN_4821 : _GEN_4821; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7516 = _GEN_774 ? _GEN_4822 : _GEN_4822; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7517 = _GEN_774 ? _GEN_4823 : _GEN_4823; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7518 = _GEN_774 ? _GEN_4824 : _GEN_4824; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7519 = _GEN_774 ? _GEN_4825 : _GEN_4825; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7520 = _GEN_774 ? _GEN_4826 : _GEN_4826; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7521 = _GEN_774 ? _GEN_4827 : _GEN_4827; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7522 = _GEN_774 ? _GEN_4828 : _GEN_4828; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7523 = _GEN_774 ? _GEN_4829 : _GEN_4829; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7524 = _GEN_774 ? _GEN_4830 : _GEN_4830; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7525 = _GEN_774 ? _GEN_4831 : _GEN_4831; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7526 = _GEN_774 ? _GEN_4832 : _GEN_4832; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7527 = _GEN_774 ? _GEN_4833 : _GEN_4833; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7528 = _GEN_774 ? _GEN_4834 : _GEN_4834; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7529 = _GEN_774 ? _GEN_4835 : _GEN_4835; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7530 = _GEN_774 ? _GEN_4836 : _GEN_4836; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7531 = _GEN_774 ? _GEN_4837 : _GEN_4837; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7532 = _GEN_774 ? _GEN_4838 : _GEN_4838; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7533 = _GEN_774 ? _GEN_4839 : _GEN_4839; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7534 = _GEN_774 ? _GEN_4840 : _GEN_4840; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7535 = _GEN_774 ? _GEN_4841 : _GEN_4841; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7536 = _GEN_774 ? _GEN_4842 : _GEN_4842; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7537 = _GEN_774 ? _GEN_4843 : _GEN_4843; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7538 = _GEN_774 ? _GEN_4844 : _GEN_4844; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7539 = _GEN_774 ? _GEN_4845 : _GEN_4845; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7540 = _GEN_774 ? _GEN_4846 : _GEN_4846; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7541 = _GEN_774 ? _GEN_4847 : _GEN_4847; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7542 = _GEN_774 ? _GEN_4848 : _GEN_4848; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7543 = _GEN_774 ? _GEN_4849 : _GEN_4849; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7544 = _GEN_774 ? _GEN_4850 : _GEN_4850; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7545 = _GEN_774 ? _GEN_4851 : _GEN_4851; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7546 = _GEN_774 ? _GEN_4852 : _GEN_4852; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7547 = _GEN_774 ? _GEN_4853 : _GEN_4853; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7548 = _GEN_774 ? _GEN_4854 : _GEN_4854; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7549 = _GEN_774 ? _GEN_4855 : _GEN_4855; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7550 = _GEN_774 ? _GEN_4856 : _GEN_4856; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7551 = _GEN_774 ? _GEN_4857 : _GEN_4857; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7552 = _GEN_774 ? _GEN_4858 : _GEN_4858; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7553 = _GEN_774 ? _GEN_4859 : _GEN_4859; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7554 = _GEN_774 ? _GEN_4860 : _GEN_4860; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7555 = _GEN_774 ? _GEN_4861 : _GEN_4861; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7556 = _GEN_774 ? _GEN_4862 : _GEN_4862; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7557 = _GEN_774 ? _GEN_4863 : _GEN_4863; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7558 = _GEN_774 ? _GEN_4864 : _GEN_4864; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7559 = _GEN_774 ? _GEN_4865 : _GEN_4865; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7560 = _GEN_774 ? _GEN_4866 : _GEN_4866; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7561 = _GEN_774 ? _GEN_4867 : _GEN_4867; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7562 = _GEN_774 ? _GEN_4868 : _GEN_4868; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7563 = _GEN_774 ? _GEN_4869 : _GEN_4869; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7564 = _GEN_774 ? _GEN_4870 : _GEN_4870; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7565 = _GEN_774 ? _GEN_4871 : _GEN_4871; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7566 = _GEN_774 ? _GEN_4872 : _GEN_4872; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7567 = _GEN_774 ? _GEN_4873 : _GEN_4873; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7568 = _GEN_774 ? _GEN_4874 : _GEN_4874; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7569 = _GEN_774 ? _GEN_4875 : _GEN_4875; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7570 = _GEN_774 ? _GEN_4876 : _GEN_4876; // @[d_cache.scala 182:47]
  wire [31:0] _GEN_7571 = _GEN_774 ? _GEN_4877 : _GEN_4877; // @[d_cache.scala 182:47]
  wire  _GEN_7572 = _GEN_774 ? _GEN_6674 : dirty_1_0; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7573 = _GEN_774 ? _GEN_6675 : dirty_1_1; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7574 = _GEN_774 ? _GEN_6676 : dirty_1_2; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7575 = _GEN_774 ? _GEN_6677 : dirty_1_3; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7576 = _GEN_774 ? _GEN_6678 : dirty_1_4; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7577 = _GEN_774 ? _GEN_6679 : dirty_1_5; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7578 = _GEN_774 ? _GEN_6680 : dirty_1_6; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7579 = _GEN_774 ? _GEN_6681 : dirty_1_7; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7580 = _GEN_774 ? _GEN_6682 : dirty_1_8; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7581 = _GEN_774 ? _GEN_6683 : dirty_1_9; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7582 = _GEN_774 ? _GEN_6684 : dirty_1_10; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7583 = _GEN_774 ? _GEN_6685 : dirty_1_11; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7584 = _GEN_774 ? _GEN_6686 : dirty_1_12; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7585 = _GEN_774 ? _GEN_6687 : dirty_1_13; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7586 = _GEN_774 ? _GEN_6688 : dirty_1_14; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7587 = _GEN_774 ? _GEN_6689 : dirty_1_15; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7588 = _GEN_774 ? _GEN_6690 : dirty_1_16; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7589 = _GEN_774 ? _GEN_6691 : dirty_1_17; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7590 = _GEN_774 ? _GEN_6692 : dirty_1_18; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7591 = _GEN_774 ? _GEN_6693 : dirty_1_19; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7592 = _GEN_774 ? _GEN_6694 : dirty_1_20; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7593 = _GEN_774 ? _GEN_6695 : dirty_1_21; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7594 = _GEN_774 ? _GEN_6696 : dirty_1_22; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7595 = _GEN_774 ? _GEN_6697 : dirty_1_23; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7596 = _GEN_774 ? _GEN_6698 : dirty_1_24; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7597 = _GEN_774 ? _GEN_6699 : dirty_1_25; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7598 = _GEN_774 ? _GEN_6700 : dirty_1_26; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7599 = _GEN_774 ? _GEN_6701 : dirty_1_27; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7600 = _GEN_774 ? _GEN_6702 : dirty_1_28; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7601 = _GEN_774 ? _GEN_6703 : dirty_1_29; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7602 = _GEN_774 ? _GEN_6704 : dirty_1_30; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7603 = _GEN_774 ? _GEN_6705 : dirty_1_31; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7604 = _GEN_774 ? _GEN_6706 : dirty_1_32; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7605 = _GEN_774 ? _GEN_6707 : dirty_1_33; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7606 = _GEN_774 ? _GEN_6708 : dirty_1_34; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7607 = _GEN_774 ? _GEN_6709 : dirty_1_35; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7608 = _GEN_774 ? _GEN_6710 : dirty_1_36; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7609 = _GEN_774 ? _GEN_6711 : dirty_1_37; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7610 = _GEN_774 ? _GEN_6712 : dirty_1_38; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7611 = _GEN_774 ? _GEN_6713 : dirty_1_39; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7612 = _GEN_774 ? _GEN_6714 : dirty_1_40; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7613 = _GEN_774 ? _GEN_6715 : dirty_1_41; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7614 = _GEN_774 ? _GEN_6716 : dirty_1_42; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7615 = _GEN_774 ? _GEN_6717 : dirty_1_43; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7616 = _GEN_774 ? _GEN_6718 : dirty_1_44; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7617 = _GEN_774 ? _GEN_6719 : dirty_1_45; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7618 = _GEN_774 ? _GEN_6720 : dirty_1_46; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7619 = _GEN_774 ? _GEN_6721 : dirty_1_47; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7620 = _GEN_774 ? _GEN_6722 : dirty_1_48; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7621 = _GEN_774 ? _GEN_6723 : dirty_1_49; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7622 = _GEN_774 ? _GEN_6724 : dirty_1_50; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7623 = _GEN_774 ? _GEN_6725 : dirty_1_51; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7624 = _GEN_774 ? _GEN_6726 : dirty_1_52; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7625 = _GEN_774 ? _GEN_6727 : dirty_1_53; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7626 = _GEN_774 ? _GEN_6728 : dirty_1_54; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7627 = _GEN_774 ? _GEN_6729 : dirty_1_55; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7628 = _GEN_774 ? _GEN_6730 : dirty_1_56; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7629 = _GEN_774 ? _GEN_6731 : dirty_1_57; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7630 = _GEN_774 ? _GEN_6732 : dirty_1_58; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7631 = _GEN_774 ? _GEN_6733 : dirty_1_59; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7632 = _GEN_774 ? _GEN_6734 : dirty_1_60; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7633 = _GEN_774 ? _GEN_6735 : dirty_1_61; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7634 = _GEN_774 ? _GEN_6736 : dirty_1_62; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7635 = _GEN_774 ? _GEN_6737 : dirty_1_63; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7636 = _GEN_774 ? _GEN_6738 : dirty_1_64; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7637 = _GEN_774 ? _GEN_6739 : dirty_1_65; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7638 = _GEN_774 ? _GEN_6740 : dirty_1_66; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7639 = _GEN_774 ? _GEN_6741 : dirty_1_67; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7640 = _GEN_774 ? _GEN_6742 : dirty_1_68; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7641 = _GEN_774 ? _GEN_6743 : dirty_1_69; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7642 = _GEN_774 ? _GEN_6744 : dirty_1_70; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7643 = _GEN_774 ? _GEN_6745 : dirty_1_71; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7644 = _GEN_774 ? _GEN_6746 : dirty_1_72; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7645 = _GEN_774 ? _GEN_6747 : dirty_1_73; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7646 = _GEN_774 ? _GEN_6748 : dirty_1_74; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7647 = _GEN_774 ? _GEN_6749 : dirty_1_75; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7648 = _GEN_774 ? _GEN_6750 : dirty_1_76; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7649 = _GEN_774 ? _GEN_6751 : dirty_1_77; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7650 = _GEN_774 ? _GEN_6752 : dirty_1_78; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7651 = _GEN_774 ? _GEN_6753 : dirty_1_79; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7652 = _GEN_774 ? _GEN_6754 : dirty_1_80; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7653 = _GEN_774 ? _GEN_6755 : dirty_1_81; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7654 = _GEN_774 ? _GEN_6756 : dirty_1_82; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7655 = _GEN_774 ? _GEN_6757 : dirty_1_83; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7656 = _GEN_774 ? _GEN_6758 : dirty_1_84; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7657 = _GEN_774 ? _GEN_6759 : dirty_1_85; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7658 = _GEN_774 ? _GEN_6760 : dirty_1_86; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7659 = _GEN_774 ? _GEN_6761 : dirty_1_87; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7660 = _GEN_774 ? _GEN_6762 : dirty_1_88; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7661 = _GEN_774 ? _GEN_6763 : dirty_1_89; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7662 = _GEN_774 ? _GEN_6764 : dirty_1_90; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7663 = _GEN_774 ? _GEN_6765 : dirty_1_91; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7664 = _GEN_774 ? _GEN_6766 : dirty_1_92; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7665 = _GEN_774 ? _GEN_6767 : dirty_1_93; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7666 = _GEN_774 ? _GEN_6768 : dirty_1_94; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7667 = _GEN_774 ? _GEN_6769 : dirty_1_95; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7668 = _GEN_774 ? _GEN_6770 : dirty_1_96; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7669 = _GEN_774 ? _GEN_6771 : dirty_1_97; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7670 = _GEN_774 ? _GEN_6772 : dirty_1_98; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7671 = _GEN_774 ? _GEN_6773 : dirty_1_99; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7672 = _GEN_774 ? _GEN_6774 : dirty_1_100; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7673 = _GEN_774 ? _GEN_6775 : dirty_1_101; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7674 = _GEN_774 ? _GEN_6776 : dirty_1_102; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7675 = _GEN_774 ? _GEN_6777 : dirty_1_103; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7676 = _GEN_774 ? _GEN_6778 : dirty_1_104; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7677 = _GEN_774 ? _GEN_6779 : dirty_1_105; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7678 = _GEN_774 ? _GEN_6780 : dirty_1_106; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7679 = _GEN_774 ? _GEN_6781 : dirty_1_107; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7680 = _GEN_774 ? _GEN_6782 : dirty_1_108; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7681 = _GEN_774 ? _GEN_6783 : dirty_1_109; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7682 = _GEN_774 ? _GEN_6784 : dirty_1_110; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7683 = _GEN_774 ? _GEN_6785 : dirty_1_111; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7684 = _GEN_774 ? _GEN_6786 : dirty_1_112; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7685 = _GEN_774 ? _GEN_6787 : dirty_1_113; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7686 = _GEN_774 ? _GEN_6788 : dirty_1_114; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7687 = _GEN_774 ? _GEN_6789 : dirty_1_115; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7688 = _GEN_774 ? _GEN_6790 : dirty_1_116; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7689 = _GEN_774 ? _GEN_6791 : dirty_1_117; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7690 = _GEN_774 ? _GEN_6792 : dirty_1_118; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7691 = _GEN_774 ? _GEN_6793 : dirty_1_119; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7692 = _GEN_774 ? _GEN_6794 : dirty_1_120; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7693 = _GEN_774 ? _GEN_6795 : dirty_1_121; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7694 = _GEN_774 ? _GEN_6796 : dirty_1_122; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7695 = _GEN_774 ? _GEN_6797 : dirty_1_123; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7696 = _GEN_774 ? _GEN_6798 : dirty_1_124; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7697 = _GEN_774 ? _GEN_6799 : dirty_1_125; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7698 = _GEN_774 ? _GEN_6800 : dirty_1_126; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7699 = _GEN_774 ? _GEN_6801 : dirty_1_127; // @[d_cache.scala 182:47 33:26]
  wire  _GEN_7700 = _GEN_774 ? _GEN_4878 : _GEN_4878; // @[d_cache.scala 182:47]
  wire  _GEN_7701 = _GEN_774 ? _GEN_4879 : _GEN_4879; // @[d_cache.scala 182:47]
  wire  _GEN_7702 = _GEN_774 ? _GEN_4880 : _GEN_4880; // @[d_cache.scala 182:47]
  wire  _GEN_7703 = _GEN_774 ? _GEN_4881 : _GEN_4881; // @[d_cache.scala 182:47]
  wire  _GEN_7704 = _GEN_774 ? _GEN_4882 : _GEN_4882; // @[d_cache.scala 182:47]
  wire  _GEN_7705 = _GEN_774 ? _GEN_4883 : _GEN_4883; // @[d_cache.scala 182:47]
  wire  _GEN_7706 = _GEN_774 ? _GEN_4884 : _GEN_4884; // @[d_cache.scala 182:47]
  wire  _GEN_7707 = _GEN_774 ? _GEN_4885 : _GEN_4885; // @[d_cache.scala 182:47]
  wire  _GEN_7708 = _GEN_774 ? _GEN_4886 : _GEN_4886; // @[d_cache.scala 182:47]
  wire  _GEN_7709 = _GEN_774 ? _GEN_4887 : _GEN_4887; // @[d_cache.scala 182:47]
  wire  _GEN_7710 = _GEN_774 ? _GEN_4888 : _GEN_4888; // @[d_cache.scala 182:47]
  wire  _GEN_7711 = _GEN_774 ? _GEN_4889 : _GEN_4889; // @[d_cache.scala 182:47]
  wire  _GEN_7712 = _GEN_774 ? _GEN_4890 : _GEN_4890; // @[d_cache.scala 182:47]
  wire  _GEN_7713 = _GEN_774 ? _GEN_4891 : _GEN_4891; // @[d_cache.scala 182:47]
  wire  _GEN_7714 = _GEN_774 ? _GEN_4892 : _GEN_4892; // @[d_cache.scala 182:47]
  wire  _GEN_7715 = _GEN_774 ? _GEN_4893 : _GEN_4893; // @[d_cache.scala 182:47]
  wire  _GEN_7716 = _GEN_774 ? _GEN_4894 : _GEN_4894; // @[d_cache.scala 182:47]
  wire  _GEN_7717 = _GEN_774 ? _GEN_4895 : _GEN_4895; // @[d_cache.scala 182:47]
  wire  _GEN_7718 = _GEN_774 ? _GEN_4896 : _GEN_4896; // @[d_cache.scala 182:47]
  wire  _GEN_7719 = _GEN_774 ? _GEN_4897 : _GEN_4897; // @[d_cache.scala 182:47]
  wire  _GEN_7720 = _GEN_774 ? _GEN_4898 : _GEN_4898; // @[d_cache.scala 182:47]
  wire  _GEN_7721 = _GEN_774 ? _GEN_4899 : _GEN_4899; // @[d_cache.scala 182:47]
  wire  _GEN_7722 = _GEN_774 ? _GEN_4900 : _GEN_4900; // @[d_cache.scala 182:47]
  wire  _GEN_7723 = _GEN_774 ? _GEN_4901 : _GEN_4901; // @[d_cache.scala 182:47]
  wire  _GEN_7724 = _GEN_774 ? _GEN_4902 : _GEN_4902; // @[d_cache.scala 182:47]
  wire  _GEN_7725 = _GEN_774 ? _GEN_4903 : _GEN_4903; // @[d_cache.scala 182:47]
  wire  _GEN_7726 = _GEN_774 ? _GEN_4904 : _GEN_4904; // @[d_cache.scala 182:47]
  wire  _GEN_7727 = _GEN_774 ? _GEN_4905 : _GEN_4905; // @[d_cache.scala 182:47]
  wire  _GEN_7728 = _GEN_774 ? _GEN_4906 : _GEN_4906; // @[d_cache.scala 182:47]
  wire  _GEN_7729 = _GEN_774 ? _GEN_4907 : _GEN_4907; // @[d_cache.scala 182:47]
  wire  _GEN_7730 = _GEN_774 ? _GEN_4908 : _GEN_4908; // @[d_cache.scala 182:47]
  wire  _GEN_7731 = _GEN_774 ? _GEN_4909 : _GEN_4909; // @[d_cache.scala 182:47]
  wire  _GEN_7732 = _GEN_774 ? _GEN_4910 : _GEN_4910; // @[d_cache.scala 182:47]
  wire  _GEN_7733 = _GEN_774 ? _GEN_4911 : _GEN_4911; // @[d_cache.scala 182:47]
  wire  _GEN_7734 = _GEN_774 ? _GEN_4912 : _GEN_4912; // @[d_cache.scala 182:47]
  wire  _GEN_7735 = _GEN_774 ? _GEN_4913 : _GEN_4913; // @[d_cache.scala 182:47]
  wire  _GEN_7736 = _GEN_774 ? _GEN_4914 : _GEN_4914; // @[d_cache.scala 182:47]
  wire  _GEN_7737 = _GEN_774 ? _GEN_4915 : _GEN_4915; // @[d_cache.scala 182:47]
  wire  _GEN_7738 = _GEN_774 ? _GEN_4916 : _GEN_4916; // @[d_cache.scala 182:47]
  wire  _GEN_7739 = _GEN_774 ? _GEN_4917 : _GEN_4917; // @[d_cache.scala 182:47]
  wire  _GEN_7740 = _GEN_774 ? _GEN_4918 : _GEN_4918; // @[d_cache.scala 182:47]
  wire  _GEN_7741 = _GEN_774 ? _GEN_4919 : _GEN_4919; // @[d_cache.scala 182:47]
  wire  _GEN_7742 = _GEN_774 ? _GEN_4920 : _GEN_4920; // @[d_cache.scala 182:47]
  wire  _GEN_7743 = _GEN_774 ? _GEN_4921 : _GEN_4921; // @[d_cache.scala 182:47]
  wire  _GEN_7744 = _GEN_774 ? _GEN_4922 : _GEN_4922; // @[d_cache.scala 182:47]
  wire  _GEN_7745 = _GEN_774 ? _GEN_4923 : _GEN_4923; // @[d_cache.scala 182:47]
  wire  _GEN_7746 = _GEN_774 ? _GEN_4924 : _GEN_4924; // @[d_cache.scala 182:47]
  wire  _GEN_7747 = _GEN_774 ? _GEN_4925 : _GEN_4925; // @[d_cache.scala 182:47]
  wire  _GEN_7748 = _GEN_774 ? _GEN_4926 : _GEN_4926; // @[d_cache.scala 182:47]
  wire  _GEN_7749 = _GEN_774 ? _GEN_4927 : _GEN_4927; // @[d_cache.scala 182:47]
  wire  _GEN_7750 = _GEN_774 ? _GEN_4928 : _GEN_4928; // @[d_cache.scala 182:47]
  wire  _GEN_7751 = _GEN_774 ? _GEN_4929 : _GEN_4929; // @[d_cache.scala 182:47]
  wire  _GEN_7752 = _GEN_774 ? _GEN_4930 : _GEN_4930; // @[d_cache.scala 182:47]
  wire  _GEN_7753 = _GEN_774 ? _GEN_4931 : _GEN_4931; // @[d_cache.scala 182:47]
  wire  _GEN_7754 = _GEN_774 ? _GEN_4932 : _GEN_4932; // @[d_cache.scala 182:47]
  wire  _GEN_7755 = _GEN_774 ? _GEN_4933 : _GEN_4933; // @[d_cache.scala 182:47]
  wire  _GEN_7756 = _GEN_774 ? _GEN_4934 : _GEN_4934; // @[d_cache.scala 182:47]
  wire  _GEN_7757 = _GEN_774 ? _GEN_4935 : _GEN_4935; // @[d_cache.scala 182:47]
  wire  _GEN_7758 = _GEN_774 ? _GEN_4936 : _GEN_4936; // @[d_cache.scala 182:47]
  wire  _GEN_7759 = _GEN_774 ? _GEN_4937 : _GEN_4937; // @[d_cache.scala 182:47]
  wire  _GEN_7760 = _GEN_774 ? _GEN_4938 : _GEN_4938; // @[d_cache.scala 182:47]
  wire  _GEN_7761 = _GEN_774 ? _GEN_4939 : _GEN_4939; // @[d_cache.scala 182:47]
  wire  _GEN_7762 = _GEN_774 ? _GEN_4940 : _GEN_4940; // @[d_cache.scala 182:47]
  wire  _GEN_7763 = _GEN_774 ? _GEN_4941 : _GEN_4941; // @[d_cache.scala 182:47]
  wire  _GEN_7764 = _GEN_774 ? _GEN_4942 : _GEN_4942; // @[d_cache.scala 182:47]
  wire  _GEN_7765 = _GEN_774 ? _GEN_4943 : _GEN_4943; // @[d_cache.scala 182:47]
  wire  _GEN_7766 = _GEN_774 ? _GEN_4944 : _GEN_4944; // @[d_cache.scala 182:47]
  wire  _GEN_7767 = _GEN_774 ? _GEN_4945 : _GEN_4945; // @[d_cache.scala 182:47]
  wire  _GEN_7768 = _GEN_774 ? _GEN_4946 : _GEN_4946; // @[d_cache.scala 182:47]
  wire  _GEN_7769 = _GEN_774 ? _GEN_4947 : _GEN_4947; // @[d_cache.scala 182:47]
  wire  _GEN_7770 = _GEN_774 ? _GEN_4948 : _GEN_4948; // @[d_cache.scala 182:47]
  wire  _GEN_7771 = _GEN_774 ? _GEN_4949 : _GEN_4949; // @[d_cache.scala 182:47]
  wire  _GEN_7772 = _GEN_774 ? _GEN_4950 : _GEN_4950; // @[d_cache.scala 182:47]
  wire  _GEN_7773 = _GEN_774 ? _GEN_4951 : _GEN_4951; // @[d_cache.scala 182:47]
  wire  _GEN_7774 = _GEN_774 ? _GEN_4952 : _GEN_4952; // @[d_cache.scala 182:47]
  wire  _GEN_7775 = _GEN_774 ? _GEN_4953 : _GEN_4953; // @[d_cache.scala 182:47]
  wire  _GEN_7776 = _GEN_774 ? _GEN_4954 : _GEN_4954; // @[d_cache.scala 182:47]
  wire  _GEN_7777 = _GEN_774 ? _GEN_4955 : _GEN_4955; // @[d_cache.scala 182:47]
  wire  _GEN_7778 = _GEN_774 ? _GEN_4956 : _GEN_4956; // @[d_cache.scala 182:47]
  wire  _GEN_7779 = _GEN_774 ? _GEN_4957 : _GEN_4957; // @[d_cache.scala 182:47]
  wire  _GEN_7780 = _GEN_774 ? _GEN_4958 : _GEN_4958; // @[d_cache.scala 182:47]
  wire  _GEN_7781 = _GEN_774 ? _GEN_4959 : _GEN_4959; // @[d_cache.scala 182:47]
  wire  _GEN_7782 = _GEN_774 ? _GEN_4960 : _GEN_4960; // @[d_cache.scala 182:47]
  wire  _GEN_7783 = _GEN_774 ? _GEN_4961 : _GEN_4961; // @[d_cache.scala 182:47]
  wire  _GEN_7784 = _GEN_774 ? _GEN_4962 : _GEN_4962; // @[d_cache.scala 182:47]
  wire  _GEN_7785 = _GEN_774 ? _GEN_4963 : _GEN_4963; // @[d_cache.scala 182:47]
  wire  _GEN_7786 = _GEN_774 ? _GEN_4964 : _GEN_4964; // @[d_cache.scala 182:47]
  wire  _GEN_7787 = _GEN_774 ? _GEN_4965 : _GEN_4965; // @[d_cache.scala 182:47]
  wire  _GEN_7788 = _GEN_774 ? _GEN_4966 : _GEN_4966; // @[d_cache.scala 182:47]
  wire  _GEN_7789 = _GEN_774 ? _GEN_4967 : _GEN_4967; // @[d_cache.scala 182:47]
  wire  _GEN_7790 = _GEN_774 ? _GEN_4968 : _GEN_4968; // @[d_cache.scala 182:47]
  wire  _GEN_7791 = _GEN_774 ? _GEN_4969 : _GEN_4969; // @[d_cache.scala 182:47]
  wire  _GEN_7792 = _GEN_774 ? _GEN_4970 : _GEN_4970; // @[d_cache.scala 182:47]
  wire  _GEN_7793 = _GEN_774 ? _GEN_4971 : _GEN_4971; // @[d_cache.scala 182:47]
  wire  _GEN_7794 = _GEN_774 ? _GEN_4972 : _GEN_4972; // @[d_cache.scala 182:47]
  wire  _GEN_7795 = _GEN_774 ? _GEN_4973 : _GEN_4973; // @[d_cache.scala 182:47]
  wire  _GEN_7796 = _GEN_774 ? _GEN_4974 : _GEN_4974; // @[d_cache.scala 182:47]
  wire  _GEN_7797 = _GEN_774 ? _GEN_4975 : _GEN_4975; // @[d_cache.scala 182:47]
  wire  _GEN_7798 = _GEN_774 ? _GEN_4976 : _GEN_4976; // @[d_cache.scala 182:47]
  wire  _GEN_7799 = _GEN_774 ? _GEN_4977 : _GEN_4977; // @[d_cache.scala 182:47]
  wire  _GEN_7800 = _GEN_774 ? _GEN_4978 : _GEN_4978; // @[d_cache.scala 182:47]
  wire  _GEN_7801 = _GEN_774 ? _GEN_4979 : _GEN_4979; // @[d_cache.scala 182:47]
  wire  _GEN_7802 = _GEN_774 ? _GEN_4980 : _GEN_4980; // @[d_cache.scala 182:47]
  wire  _GEN_7803 = _GEN_774 ? _GEN_4981 : _GEN_4981; // @[d_cache.scala 182:47]
  wire  _GEN_7804 = _GEN_774 ? _GEN_4982 : _GEN_4982; // @[d_cache.scala 182:47]
  wire  _GEN_7805 = _GEN_774 ? _GEN_4983 : _GEN_4983; // @[d_cache.scala 182:47]
  wire  _GEN_7806 = _GEN_774 ? _GEN_4984 : _GEN_4984; // @[d_cache.scala 182:47]
  wire  _GEN_7807 = _GEN_774 ? _GEN_4985 : _GEN_4985; // @[d_cache.scala 182:47]
  wire  _GEN_7808 = _GEN_774 ? _GEN_4986 : _GEN_4986; // @[d_cache.scala 182:47]
  wire  _GEN_7809 = _GEN_774 ? _GEN_4987 : _GEN_4987; // @[d_cache.scala 182:47]
  wire  _GEN_7810 = _GEN_774 ? _GEN_4988 : _GEN_4988; // @[d_cache.scala 182:47]
  wire  _GEN_7811 = _GEN_774 ? _GEN_4989 : _GEN_4989; // @[d_cache.scala 182:47]
  wire  _GEN_7812 = _GEN_774 ? _GEN_4990 : _GEN_4990; // @[d_cache.scala 182:47]
  wire  _GEN_7813 = _GEN_774 ? _GEN_4991 : _GEN_4991; // @[d_cache.scala 182:47]
  wire  _GEN_7814 = _GEN_774 ? _GEN_4992 : _GEN_4992; // @[d_cache.scala 182:47]
  wire  _GEN_7815 = _GEN_774 ? _GEN_4993 : _GEN_4993; // @[d_cache.scala 182:47]
  wire  _GEN_7816 = _GEN_774 ? _GEN_4994 : _GEN_4994; // @[d_cache.scala 182:47]
  wire  _GEN_7817 = _GEN_774 ? _GEN_4995 : _GEN_4995; // @[d_cache.scala 182:47]
  wire  _GEN_7818 = _GEN_774 ? _GEN_4996 : _GEN_4996; // @[d_cache.scala 182:47]
  wire  _GEN_7819 = _GEN_774 ? _GEN_4997 : _GEN_4997; // @[d_cache.scala 182:47]
  wire  _GEN_7820 = _GEN_774 ? _GEN_4998 : _GEN_4998; // @[d_cache.scala 182:47]
  wire  _GEN_7821 = _GEN_774 ? _GEN_4999 : _GEN_4999; // @[d_cache.scala 182:47]
  wire  _GEN_7822 = _GEN_774 ? _GEN_5000 : _GEN_5000; // @[d_cache.scala 182:47]
  wire  _GEN_7823 = _GEN_774 ? _GEN_5001 : _GEN_5001; // @[d_cache.scala 182:47]
  wire  _GEN_7824 = _GEN_774 ? _GEN_5002 : _GEN_5002; // @[d_cache.scala 182:47]
  wire  _GEN_7825 = _GEN_774 ? _GEN_5003 : _GEN_5003; // @[d_cache.scala 182:47]
  wire  _GEN_7826 = _GEN_774 ? _GEN_5004 : _GEN_5004; // @[d_cache.scala 182:47]
  wire  _GEN_7827 = _GEN_774 ? _GEN_5005 : _GEN_5005; // @[d_cache.scala 182:47]
  wire [2:0] _GEN_7828 = _GEN_774 ? 3'h6 : 3'h7; // @[d_cache.scala 182:47 189:31 192:31]
  wire [63:0] _GEN_7830 = ~quene ? _GEN_5902 : _GEN_7314; // @[d_cache.scala 163:34]
  wire [41:0] _GEN_7831 = ~quene ? _GEN_5903 : _GEN_7315; // @[d_cache.scala 163:34]
  wire [63:0] _GEN_7832 = ~quene ? _GEN_5904 : ram_0_0; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7833 = ~quene ? _GEN_5905 : ram_0_1; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7834 = ~quene ? _GEN_5906 : ram_0_2; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7835 = ~quene ? _GEN_5907 : ram_0_3; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7836 = ~quene ? _GEN_5908 : ram_0_4; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7837 = ~quene ? _GEN_5909 : ram_0_5; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7838 = ~quene ? _GEN_5910 : ram_0_6; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7839 = ~quene ? _GEN_5911 : ram_0_7; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7840 = ~quene ? _GEN_5912 : ram_0_8; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7841 = ~quene ? _GEN_5913 : ram_0_9; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7842 = ~quene ? _GEN_5914 : ram_0_10; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7843 = ~quene ? _GEN_5915 : ram_0_11; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7844 = ~quene ? _GEN_5916 : ram_0_12; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7845 = ~quene ? _GEN_5917 : ram_0_13; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7846 = ~quene ? _GEN_5918 : ram_0_14; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7847 = ~quene ? _GEN_5919 : ram_0_15; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7848 = ~quene ? _GEN_5920 : ram_0_16; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7849 = ~quene ? _GEN_5921 : ram_0_17; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7850 = ~quene ? _GEN_5922 : ram_0_18; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7851 = ~quene ? _GEN_5923 : ram_0_19; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7852 = ~quene ? _GEN_5924 : ram_0_20; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7853 = ~quene ? _GEN_5925 : ram_0_21; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7854 = ~quene ? _GEN_5926 : ram_0_22; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7855 = ~quene ? _GEN_5927 : ram_0_23; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7856 = ~quene ? _GEN_5928 : ram_0_24; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7857 = ~quene ? _GEN_5929 : ram_0_25; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7858 = ~quene ? _GEN_5930 : ram_0_26; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7859 = ~quene ? _GEN_5931 : ram_0_27; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7860 = ~quene ? _GEN_5932 : ram_0_28; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7861 = ~quene ? _GEN_5933 : ram_0_29; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7862 = ~quene ? _GEN_5934 : ram_0_30; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7863 = ~quene ? _GEN_5935 : ram_0_31; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7864 = ~quene ? _GEN_5936 : ram_0_32; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7865 = ~quene ? _GEN_5937 : ram_0_33; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7866 = ~quene ? _GEN_5938 : ram_0_34; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7867 = ~quene ? _GEN_5939 : ram_0_35; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7868 = ~quene ? _GEN_5940 : ram_0_36; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7869 = ~quene ? _GEN_5941 : ram_0_37; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7870 = ~quene ? _GEN_5942 : ram_0_38; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7871 = ~quene ? _GEN_5943 : ram_0_39; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7872 = ~quene ? _GEN_5944 : ram_0_40; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7873 = ~quene ? _GEN_5945 : ram_0_41; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7874 = ~quene ? _GEN_5946 : ram_0_42; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7875 = ~quene ? _GEN_5947 : ram_0_43; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7876 = ~quene ? _GEN_5948 : ram_0_44; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7877 = ~quene ? _GEN_5949 : ram_0_45; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7878 = ~quene ? _GEN_5950 : ram_0_46; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7879 = ~quene ? _GEN_5951 : ram_0_47; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7880 = ~quene ? _GEN_5952 : ram_0_48; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7881 = ~quene ? _GEN_5953 : ram_0_49; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7882 = ~quene ? _GEN_5954 : ram_0_50; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7883 = ~quene ? _GEN_5955 : ram_0_51; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7884 = ~quene ? _GEN_5956 : ram_0_52; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7885 = ~quene ? _GEN_5957 : ram_0_53; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7886 = ~quene ? _GEN_5958 : ram_0_54; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7887 = ~quene ? _GEN_5959 : ram_0_55; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7888 = ~quene ? _GEN_5960 : ram_0_56; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7889 = ~quene ? _GEN_5961 : ram_0_57; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7890 = ~quene ? _GEN_5962 : ram_0_58; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7891 = ~quene ? _GEN_5963 : ram_0_59; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7892 = ~quene ? _GEN_5964 : ram_0_60; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7893 = ~quene ? _GEN_5965 : ram_0_61; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7894 = ~quene ? _GEN_5966 : ram_0_62; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7895 = ~quene ? _GEN_5967 : ram_0_63; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7896 = ~quene ? _GEN_5968 : ram_0_64; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7897 = ~quene ? _GEN_5969 : ram_0_65; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7898 = ~quene ? _GEN_5970 : ram_0_66; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7899 = ~quene ? _GEN_5971 : ram_0_67; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7900 = ~quene ? _GEN_5972 : ram_0_68; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7901 = ~quene ? _GEN_5973 : ram_0_69; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7902 = ~quene ? _GEN_5974 : ram_0_70; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7903 = ~quene ? _GEN_5975 : ram_0_71; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7904 = ~quene ? _GEN_5976 : ram_0_72; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7905 = ~quene ? _GEN_5977 : ram_0_73; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7906 = ~quene ? _GEN_5978 : ram_0_74; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7907 = ~quene ? _GEN_5979 : ram_0_75; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7908 = ~quene ? _GEN_5980 : ram_0_76; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7909 = ~quene ? _GEN_5981 : ram_0_77; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7910 = ~quene ? _GEN_5982 : ram_0_78; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7911 = ~quene ? _GEN_5983 : ram_0_79; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7912 = ~quene ? _GEN_5984 : ram_0_80; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7913 = ~quene ? _GEN_5985 : ram_0_81; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7914 = ~quene ? _GEN_5986 : ram_0_82; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7915 = ~quene ? _GEN_5987 : ram_0_83; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7916 = ~quene ? _GEN_5988 : ram_0_84; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7917 = ~quene ? _GEN_5989 : ram_0_85; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7918 = ~quene ? _GEN_5990 : ram_0_86; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7919 = ~quene ? _GEN_5991 : ram_0_87; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7920 = ~quene ? _GEN_5992 : ram_0_88; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7921 = ~quene ? _GEN_5993 : ram_0_89; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7922 = ~quene ? _GEN_5994 : ram_0_90; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7923 = ~quene ? _GEN_5995 : ram_0_91; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7924 = ~quene ? _GEN_5996 : ram_0_92; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7925 = ~quene ? _GEN_5997 : ram_0_93; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7926 = ~quene ? _GEN_5998 : ram_0_94; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7927 = ~quene ? _GEN_5999 : ram_0_95; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7928 = ~quene ? _GEN_6000 : ram_0_96; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7929 = ~quene ? _GEN_6001 : ram_0_97; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7930 = ~quene ? _GEN_6002 : ram_0_98; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7931 = ~quene ? _GEN_6003 : ram_0_99; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7932 = ~quene ? _GEN_6004 : ram_0_100; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7933 = ~quene ? _GEN_6005 : ram_0_101; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7934 = ~quene ? _GEN_6006 : ram_0_102; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7935 = ~quene ? _GEN_6007 : ram_0_103; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7936 = ~quene ? _GEN_6008 : ram_0_104; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7937 = ~quene ? _GEN_6009 : ram_0_105; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7938 = ~quene ? _GEN_6010 : ram_0_106; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7939 = ~quene ? _GEN_6011 : ram_0_107; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7940 = ~quene ? _GEN_6012 : ram_0_108; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7941 = ~quene ? _GEN_6013 : ram_0_109; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7942 = ~quene ? _GEN_6014 : ram_0_110; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7943 = ~quene ? _GEN_6015 : ram_0_111; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7944 = ~quene ? _GEN_6016 : ram_0_112; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7945 = ~quene ? _GEN_6017 : ram_0_113; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7946 = ~quene ? _GEN_6018 : ram_0_114; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7947 = ~quene ? _GEN_6019 : ram_0_115; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7948 = ~quene ? _GEN_6020 : ram_0_116; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7949 = ~quene ? _GEN_6021 : ram_0_117; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7950 = ~quene ? _GEN_6022 : ram_0_118; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7951 = ~quene ? _GEN_6023 : ram_0_119; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7952 = ~quene ? _GEN_6024 : ram_0_120; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7953 = ~quene ? _GEN_6025 : ram_0_121; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7954 = ~quene ? _GEN_6026 : ram_0_122; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7955 = ~quene ? _GEN_6027 : ram_0_123; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7956 = ~quene ? _GEN_6028 : ram_0_124; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7957 = ~quene ? _GEN_6029 : ram_0_125; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7958 = ~quene ? _GEN_6030 : ram_0_126; // @[d_cache.scala 163:34 19:24]
  wire [63:0] _GEN_7959 = ~quene ? _GEN_6031 : ram_0_127; // @[d_cache.scala 163:34 19:24]
  wire [31:0] _GEN_7960 = ~quene ? _GEN_6032 : tag_0_0; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7961 = ~quene ? _GEN_6033 : tag_0_1; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7962 = ~quene ? _GEN_6034 : tag_0_2; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7963 = ~quene ? _GEN_6035 : tag_0_3; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7964 = ~quene ? _GEN_6036 : tag_0_4; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7965 = ~quene ? _GEN_6037 : tag_0_5; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7966 = ~quene ? _GEN_6038 : tag_0_6; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7967 = ~quene ? _GEN_6039 : tag_0_7; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7968 = ~quene ? _GEN_6040 : tag_0_8; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7969 = ~quene ? _GEN_6041 : tag_0_9; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7970 = ~quene ? _GEN_6042 : tag_0_10; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7971 = ~quene ? _GEN_6043 : tag_0_11; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7972 = ~quene ? _GEN_6044 : tag_0_12; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7973 = ~quene ? _GEN_6045 : tag_0_13; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7974 = ~quene ? _GEN_6046 : tag_0_14; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7975 = ~quene ? _GEN_6047 : tag_0_15; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7976 = ~quene ? _GEN_6048 : tag_0_16; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7977 = ~quene ? _GEN_6049 : tag_0_17; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7978 = ~quene ? _GEN_6050 : tag_0_18; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7979 = ~quene ? _GEN_6051 : tag_0_19; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7980 = ~quene ? _GEN_6052 : tag_0_20; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7981 = ~quene ? _GEN_6053 : tag_0_21; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7982 = ~quene ? _GEN_6054 : tag_0_22; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7983 = ~quene ? _GEN_6055 : tag_0_23; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7984 = ~quene ? _GEN_6056 : tag_0_24; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7985 = ~quene ? _GEN_6057 : tag_0_25; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7986 = ~quene ? _GEN_6058 : tag_0_26; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7987 = ~quene ? _GEN_6059 : tag_0_27; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7988 = ~quene ? _GEN_6060 : tag_0_28; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7989 = ~quene ? _GEN_6061 : tag_0_29; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7990 = ~quene ? _GEN_6062 : tag_0_30; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7991 = ~quene ? _GEN_6063 : tag_0_31; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7992 = ~quene ? _GEN_6064 : tag_0_32; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7993 = ~quene ? _GEN_6065 : tag_0_33; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7994 = ~quene ? _GEN_6066 : tag_0_34; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7995 = ~quene ? _GEN_6067 : tag_0_35; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7996 = ~quene ? _GEN_6068 : tag_0_36; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7997 = ~quene ? _GEN_6069 : tag_0_37; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7998 = ~quene ? _GEN_6070 : tag_0_38; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_7999 = ~quene ? _GEN_6071 : tag_0_39; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8000 = ~quene ? _GEN_6072 : tag_0_40; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8001 = ~quene ? _GEN_6073 : tag_0_41; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8002 = ~quene ? _GEN_6074 : tag_0_42; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8003 = ~quene ? _GEN_6075 : tag_0_43; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8004 = ~quene ? _GEN_6076 : tag_0_44; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8005 = ~quene ? _GEN_6077 : tag_0_45; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8006 = ~quene ? _GEN_6078 : tag_0_46; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8007 = ~quene ? _GEN_6079 : tag_0_47; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8008 = ~quene ? _GEN_6080 : tag_0_48; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8009 = ~quene ? _GEN_6081 : tag_0_49; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8010 = ~quene ? _GEN_6082 : tag_0_50; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8011 = ~quene ? _GEN_6083 : tag_0_51; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8012 = ~quene ? _GEN_6084 : tag_0_52; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8013 = ~quene ? _GEN_6085 : tag_0_53; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8014 = ~quene ? _GEN_6086 : tag_0_54; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8015 = ~quene ? _GEN_6087 : tag_0_55; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8016 = ~quene ? _GEN_6088 : tag_0_56; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8017 = ~quene ? _GEN_6089 : tag_0_57; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8018 = ~quene ? _GEN_6090 : tag_0_58; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8019 = ~quene ? _GEN_6091 : tag_0_59; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8020 = ~quene ? _GEN_6092 : tag_0_60; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8021 = ~quene ? _GEN_6093 : tag_0_61; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8022 = ~quene ? _GEN_6094 : tag_0_62; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8023 = ~quene ? _GEN_6095 : tag_0_63; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8024 = ~quene ? _GEN_6096 : tag_0_64; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8025 = ~quene ? _GEN_6097 : tag_0_65; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8026 = ~quene ? _GEN_6098 : tag_0_66; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8027 = ~quene ? _GEN_6099 : tag_0_67; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8028 = ~quene ? _GEN_6100 : tag_0_68; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8029 = ~quene ? _GEN_6101 : tag_0_69; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8030 = ~quene ? _GEN_6102 : tag_0_70; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8031 = ~quene ? _GEN_6103 : tag_0_71; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8032 = ~quene ? _GEN_6104 : tag_0_72; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8033 = ~quene ? _GEN_6105 : tag_0_73; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8034 = ~quene ? _GEN_6106 : tag_0_74; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8035 = ~quene ? _GEN_6107 : tag_0_75; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8036 = ~quene ? _GEN_6108 : tag_0_76; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8037 = ~quene ? _GEN_6109 : tag_0_77; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8038 = ~quene ? _GEN_6110 : tag_0_78; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8039 = ~quene ? _GEN_6111 : tag_0_79; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8040 = ~quene ? _GEN_6112 : tag_0_80; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8041 = ~quene ? _GEN_6113 : tag_0_81; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8042 = ~quene ? _GEN_6114 : tag_0_82; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8043 = ~quene ? _GEN_6115 : tag_0_83; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8044 = ~quene ? _GEN_6116 : tag_0_84; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8045 = ~quene ? _GEN_6117 : tag_0_85; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8046 = ~quene ? _GEN_6118 : tag_0_86; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8047 = ~quene ? _GEN_6119 : tag_0_87; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8048 = ~quene ? _GEN_6120 : tag_0_88; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8049 = ~quene ? _GEN_6121 : tag_0_89; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8050 = ~quene ? _GEN_6122 : tag_0_90; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8051 = ~quene ? _GEN_6123 : tag_0_91; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8052 = ~quene ? _GEN_6124 : tag_0_92; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8053 = ~quene ? _GEN_6125 : tag_0_93; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8054 = ~quene ? _GEN_6126 : tag_0_94; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8055 = ~quene ? _GEN_6127 : tag_0_95; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8056 = ~quene ? _GEN_6128 : tag_0_96; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8057 = ~quene ? _GEN_6129 : tag_0_97; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8058 = ~quene ? _GEN_6130 : tag_0_98; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8059 = ~quene ? _GEN_6131 : tag_0_99; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8060 = ~quene ? _GEN_6132 : tag_0_100; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8061 = ~quene ? _GEN_6133 : tag_0_101; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8062 = ~quene ? _GEN_6134 : tag_0_102; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8063 = ~quene ? _GEN_6135 : tag_0_103; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8064 = ~quene ? _GEN_6136 : tag_0_104; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8065 = ~quene ? _GEN_6137 : tag_0_105; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8066 = ~quene ? _GEN_6138 : tag_0_106; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8067 = ~quene ? _GEN_6139 : tag_0_107; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8068 = ~quene ? _GEN_6140 : tag_0_108; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8069 = ~quene ? _GEN_6141 : tag_0_109; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8070 = ~quene ? _GEN_6142 : tag_0_110; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8071 = ~quene ? _GEN_6143 : tag_0_111; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8072 = ~quene ? _GEN_6144 : tag_0_112; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8073 = ~quene ? _GEN_6145 : tag_0_113; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8074 = ~quene ? _GEN_6146 : tag_0_114; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8075 = ~quene ? _GEN_6147 : tag_0_115; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8076 = ~quene ? _GEN_6148 : tag_0_116; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8077 = ~quene ? _GEN_6149 : tag_0_117; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8078 = ~quene ? _GEN_6150 : tag_0_118; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8079 = ~quene ? _GEN_6151 : tag_0_119; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8080 = ~quene ? _GEN_6152 : tag_0_120; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8081 = ~quene ? _GEN_6153 : tag_0_121; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8082 = ~quene ? _GEN_6154 : tag_0_122; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8083 = ~quene ? _GEN_6155 : tag_0_123; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8084 = ~quene ? _GEN_6156 : tag_0_124; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8085 = ~quene ? _GEN_6157 : tag_0_125; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8086 = ~quene ? _GEN_6158 : tag_0_126; // @[d_cache.scala 163:34 28:24]
  wire [31:0] _GEN_8087 = ~quene ? _GEN_6159 : tag_0_127; // @[d_cache.scala 163:34 28:24]
  wire  _GEN_8088 = ~quene ? _GEN_6160 : dirty_0_0; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8089 = ~quene ? _GEN_6161 : dirty_0_1; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8090 = ~quene ? _GEN_6162 : dirty_0_2; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8091 = ~quene ? _GEN_6163 : dirty_0_3; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8092 = ~quene ? _GEN_6164 : dirty_0_4; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8093 = ~quene ? _GEN_6165 : dirty_0_5; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8094 = ~quene ? _GEN_6166 : dirty_0_6; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8095 = ~quene ? _GEN_6167 : dirty_0_7; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8096 = ~quene ? _GEN_6168 : dirty_0_8; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8097 = ~quene ? _GEN_6169 : dirty_0_9; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8098 = ~quene ? _GEN_6170 : dirty_0_10; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8099 = ~quene ? _GEN_6171 : dirty_0_11; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8100 = ~quene ? _GEN_6172 : dirty_0_12; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8101 = ~quene ? _GEN_6173 : dirty_0_13; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8102 = ~quene ? _GEN_6174 : dirty_0_14; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8103 = ~quene ? _GEN_6175 : dirty_0_15; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8104 = ~quene ? _GEN_6176 : dirty_0_16; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8105 = ~quene ? _GEN_6177 : dirty_0_17; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8106 = ~quene ? _GEN_6178 : dirty_0_18; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8107 = ~quene ? _GEN_6179 : dirty_0_19; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8108 = ~quene ? _GEN_6180 : dirty_0_20; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8109 = ~quene ? _GEN_6181 : dirty_0_21; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8110 = ~quene ? _GEN_6182 : dirty_0_22; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8111 = ~quene ? _GEN_6183 : dirty_0_23; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8112 = ~quene ? _GEN_6184 : dirty_0_24; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8113 = ~quene ? _GEN_6185 : dirty_0_25; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8114 = ~quene ? _GEN_6186 : dirty_0_26; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8115 = ~quene ? _GEN_6187 : dirty_0_27; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8116 = ~quene ? _GEN_6188 : dirty_0_28; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8117 = ~quene ? _GEN_6189 : dirty_0_29; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8118 = ~quene ? _GEN_6190 : dirty_0_30; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8119 = ~quene ? _GEN_6191 : dirty_0_31; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8120 = ~quene ? _GEN_6192 : dirty_0_32; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8121 = ~quene ? _GEN_6193 : dirty_0_33; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8122 = ~quene ? _GEN_6194 : dirty_0_34; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8123 = ~quene ? _GEN_6195 : dirty_0_35; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8124 = ~quene ? _GEN_6196 : dirty_0_36; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8125 = ~quene ? _GEN_6197 : dirty_0_37; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8126 = ~quene ? _GEN_6198 : dirty_0_38; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8127 = ~quene ? _GEN_6199 : dirty_0_39; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8128 = ~quene ? _GEN_6200 : dirty_0_40; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8129 = ~quene ? _GEN_6201 : dirty_0_41; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8130 = ~quene ? _GEN_6202 : dirty_0_42; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8131 = ~quene ? _GEN_6203 : dirty_0_43; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8132 = ~quene ? _GEN_6204 : dirty_0_44; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8133 = ~quene ? _GEN_6205 : dirty_0_45; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8134 = ~quene ? _GEN_6206 : dirty_0_46; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8135 = ~quene ? _GEN_6207 : dirty_0_47; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8136 = ~quene ? _GEN_6208 : dirty_0_48; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8137 = ~quene ? _GEN_6209 : dirty_0_49; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8138 = ~quene ? _GEN_6210 : dirty_0_50; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8139 = ~quene ? _GEN_6211 : dirty_0_51; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8140 = ~quene ? _GEN_6212 : dirty_0_52; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8141 = ~quene ? _GEN_6213 : dirty_0_53; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8142 = ~quene ? _GEN_6214 : dirty_0_54; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8143 = ~quene ? _GEN_6215 : dirty_0_55; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8144 = ~quene ? _GEN_6216 : dirty_0_56; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8145 = ~quene ? _GEN_6217 : dirty_0_57; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8146 = ~quene ? _GEN_6218 : dirty_0_58; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8147 = ~quene ? _GEN_6219 : dirty_0_59; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8148 = ~quene ? _GEN_6220 : dirty_0_60; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8149 = ~quene ? _GEN_6221 : dirty_0_61; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8150 = ~quene ? _GEN_6222 : dirty_0_62; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8151 = ~quene ? _GEN_6223 : dirty_0_63; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8152 = ~quene ? _GEN_6224 : dirty_0_64; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8153 = ~quene ? _GEN_6225 : dirty_0_65; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8154 = ~quene ? _GEN_6226 : dirty_0_66; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8155 = ~quene ? _GEN_6227 : dirty_0_67; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8156 = ~quene ? _GEN_6228 : dirty_0_68; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8157 = ~quene ? _GEN_6229 : dirty_0_69; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8158 = ~quene ? _GEN_6230 : dirty_0_70; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8159 = ~quene ? _GEN_6231 : dirty_0_71; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8160 = ~quene ? _GEN_6232 : dirty_0_72; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8161 = ~quene ? _GEN_6233 : dirty_0_73; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8162 = ~quene ? _GEN_6234 : dirty_0_74; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8163 = ~quene ? _GEN_6235 : dirty_0_75; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8164 = ~quene ? _GEN_6236 : dirty_0_76; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8165 = ~quene ? _GEN_6237 : dirty_0_77; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8166 = ~quene ? _GEN_6238 : dirty_0_78; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8167 = ~quene ? _GEN_6239 : dirty_0_79; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8168 = ~quene ? _GEN_6240 : dirty_0_80; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8169 = ~quene ? _GEN_6241 : dirty_0_81; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8170 = ~quene ? _GEN_6242 : dirty_0_82; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8171 = ~quene ? _GEN_6243 : dirty_0_83; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8172 = ~quene ? _GEN_6244 : dirty_0_84; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8173 = ~quene ? _GEN_6245 : dirty_0_85; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8174 = ~quene ? _GEN_6246 : dirty_0_86; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8175 = ~quene ? _GEN_6247 : dirty_0_87; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8176 = ~quene ? _GEN_6248 : dirty_0_88; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8177 = ~quene ? _GEN_6249 : dirty_0_89; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8178 = ~quene ? _GEN_6250 : dirty_0_90; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8179 = ~quene ? _GEN_6251 : dirty_0_91; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8180 = ~quene ? _GEN_6252 : dirty_0_92; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8181 = ~quene ? _GEN_6253 : dirty_0_93; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8182 = ~quene ? _GEN_6254 : dirty_0_94; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8183 = ~quene ? _GEN_6255 : dirty_0_95; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8184 = ~quene ? _GEN_6256 : dirty_0_96; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8185 = ~quene ? _GEN_6257 : dirty_0_97; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8186 = ~quene ? _GEN_6258 : dirty_0_98; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8187 = ~quene ? _GEN_6259 : dirty_0_99; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8188 = ~quene ? _GEN_6260 : dirty_0_100; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8189 = ~quene ? _GEN_6261 : dirty_0_101; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8190 = ~quene ? _GEN_6262 : dirty_0_102; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8191 = ~quene ? _GEN_6263 : dirty_0_103; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8192 = ~quene ? _GEN_6264 : dirty_0_104; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8193 = ~quene ? _GEN_6265 : dirty_0_105; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8194 = ~quene ? _GEN_6266 : dirty_0_106; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8195 = ~quene ? _GEN_6267 : dirty_0_107; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8196 = ~quene ? _GEN_6268 : dirty_0_108; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8197 = ~quene ? _GEN_6269 : dirty_0_109; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8198 = ~quene ? _GEN_6270 : dirty_0_110; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8199 = ~quene ? _GEN_6271 : dirty_0_111; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8200 = ~quene ? _GEN_6272 : dirty_0_112; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8201 = ~quene ? _GEN_6273 : dirty_0_113; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8202 = ~quene ? _GEN_6274 : dirty_0_114; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8203 = ~quene ? _GEN_6275 : dirty_0_115; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8204 = ~quene ? _GEN_6276 : dirty_0_116; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8205 = ~quene ? _GEN_6277 : dirty_0_117; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8206 = ~quene ? _GEN_6278 : dirty_0_118; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8207 = ~quene ? _GEN_6279 : dirty_0_119; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8208 = ~quene ? _GEN_6280 : dirty_0_120; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8209 = ~quene ? _GEN_6281 : dirty_0_121; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8210 = ~quene ? _GEN_6282 : dirty_0_122; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8211 = ~quene ? _GEN_6283 : dirty_0_123; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8212 = ~quene ? _GEN_6284 : dirty_0_124; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8213 = ~quene ? _GEN_6285 : dirty_0_125; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8214 = ~quene ? _GEN_6286 : dirty_0_126; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8215 = ~quene ? _GEN_6287 : dirty_0_127; // @[d_cache.scala 163:34 32:26]
  wire  _GEN_8216 = ~quene ? _GEN_6288 : valid_0_0; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8217 = ~quene ? _GEN_6289 : valid_0_1; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8218 = ~quene ? _GEN_6290 : valid_0_2; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8219 = ~quene ? _GEN_6291 : valid_0_3; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8220 = ~quene ? _GEN_6292 : valid_0_4; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8221 = ~quene ? _GEN_6293 : valid_0_5; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8222 = ~quene ? _GEN_6294 : valid_0_6; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8223 = ~quene ? _GEN_6295 : valid_0_7; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8224 = ~quene ? _GEN_6296 : valid_0_8; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8225 = ~quene ? _GEN_6297 : valid_0_9; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8226 = ~quene ? _GEN_6298 : valid_0_10; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8227 = ~quene ? _GEN_6299 : valid_0_11; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8228 = ~quene ? _GEN_6300 : valid_0_12; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8229 = ~quene ? _GEN_6301 : valid_0_13; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8230 = ~quene ? _GEN_6302 : valid_0_14; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8231 = ~quene ? _GEN_6303 : valid_0_15; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8232 = ~quene ? _GEN_6304 : valid_0_16; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8233 = ~quene ? _GEN_6305 : valid_0_17; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8234 = ~quene ? _GEN_6306 : valid_0_18; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8235 = ~quene ? _GEN_6307 : valid_0_19; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8236 = ~quene ? _GEN_6308 : valid_0_20; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8237 = ~quene ? _GEN_6309 : valid_0_21; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8238 = ~quene ? _GEN_6310 : valid_0_22; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8239 = ~quene ? _GEN_6311 : valid_0_23; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8240 = ~quene ? _GEN_6312 : valid_0_24; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8241 = ~quene ? _GEN_6313 : valid_0_25; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8242 = ~quene ? _GEN_6314 : valid_0_26; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8243 = ~quene ? _GEN_6315 : valid_0_27; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8244 = ~quene ? _GEN_6316 : valid_0_28; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8245 = ~quene ? _GEN_6317 : valid_0_29; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8246 = ~quene ? _GEN_6318 : valid_0_30; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8247 = ~quene ? _GEN_6319 : valid_0_31; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8248 = ~quene ? _GEN_6320 : valid_0_32; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8249 = ~quene ? _GEN_6321 : valid_0_33; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8250 = ~quene ? _GEN_6322 : valid_0_34; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8251 = ~quene ? _GEN_6323 : valid_0_35; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8252 = ~quene ? _GEN_6324 : valid_0_36; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8253 = ~quene ? _GEN_6325 : valid_0_37; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8254 = ~quene ? _GEN_6326 : valid_0_38; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8255 = ~quene ? _GEN_6327 : valid_0_39; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8256 = ~quene ? _GEN_6328 : valid_0_40; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8257 = ~quene ? _GEN_6329 : valid_0_41; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8258 = ~quene ? _GEN_6330 : valid_0_42; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8259 = ~quene ? _GEN_6331 : valid_0_43; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8260 = ~quene ? _GEN_6332 : valid_0_44; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8261 = ~quene ? _GEN_6333 : valid_0_45; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8262 = ~quene ? _GEN_6334 : valid_0_46; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8263 = ~quene ? _GEN_6335 : valid_0_47; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8264 = ~quene ? _GEN_6336 : valid_0_48; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8265 = ~quene ? _GEN_6337 : valid_0_49; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8266 = ~quene ? _GEN_6338 : valid_0_50; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8267 = ~quene ? _GEN_6339 : valid_0_51; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8268 = ~quene ? _GEN_6340 : valid_0_52; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8269 = ~quene ? _GEN_6341 : valid_0_53; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8270 = ~quene ? _GEN_6342 : valid_0_54; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8271 = ~quene ? _GEN_6343 : valid_0_55; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8272 = ~quene ? _GEN_6344 : valid_0_56; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8273 = ~quene ? _GEN_6345 : valid_0_57; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8274 = ~quene ? _GEN_6346 : valid_0_58; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8275 = ~quene ? _GEN_6347 : valid_0_59; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8276 = ~quene ? _GEN_6348 : valid_0_60; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8277 = ~quene ? _GEN_6349 : valid_0_61; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8278 = ~quene ? _GEN_6350 : valid_0_62; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8279 = ~quene ? _GEN_6351 : valid_0_63; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8280 = ~quene ? _GEN_6352 : valid_0_64; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8281 = ~quene ? _GEN_6353 : valid_0_65; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8282 = ~quene ? _GEN_6354 : valid_0_66; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8283 = ~quene ? _GEN_6355 : valid_0_67; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8284 = ~quene ? _GEN_6356 : valid_0_68; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8285 = ~quene ? _GEN_6357 : valid_0_69; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8286 = ~quene ? _GEN_6358 : valid_0_70; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8287 = ~quene ? _GEN_6359 : valid_0_71; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8288 = ~quene ? _GEN_6360 : valid_0_72; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8289 = ~quene ? _GEN_6361 : valid_0_73; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8290 = ~quene ? _GEN_6362 : valid_0_74; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8291 = ~quene ? _GEN_6363 : valid_0_75; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8292 = ~quene ? _GEN_6364 : valid_0_76; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8293 = ~quene ? _GEN_6365 : valid_0_77; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8294 = ~quene ? _GEN_6366 : valid_0_78; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8295 = ~quene ? _GEN_6367 : valid_0_79; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8296 = ~quene ? _GEN_6368 : valid_0_80; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8297 = ~quene ? _GEN_6369 : valid_0_81; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8298 = ~quene ? _GEN_6370 : valid_0_82; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8299 = ~quene ? _GEN_6371 : valid_0_83; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8300 = ~quene ? _GEN_6372 : valid_0_84; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8301 = ~quene ? _GEN_6373 : valid_0_85; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8302 = ~quene ? _GEN_6374 : valid_0_86; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8303 = ~quene ? _GEN_6375 : valid_0_87; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8304 = ~quene ? _GEN_6376 : valid_0_88; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8305 = ~quene ? _GEN_6377 : valid_0_89; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8306 = ~quene ? _GEN_6378 : valid_0_90; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8307 = ~quene ? _GEN_6379 : valid_0_91; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8308 = ~quene ? _GEN_6380 : valid_0_92; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8309 = ~quene ? _GEN_6381 : valid_0_93; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8310 = ~quene ? _GEN_6382 : valid_0_94; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8311 = ~quene ? _GEN_6383 : valid_0_95; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8312 = ~quene ? _GEN_6384 : valid_0_96; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8313 = ~quene ? _GEN_6385 : valid_0_97; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8314 = ~quene ? _GEN_6386 : valid_0_98; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8315 = ~quene ? _GEN_6387 : valid_0_99; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8316 = ~quene ? _GEN_6388 : valid_0_100; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8317 = ~quene ? _GEN_6389 : valid_0_101; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8318 = ~quene ? _GEN_6390 : valid_0_102; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8319 = ~quene ? _GEN_6391 : valid_0_103; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8320 = ~quene ? _GEN_6392 : valid_0_104; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8321 = ~quene ? _GEN_6393 : valid_0_105; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8322 = ~quene ? _GEN_6394 : valid_0_106; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8323 = ~quene ? _GEN_6395 : valid_0_107; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8324 = ~quene ? _GEN_6396 : valid_0_108; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8325 = ~quene ? _GEN_6397 : valid_0_109; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8326 = ~quene ? _GEN_6398 : valid_0_110; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8327 = ~quene ? _GEN_6399 : valid_0_111; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8328 = ~quene ? _GEN_6400 : valid_0_112; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8329 = ~quene ? _GEN_6401 : valid_0_113; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8330 = ~quene ? _GEN_6402 : valid_0_114; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8331 = ~quene ? _GEN_6403 : valid_0_115; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8332 = ~quene ? _GEN_6404 : valid_0_116; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8333 = ~quene ? _GEN_6405 : valid_0_117; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8334 = ~quene ? _GEN_6406 : valid_0_118; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8335 = ~quene ? _GEN_6407 : valid_0_119; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8336 = ~quene ? _GEN_6408 : valid_0_120; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8337 = ~quene ? _GEN_6409 : valid_0_121; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8338 = ~quene ? _GEN_6410 : valid_0_122; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8339 = ~quene ? _GEN_6411 : valid_0_123; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8340 = ~quene ? _GEN_6412 : valid_0_124; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8341 = ~quene ? _GEN_6413 : valid_0_125; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8342 = ~quene ? _GEN_6414 : valid_0_126; // @[d_cache.scala 163:34 30:26]
  wire  _GEN_8343 = ~quene ? _GEN_6415 : valid_0_127; // @[d_cache.scala 163:34 30:26]
  wire [2:0] _GEN_8344 = ~quene ? _GEN_6416 : _GEN_7828; // @[d_cache.scala 163:34]
  wire [63:0] _GEN_8346 = ~quene ? ram_1_0 : _GEN_7316; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8347 = ~quene ? ram_1_1 : _GEN_7317; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8348 = ~quene ? ram_1_2 : _GEN_7318; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8349 = ~quene ? ram_1_3 : _GEN_7319; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8350 = ~quene ? ram_1_4 : _GEN_7320; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8351 = ~quene ? ram_1_5 : _GEN_7321; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8352 = ~quene ? ram_1_6 : _GEN_7322; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8353 = ~quene ? ram_1_7 : _GEN_7323; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8354 = ~quene ? ram_1_8 : _GEN_7324; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8355 = ~quene ? ram_1_9 : _GEN_7325; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8356 = ~quene ? ram_1_10 : _GEN_7326; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8357 = ~quene ? ram_1_11 : _GEN_7327; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8358 = ~quene ? ram_1_12 : _GEN_7328; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8359 = ~quene ? ram_1_13 : _GEN_7329; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8360 = ~quene ? ram_1_14 : _GEN_7330; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8361 = ~quene ? ram_1_15 : _GEN_7331; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8362 = ~quene ? ram_1_16 : _GEN_7332; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8363 = ~quene ? ram_1_17 : _GEN_7333; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8364 = ~quene ? ram_1_18 : _GEN_7334; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8365 = ~quene ? ram_1_19 : _GEN_7335; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8366 = ~quene ? ram_1_20 : _GEN_7336; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8367 = ~quene ? ram_1_21 : _GEN_7337; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8368 = ~quene ? ram_1_22 : _GEN_7338; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8369 = ~quene ? ram_1_23 : _GEN_7339; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8370 = ~quene ? ram_1_24 : _GEN_7340; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8371 = ~quene ? ram_1_25 : _GEN_7341; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8372 = ~quene ? ram_1_26 : _GEN_7342; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8373 = ~quene ? ram_1_27 : _GEN_7343; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8374 = ~quene ? ram_1_28 : _GEN_7344; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8375 = ~quene ? ram_1_29 : _GEN_7345; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8376 = ~quene ? ram_1_30 : _GEN_7346; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8377 = ~quene ? ram_1_31 : _GEN_7347; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8378 = ~quene ? ram_1_32 : _GEN_7348; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8379 = ~quene ? ram_1_33 : _GEN_7349; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8380 = ~quene ? ram_1_34 : _GEN_7350; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8381 = ~quene ? ram_1_35 : _GEN_7351; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8382 = ~quene ? ram_1_36 : _GEN_7352; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8383 = ~quene ? ram_1_37 : _GEN_7353; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8384 = ~quene ? ram_1_38 : _GEN_7354; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8385 = ~quene ? ram_1_39 : _GEN_7355; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8386 = ~quene ? ram_1_40 : _GEN_7356; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8387 = ~quene ? ram_1_41 : _GEN_7357; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8388 = ~quene ? ram_1_42 : _GEN_7358; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8389 = ~quene ? ram_1_43 : _GEN_7359; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8390 = ~quene ? ram_1_44 : _GEN_7360; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8391 = ~quene ? ram_1_45 : _GEN_7361; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8392 = ~quene ? ram_1_46 : _GEN_7362; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8393 = ~quene ? ram_1_47 : _GEN_7363; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8394 = ~quene ? ram_1_48 : _GEN_7364; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8395 = ~quene ? ram_1_49 : _GEN_7365; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8396 = ~quene ? ram_1_50 : _GEN_7366; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8397 = ~quene ? ram_1_51 : _GEN_7367; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8398 = ~quene ? ram_1_52 : _GEN_7368; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8399 = ~quene ? ram_1_53 : _GEN_7369; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8400 = ~quene ? ram_1_54 : _GEN_7370; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8401 = ~quene ? ram_1_55 : _GEN_7371; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8402 = ~quene ? ram_1_56 : _GEN_7372; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8403 = ~quene ? ram_1_57 : _GEN_7373; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8404 = ~quene ? ram_1_58 : _GEN_7374; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8405 = ~quene ? ram_1_59 : _GEN_7375; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8406 = ~quene ? ram_1_60 : _GEN_7376; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8407 = ~quene ? ram_1_61 : _GEN_7377; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8408 = ~quene ? ram_1_62 : _GEN_7378; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8409 = ~quene ? ram_1_63 : _GEN_7379; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8410 = ~quene ? ram_1_64 : _GEN_7380; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8411 = ~quene ? ram_1_65 : _GEN_7381; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8412 = ~quene ? ram_1_66 : _GEN_7382; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8413 = ~quene ? ram_1_67 : _GEN_7383; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8414 = ~quene ? ram_1_68 : _GEN_7384; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8415 = ~quene ? ram_1_69 : _GEN_7385; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8416 = ~quene ? ram_1_70 : _GEN_7386; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8417 = ~quene ? ram_1_71 : _GEN_7387; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8418 = ~quene ? ram_1_72 : _GEN_7388; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8419 = ~quene ? ram_1_73 : _GEN_7389; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8420 = ~quene ? ram_1_74 : _GEN_7390; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8421 = ~quene ? ram_1_75 : _GEN_7391; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8422 = ~quene ? ram_1_76 : _GEN_7392; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8423 = ~quene ? ram_1_77 : _GEN_7393; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8424 = ~quene ? ram_1_78 : _GEN_7394; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8425 = ~quene ? ram_1_79 : _GEN_7395; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8426 = ~quene ? ram_1_80 : _GEN_7396; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8427 = ~quene ? ram_1_81 : _GEN_7397; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8428 = ~quene ? ram_1_82 : _GEN_7398; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8429 = ~quene ? ram_1_83 : _GEN_7399; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8430 = ~quene ? ram_1_84 : _GEN_7400; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8431 = ~quene ? ram_1_85 : _GEN_7401; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8432 = ~quene ? ram_1_86 : _GEN_7402; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8433 = ~quene ? ram_1_87 : _GEN_7403; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8434 = ~quene ? ram_1_88 : _GEN_7404; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8435 = ~quene ? ram_1_89 : _GEN_7405; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8436 = ~quene ? ram_1_90 : _GEN_7406; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8437 = ~quene ? ram_1_91 : _GEN_7407; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8438 = ~quene ? ram_1_92 : _GEN_7408; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8439 = ~quene ? ram_1_93 : _GEN_7409; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8440 = ~quene ? ram_1_94 : _GEN_7410; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8441 = ~quene ? ram_1_95 : _GEN_7411; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8442 = ~quene ? ram_1_96 : _GEN_7412; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8443 = ~quene ? ram_1_97 : _GEN_7413; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8444 = ~quene ? ram_1_98 : _GEN_7414; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8445 = ~quene ? ram_1_99 : _GEN_7415; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8446 = ~quene ? ram_1_100 : _GEN_7416; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8447 = ~quene ? ram_1_101 : _GEN_7417; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8448 = ~quene ? ram_1_102 : _GEN_7418; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8449 = ~quene ? ram_1_103 : _GEN_7419; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8450 = ~quene ? ram_1_104 : _GEN_7420; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8451 = ~quene ? ram_1_105 : _GEN_7421; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8452 = ~quene ? ram_1_106 : _GEN_7422; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8453 = ~quene ? ram_1_107 : _GEN_7423; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8454 = ~quene ? ram_1_108 : _GEN_7424; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8455 = ~quene ? ram_1_109 : _GEN_7425; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8456 = ~quene ? ram_1_110 : _GEN_7426; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8457 = ~quene ? ram_1_111 : _GEN_7427; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8458 = ~quene ? ram_1_112 : _GEN_7428; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8459 = ~quene ? ram_1_113 : _GEN_7429; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8460 = ~quene ? ram_1_114 : _GEN_7430; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8461 = ~quene ? ram_1_115 : _GEN_7431; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8462 = ~quene ? ram_1_116 : _GEN_7432; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8463 = ~quene ? ram_1_117 : _GEN_7433; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8464 = ~quene ? ram_1_118 : _GEN_7434; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8465 = ~quene ? ram_1_119 : _GEN_7435; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8466 = ~quene ? ram_1_120 : _GEN_7436; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8467 = ~quene ? ram_1_121 : _GEN_7437; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8468 = ~quene ? ram_1_122 : _GEN_7438; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8469 = ~quene ? ram_1_123 : _GEN_7439; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8470 = ~quene ? ram_1_124 : _GEN_7440; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8471 = ~quene ? ram_1_125 : _GEN_7441; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8472 = ~quene ? ram_1_126 : _GEN_7442; // @[d_cache.scala 163:34 20:24]
  wire [63:0] _GEN_8473 = ~quene ? ram_1_127 : _GEN_7443; // @[d_cache.scala 163:34 20:24]
  wire [31:0] _GEN_8474 = ~quene ? tag_1_0 : _GEN_7444; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8475 = ~quene ? tag_1_1 : _GEN_7445; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8476 = ~quene ? tag_1_2 : _GEN_7446; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8477 = ~quene ? tag_1_3 : _GEN_7447; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8478 = ~quene ? tag_1_4 : _GEN_7448; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8479 = ~quene ? tag_1_5 : _GEN_7449; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8480 = ~quene ? tag_1_6 : _GEN_7450; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8481 = ~quene ? tag_1_7 : _GEN_7451; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8482 = ~quene ? tag_1_8 : _GEN_7452; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8483 = ~quene ? tag_1_9 : _GEN_7453; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8484 = ~quene ? tag_1_10 : _GEN_7454; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8485 = ~quene ? tag_1_11 : _GEN_7455; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8486 = ~quene ? tag_1_12 : _GEN_7456; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8487 = ~quene ? tag_1_13 : _GEN_7457; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8488 = ~quene ? tag_1_14 : _GEN_7458; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8489 = ~quene ? tag_1_15 : _GEN_7459; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8490 = ~quene ? tag_1_16 : _GEN_7460; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8491 = ~quene ? tag_1_17 : _GEN_7461; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8492 = ~quene ? tag_1_18 : _GEN_7462; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8493 = ~quene ? tag_1_19 : _GEN_7463; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8494 = ~quene ? tag_1_20 : _GEN_7464; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8495 = ~quene ? tag_1_21 : _GEN_7465; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8496 = ~quene ? tag_1_22 : _GEN_7466; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8497 = ~quene ? tag_1_23 : _GEN_7467; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8498 = ~quene ? tag_1_24 : _GEN_7468; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8499 = ~quene ? tag_1_25 : _GEN_7469; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8500 = ~quene ? tag_1_26 : _GEN_7470; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8501 = ~quene ? tag_1_27 : _GEN_7471; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8502 = ~quene ? tag_1_28 : _GEN_7472; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8503 = ~quene ? tag_1_29 : _GEN_7473; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8504 = ~quene ? tag_1_30 : _GEN_7474; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8505 = ~quene ? tag_1_31 : _GEN_7475; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8506 = ~quene ? tag_1_32 : _GEN_7476; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8507 = ~quene ? tag_1_33 : _GEN_7477; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8508 = ~quene ? tag_1_34 : _GEN_7478; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8509 = ~quene ? tag_1_35 : _GEN_7479; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8510 = ~quene ? tag_1_36 : _GEN_7480; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8511 = ~quene ? tag_1_37 : _GEN_7481; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8512 = ~quene ? tag_1_38 : _GEN_7482; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8513 = ~quene ? tag_1_39 : _GEN_7483; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8514 = ~quene ? tag_1_40 : _GEN_7484; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8515 = ~quene ? tag_1_41 : _GEN_7485; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8516 = ~quene ? tag_1_42 : _GEN_7486; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8517 = ~quene ? tag_1_43 : _GEN_7487; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8518 = ~quene ? tag_1_44 : _GEN_7488; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8519 = ~quene ? tag_1_45 : _GEN_7489; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8520 = ~quene ? tag_1_46 : _GEN_7490; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8521 = ~quene ? tag_1_47 : _GEN_7491; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8522 = ~quene ? tag_1_48 : _GEN_7492; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8523 = ~quene ? tag_1_49 : _GEN_7493; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8524 = ~quene ? tag_1_50 : _GEN_7494; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8525 = ~quene ? tag_1_51 : _GEN_7495; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8526 = ~quene ? tag_1_52 : _GEN_7496; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8527 = ~quene ? tag_1_53 : _GEN_7497; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8528 = ~quene ? tag_1_54 : _GEN_7498; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8529 = ~quene ? tag_1_55 : _GEN_7499; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8530 = ~quene ? tag_1_56 : _GEN_7500; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8531 = ~quene ? tag_1_57 : _GEN_7501; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8532 = ~quene ? tag_1_58 : _GEN_7502; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8533 = ~quene ? tag_1_59 : _GEN_7503; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8534 = ~quene ? tag_1_60 : _GEN_7504; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8535 = ~quene ? tag_1_61 : _GEN_7505; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8536 = ~quene ? tag_1_62 : _GEN_7506; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8537 = ~quene ? tag_1_63 : _GEN_7507; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8538 = ~quene ? tag_1_64 : _GEN_7508; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8539 = ~quene ? tag_1_65 : _GEN_7509; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8540 = ~quene ? tag_1_66 : _GEN_7510; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8541 = ~quene ? tag_1_67 : _GEN_7511; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8542 = ~quene ? tag_1_68 : _GEN_7512; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8543 = ~quene ? tag_1_69 : _GEN_7513; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8544 = ~quene ? tag_1_70 : _GEN_7514; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8545 = ~quene ? tag_1_71 : _GEN_7515; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8546 = ~quene ? tag_1_72 : _GEN_7516; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8547 = ~quene ? tag_1_73 : _GEN_7517; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8548 = ~quene ? tag_1_74 : _GEN_7518; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8549 = ~quene ? tag_1_75 : _GEN_7519; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8550 = ~quene ? tag_1_76 : _GEN_7520; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8551 = ~quene ? tag_1_77 : _GEN_7521; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8552 = ~quene ? tag_1_78 : _GEN_7522; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8553 = ~quene ? tag_1_79 : _GEN_7523; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8554 = ~quene ? tag_1_80 : _GEN_7524; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8555 = ~quene ? tag_1_81 : _GEN_7525; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8556 = ~quene ? tag_1_82 : _GEN_7526; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8557 = ~quene ? tag_1_83 : _GEN_7527; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8558 = ~quene ? tag_1_84 : _GEN_7528; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8559 = ~quene ? tag_1_85 : _GEN_7529; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8560 = ~quene ? tag_1_86 : _GEN_7530; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8561 = ~quene ? tag_1_87 : _GEN_7531; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8562 = ~quene ? tag_1_88 : _GEN_7532; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8563 = ~quene ? tag_1_89 : _GEN_7533; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8564 = ~quene ? tag_1_90 : _GEN_7534; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8565 = ~quene ? tag_1_91 : _GEN_7535; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8566 = ~quene ? tag_1_92 : _GEN_7536; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8567 = ~quene ? tag_1_93 : _GEN_7537; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8568 = ~quene ? tag_1_94 : _GEN_7538; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8569 = ~quene ? tag_1_95 : _GEN_7539; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8570 = ~quene ? tag_1_96 : _GEN_7540; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8571 = ~quene ? tag_1_97 : _GEN_7541; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8572 = ~quene ? tag_1_98 : _GEN_7542; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8573 = ~quene ? tag_1_99 : _GEN_7543; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8574 = ~quene ? tag_1_100 : _GEN_7544; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8575 = ~quene ? tag_1_101 : _GEN_7545; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8576 = ~quene ? tag_1_102 : _GEN_7546; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8577 = ~quene ? tag_1_103 : _GEN_7547; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8578 = ~quene ? tag_1_104 : _GEN_7548; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8579 = ~quene ? tag_1_105 : _GEN_7549; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8580 = ~quene ? tag_1_106 : _GEN_7550; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8581 = ~quene ? tag_1_107 : _GEN_7551; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8582 = ~quene ? tag_1_108 : _GEN_7552; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8583 = ~quene ? tag_1_109 : _GEN_7553; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8584 = ~quene ? tag_1_110 : _GEN_7554; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8585 = ~quene ? tag_1_111 : _GEN_7555; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8586 = ~quene ? tag_1_112 : _GEN_7556; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8587 = ~quene ? tag_1_113 : _GEN_7557; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8588 = ~quene ? tag_1_114 : _GEN_7558; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8589 = ~quene ? tag_1_115 : _GEN_7559; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8590 = ~quene ? tag_1_116 : _GEN_7560; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8591 = ~quene ? tag_1_117 : _GEN_7561; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8592 = ~quene ? tag_1_118 : _GEN_7562; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8593 = ~quene ? tag_1_119 : _GEN_7563; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8594 = ~quene ? tag_1_120 : _GEN_7564; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8595 = ~quene ? tag_1_121 : _GEN_7565; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8596 = ~quene ? tag_1_122 : _GEN_7566; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8597 = ~quene ? tag_1_123 : _GEN_7567; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8598 = ~quene ? tag_1_124 : _GEN_7568; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8599 = ~quene ? tag_1_125 : _GEN_7569; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8600 = ~quene ? tag_1_126 : _GEN_7570; // @[d_cache.scala 163:34 29:24]
  wire [31:0] _GEN_8601 = ~quene ? tag_1_127 : _GEN_7571; // @[d_cache.scala 163:34 29:24]
  wire  _GEN_8602 = ~quene ? dirty_1_0 : _GEN_7572; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8603 = ~quene ? dirty_1_1 : _GEN_7573; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8604 = ~quene ? dirty_1_2 : _GEN_7574; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8605 = ~quene ? dirty_1_3 : _GEN_7575; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8606 = ~quene ? dirty_1_4 : _GEN_7576; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8607 = ~quene ? dirty_1_5 : _GEN_7577; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8608 = ~quene ? dirty_1_6 : _GEN_7578; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8609 = ~quene ? dirty_1_7 : _GEN_7579; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8610 = ~quene ? dirty_1_8 : _GEN_7580; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8611 = ~quene ? dirty_1_9 : _GEN_7581; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8612 = ~quene ? dirty_1_10 : _GEN_7582; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8613 = ~quene ? dirty_1_11 : _GEN_7583; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8614 = ~quene ? dirty_1_12 : _GEN_7584; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8615 = ~quene ? dirty_1_13 : _GEN_7585; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8616 = ~quene ? dirty_1_14 : _GEN_7586; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8617 = ~quene ? dirty_1_15 : _GEN_7587; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8618 = ~quene ? dirty_1_16 : _GEN_7588; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8619 = ~quene ? dirty_1_17 : _GEN_7589; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8620 = ~quene ? dirty_1_18 : _GEN_7590; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8621 = ~quene ? dirty_1_19 : _GEN_7591; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8622 = ~quene ? dirty_1_20 : _GEN_7592; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8623 = ~quene ? dirty_1_21 : _GEN_7593; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8624 = ~quene ? dirty_1_22 : _GEN_7594; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8625 = ~quene ? dirty_1_23 : _GEN_7595; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8626 = ~quene ? dirty_1_24 : _GEN_7596; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8627 = ~quene ? dirty_1_25 : _GEN_7597; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8628 = ~quene ? dirty_1_26 : _GEN_7598; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8629 = ~quene ? dirty_1_27 : _GEN_7599; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8630 = ~quene ? dirty_1_28 : _GEN_7600; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8631 = ~quene ? dirty_1_29 : _GEN_7601; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8632 = ~quene ? dirty_1_30 : _GEN_7602; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8633 = ~quene ? dirty_1_31 : _GEN_7603; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8634 = ~quene ? dirty_1_32 : _GEN_7604; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8635 = ~quene ? dirty_1_33 : _GEN_7605; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8636 = ~quene ? dirty_1_34 : _GEN_7606; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8637 = ~quene ? dirty_1_35 : _GEN_7607; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8638 = ~quene ? dirty_1_36 : _GEN_7608; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8639 = ~quene ? dirty_1_37 : _GEN_7609; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8640 = ~quene ? dirty_1_38 : _GEN_7610; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8641 = ~quene ? dirty_1_39 : _GEN_7611; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8642 = ~quene ? dirty_1_40 : _GEN_7612; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8643 = ~quene ? dirty_1_41 : _GEN_7613; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8644 = ~quene ? dirty_1_42 : _GEN_7614; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8645 = ~quene ? dirty_1_43 : _GEN_7615; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8646 = ~quene ? dirty_1_44 : _GEN_7616; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8647 = ~quene ? dirty_1_45 : _GEN_7617; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8648 = ~quene ? dirty_1_46 : _GEN_7618; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8649 = ~quene ? dirty_1_47 : _GEN_7619; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8650 = ~quene ? dirty_1_48 : _GEN_7620; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8651 = ~quene ? dirty_1_49 : _GEN_7621; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8652 = ~quene ? dirty_1_50 : _GEN_7622; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8653 = ~quene ? dirty_1_51 : _GEN_7623; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8654 = ~quene ? dirty_1_52 : _GEN_7624; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8655 = ~quene ? dirty_1_53 : _GEN_7625; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8656 = ~quene ? dirty_1_54 : _GEN_7626; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8657 = ~quene ? dirty_1_55 : _GEN_7627; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8658 = ~quene ? dirty_1_56 : _GEN_7628; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8659 = ~quene ? dirty_1_57 : _GEN_7629; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8660 = ~quene ? dirty_1_58 : _GEN_7630; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8661 = ~quene ? dirty_1_59 : _GEN_7631; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8662 = ~quene ? dirty_1_60 : _GEN_7632; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8663 = ~quene ? dirty_1_61 : _GEN_7633; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8664 = ~quene ? dirty_1_62 : _GEN_7634; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8665 = ~quene ? dirty_1_63 : _GEN_7635; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8666 = ~quene ? dirty_1_64 : _GEN_7636; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8667 = ~quene ? dirty_1_65 : _GEN_7637; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8668 = ~quene ? dirty_1_66 : _GEN_7638; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8669 = ~quene ? dirty_1_67 : _GEN_7639; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8670 = ~quene ? dirty_1_68 : _GEN_7640; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8671 = ~quene ? dirty_1_69 : _GEN_7641; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8672 = ~quene ? dirty_1_70 : _GEN_7642; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8673 = ~quene ? dirty_1_71 : _GEN_7643; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8674 = ~quene ? dirty_1_72 : _GEN_7644; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8675 = ~quene ? dirty_1_73 : _GEN_7645; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8676 = ~quene ? dirty_1_74 : _GEN_7646; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8677 = ~quene ? dirty_1_75 : _GEN_7647; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8678 = ~quene ? dirty_1_76 : _GEN_7648; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8679 = ~quene ? dirty_1_77 : _GEN_7649; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8680 = ~quene ? dirty_1_78 : _GEN_7650; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8681 = ~quene ? dirty_1_79 : _GEN_7651; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8682 = ~quene ? dirty_1_80 : _GEN_7652; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8683 = ~quene ? dirty_1_81 : _GEN_7653; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8684 = ~quene ? dirty_1_82 : _GEN_7654; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8685 = ~quene ? dirty_1_83 : _GEN_7655; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8686 = ~quene ? dirty_1_84 : _GEN_7656; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8687 = ~quene ? dirty_1_85 : _GEN_7657; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8688 = ~quene ? dirty_1_86 : _GEN_7658; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8689 = ~quene ? dirty_1_87 : _GEN_7659; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8690 = ~quene ? dirty_1_88 : _GEN_7660; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8691 = ~quene ? dirty_1_89 : _GEN_7661; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8692 = ~quene ? dirty_1_90 : _GEN_7662; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8693 = ~quene ? dirty_1_91 : _GEN_7663; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8694 = ~quene ? dirty_1_92 : _GEN_7664; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8695 = ~quene ? dirty_1_93 : _GEN_7665; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8696 = ~quene ? dirty_1_94 : _GEN_7666; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8697 = ~quene ? dirty_1_95 : _GEN_7667; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8698 = ~quene ? dirty_1_96 : _GEN_7668; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8699 = ~quene ? dirty_1_97 : _GEN_7669; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8700 = ~quene ? dirty_1_98 : _GEN_7670; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8701 = ~quene ? dirty_1_99 : _GEN_7671; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8702 = ~quene ? dirty_1_100 : _GEN_7672; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8703 = ~quene ? dirty_1_101 : _GEN_7673; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8704 = ~quene ? dirty_1_102 : _GEN_7674; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8705 = ~quene ? dirty_1_103 : _GEN_7675; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8706 = ~quene ? dirty_1_104 : _GEN_7676; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8707 = ~quene ? dirty_1_105 : _GEN_7677; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8708 = ~quene ? dirty_1_106 : _GEN_7678; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8709 = ~quene ? dirty_1_107 : _GEN_7679; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8710 = ~quene ? dirty_1_108 : _GEN_7680; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8711 = ~quene ? dirty_1_109 : _GEN_7681; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8712 = ~quene ? dirty_1_110 : _GEN_7682; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8713 = ~quene ? dirty_1_111 : _GEN_7683; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8714 = ~quene ? dirty_1_112 : _GEN_7684; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8715 = ~quene ? dirty_1_113 : _GEN_7685; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8716 = ~quene ? dirty_1_114 : _GEN_7686; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8717 = ~quene ? dirty_1_115 : _GEN_7687; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8718 = ~quene ? dirty_1_116 : _GEN_7688; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8719 = ~quene ? dirty_1_117 : _GEN_7689; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8720 = ~quene ? dirty_1_118 : _GEN_7690; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8721 = ~quene ? dirty_1_119 : _GEN_7691; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8722 = ~quene ? dirty_1_120 : _GEN_7692; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8723 = ~quene ? dirty_1_121 : _GEN_7693; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8724 = ~quene ? dirty_1_122 : _GEN_7694; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8725 = ~quene ? dirty_1_123 : _GEN_7695; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8726 = ~quene ? dirty_1_124 : _GEN_7696; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8727 = ~quene ? dirty_1_125 : _GEN_7697; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8728 = ~quene ? dirty_1_126 : _GEN_7698; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8729 = ~quene ? dirty_1_127 : _GEN_7699; // @[d_cache.scala 163:34 33:26]
  wire  _GEN_8730 = ~quene ? valid_1_0 : _GEN_7700; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8731 = ~quene ? valid_1_1 : _GEN_7701; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8732 = ~quene ? valid_1_2 : _GEN_7702; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8733 = ~quene ? valid_1_3 : _GEN_7703; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8734 = ~quene ? valid_1_4 : _GEN_7704; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8735 = ~quene ? valid_1_5 : _GEN_7705; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8736 = ~quene ? valid_1_6 : _GEN_7706; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8737 = ~quene ? valid_1_7 : _GEN_7707; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8738 = ~quene ? valid_1_8 : _GEN_7708; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8739 = ~quene ? valid_1_9 : _GEN_7709; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8740 = ~quene ? valid_1_10 : _GEN_7710; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8741 = ~quene ? valid_1_11 : _GEN_7711; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8742 = ~quene ? valid_1_12 : _GEN_7712; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8743 = ~quene ? valid_1_13 : _GEN_7713; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8744 = ~quene ? valid_1_14 : _GEN_7714; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8745 = ~quene ? valid_1_15 : _GEN_7715; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8746 = ~quene ? valid_1_16 : _GEN_7716; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8747 = ~quene ? valid_1_17 : _GEN_7717; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8748 = ~quene ? valid_1_18 : _GEN_7718; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8749 = ~quene ? valid_1_19 : _GEN_7719; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8750 = ~quene ? valid_1_20 : _GEN_7720; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8751 = ~quene ? valid_1_21 : _GEN_7721; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8752 = ~quene ? valid_1_22 : _GEN_7722; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8753 = ~quene ? valid_1_23 : _GEN_7723; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8754 = ~quene ? valid_1_24 : _GEN_7724; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8755 = ~quene ? valid_1_25 : _GEN_7725; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8756 = ~quene ? valid_1_26 : _GEN_7726; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8757 = ~quene ? valid_1_27 : _GEN_7727; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8758 = ~quene ? valid_1_28 : _GEN_7728; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8759 = ~quene ? valid_1_29 : _GEN_7729; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8760 = ~quene ? valid_1_30 : _GEN_7730; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8761 = ~quene ? valid_1_31 : _GEN_7731; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8762 = ~quene ? valid_1_32 : _GEN_7732; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8763 = ~quene ? valid_1_33 : _GEN_7733; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8764 = ~quene ? valid_1_34 : _GEN_7734; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8765 = ~quene ? valid_1_35 : _GEN_7735; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8766 = ~quene ? valid_1_36 : _GEN_7736; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8767 = ~quene ? valid_1_37 : _GEN_7737; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8768 = ~quene ? valid_1_38 : _GEN_7738; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8769 = ~quene ? valid_1_39 : _GEN_7739; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8770 = ~quene ? valid_1_40 : _GEN_7740; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8771 = ~quene ? valid_1_41 : _GEN_7741; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8772 = ~quene ? valid_1_42 : _GEN_7742; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8773 = ~quene ? valid_1_43 : _GEN_7743; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8774 = ~quene ? valid_1_44 : _GEN_7744; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8775 = ~quene ? valid_1_45 : _GEN_7745; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8776 = ~quene ? valid_1_46 : _GEN_7746; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8777 = ~quene ? valid_1_47 : _GEN_7747; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8778 = ~quene ? valid_1_48 : _GEN_7748; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8779 = ~quene ? valid_1_49 : _GEN_7749; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8780 = ~quene ? valid_1_50 : _GEN_7750; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8781 = ~quene ? valid_1_51 : _GEN_7751; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8782 = ~quene ? valid_1_52 : _GEN_7752; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8783 = ~quene ? valid_1_53 : _GEN_7753; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8784 = ~quene ? valid_1_54 : _GEN_7754; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8785 = ~quene ? valid_1_55 : _GEN_7755; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8786 = ~quene ? valid_1_56 : _GEN_7756; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8787 = ~quene ? valid_1_57 : _GEN_7757; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8788 = ~quene ? valid_1_58 : _GEN_7758; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8789 = ~quene ? valid_1_59 : _GEN_7759; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8790 = ~quene ? valid_1_60 : _GEN_7760; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8791 = ~quene ? valid_1_61 : _GEN_7761; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8792 = ~quene ? valid_1_62 : _GEN_7762; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8793 = ~quene ? valid_1_63 : _GEN_7763; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8794 = ~quene ? valid_1_64 : _GEN_7764; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8795 = ~quene ? valid_1_65 : _GEN_7765; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8796 = ~quene ? valid_1_66 : _GEN_7766; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8797 = ~quene ? valid_1_67 : _GEN_7767; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8798 = ~quene ? valid_1_68 : _GEN_7768; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8799 = ~quene ? valid_1_69 : _GEN_7769; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8800 = ~quene ? valid_1_70 : _GEN_7770; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8801 = ~quene ? valid_1_71 : _GEN_7771; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8802 = ~quene ? valid_1_72 : _GEN_7772; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8803 = ~quene ? valid_1_73 : _GEN_7773; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8804 = ~quene ? valid_1_74 : _GEN_7774; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8805 = ~quene ? valid_1_75 : _GEN_7775; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8806 = ~quene ? valid_1_76 : _GEN_7776; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8807 = ~quene ? valid_1_77 : _GEN_7777; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8808 = ~quene ? valid_1_78 : _GEN_7778; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8809 = ~quene ? valid_1_79 : _GEN_7779; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8810 = ~quene ? valid_1_80 : _GEN_7780; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8811 = ~quene ? valid_1_81 : _GEN_7781; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8812 = ~quene ? valid_1_82 : _GEN_7782; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8813 = ~quene ? valid_1_83 : _GEN_7783; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8814 = ~quene ? valid_1_84 : _GEN_7784; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8815 = ~quene ? valid_1_85 : _GEN_7785; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8816 = ~quene ? valid_1_86 : _GEN_7786; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8817 = ~quene ? valid_1_87 : _GEN_7787; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8818 = ~quene ? valid_1_88 : _GEN_7788; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8819 = ~quene ? valid_1_89 : _GEN_7789; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8820 = ~quene ? valid_1_90 : _GEN_7790; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8821 = ~quene ? valid_1_91 : _GEN_7791; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8822 = ~quene ? valid_1_92 : _GEN_7792; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8823 = ~quene ? valid_1_93 : _GEN_7793; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8824 = ~quene ? valid_1_94 : _GEN_7794; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8825 = ~quene ? valid_1_95 : _GEN_7795; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8826 = ~quene ? valid_1_96 : _GEN_7796; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8827 = ~quene ? valid_1_97 : _GEN_7797; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8828 = ~quene ? valid_1_98 : _GEN_7798; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8829 = ~quene ? valid_1_99 : _GEN_7799; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8830 = ~quene ? valid_1_100 : _GEN_7800; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8831 = ~quene ? valid_1_101 : _GEN_7801; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8832 = ~quene ? valid_1_102 : _GEN_7802; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8833 = ~quene ? valid_1_103 : _GEN_7803; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8834 = ~quene ? valid_1_104 : _GEN_7804; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8835 = ~quene ? valid_1_105 : _GEN_7805; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8836 = ~quene ? valid_1_106 : _GEN_7806; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8837 = ~quene ? valid_1_107 : _GEN_7807; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8838 = ~quene ? valid_1_108 : _GEN_7808; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8839 = ~quene ? valid_1_109 : _GEN_7809; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8840 = ~quene ? valid_1_110 : _GEN_7810; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8841 = ~quene ? valid_1_111 : _GEN_7811; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8842 = ~quene ? valid_1_112 : _GEN_7812; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8843 = ~quene ? valid_1_113 : _GEN_7813; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8844 = ~quene ? valid_1_114 : _GEN_7814; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8845 = ~quene ? valid_1_115 : _GEN_7815; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8846 = ~quene ? valid_1_116 : _GEN_7816; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8847 = ~quene ? valid_1_117 : _GEN_7817; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8848 = ~quene ? valid_1_118 : _GEN_7818; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8849 = ~quene ? valid_1_119 : _GEN_7819; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8850 = ~quene ? valid_1_120 : _GEN_7820; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8851 = ~quene ? valid_1_121 : _GEN_7821; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8852 = ~quene ? valid_1_122 : _GEN_7822; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8853 = ~quene ? valid_1_123 : _GEN_7823; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8854 = ~quene ? valid_1_124 : _GEN_7824; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8855 = ~quene ? valid_1_125 : _GEN_7825; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8856 = ~quene ? valid_1_126 : _GEN_7826; // @[d_cache.scala 163:34 31:26]
  wire  _GEN_8857 = ~quene ? valid_1_127 : _GEN_7827; // @[d_cache.scala 163:34 31:26]
  wire [2:0] _GEN_8858 = unuse_way == 2'h2 ? 3'h7 : _GEN_8344; // @[d_cache.scala 156:40 157:23]
  wire [63:0] _GEN_8859 = unuse_way == 2'h2 ? _GEN_4622 : _GEN_8346; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8860 = unuse_way == 2'h2 ? _GEN_4623 : _GEN_8347; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8861 = unuse_way == 2'h2 ? _GEN_4624 : _GEN_8348; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8862 = unuse_way == 2'h2 ? _GEN_4625 : _GEN_8349; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8863 = unuse_way == 2'h2 ? _GEN_4626 : _GEN_8350; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8864 = unuse_way == 2'h2 ? _GEN_4627 : _GEN_8351; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8865 = unuse_way == 2'h2 ? _GEN_4628 : _GEN_8352; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8866 = unuse_way == 2'h2 ? _GEN_4629 : _GEN_8353; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8867 = unuse_way == 2'h2 ? _GEN_4630 : _GEN_8354; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8868 = unuse_way == 2'h2 ? _GEN_4631 : _GEN_8355; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8869 = unuse_way == 2'h2 ? _GEN_4632 : _GEN_8356; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8870 = unuse_way == 2'h2 ? _GEN_4633 : _GEN_8357; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8871 = unuse_way == 2'h2 ? _GEN_4634 : _GEN_8358; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8872 = unuse_way == 2'h2 ? _GEN_4635 : _GEN_8359; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8873 = unuse_way == 2'h2 ? _GEN_4636 : _GEN_8360; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8874 = unuse_way == 2'h2 ? _GEN_4637 : _GEN_8361; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8875 = unuse_way == 2'h2 ? _GEN_4638 : _GEN_8362; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8876 = unuse_way == 2'h2 ? _GEN_4639 : _GEN_8363; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8877 = unuse_way == 2'h2 ? _GEN_4640 : _GEN_8364; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8878 = unuse_way == 2'h2 ? _GEN_4641 : _GEN_8365; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8879 = unuse_way == 2'h2 ? _GEN_4642 : _GEN_8366; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8880 = unuse_way == 2'h2 ? _GEN_4643 : _GEN_8367; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8881 = unuse_way == 2'h2 ? _GEN_4644 : _GEN_8368; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8882 = unuse_way == 2'h2 ? _GEN_4645 : _GEN_8369; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8883 = unuse_way == 2'h2 ? _GEN_4646 : _GEN_8370; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8884 = unuse_way == 2'h2 ? _GEN_4647 : _GEN_8371; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8885 = unuse_way == 2'h2 ? _GEN_4648 : _GEN_8372; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8886 = unuse_way == 2'h2 ? _GEN_4649 : _GEN_8373; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8887 = unuse_way == 2'h2 ? _GEN_4650 : _GEN_8374; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8888 = unuse_way == 2'h2 ? _GEN_4651 : _GEN_8375; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8889 = unuse_way == 2'h2 ? _GEN_4652 : _GEN_8376; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8890 = unuse_way == 2'h2 ? _GEN_4653 : _GEN_8377; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8891 = unuse_way == 2'h2 ? _GEN_4654 : _GEN_8378; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8892 = unuse_way == 2'h2 ? _GEN_4655 : _GEN_8379; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8893 = unuse_way == 2'h2 ? _GEN_4656 : _GEN_8380; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8894 = unuse_way == 2'h2 ? _GEN_4657 : _GEN_8381; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8895 = unuse_way == 2'h2 ? _GEN_4658 : _GEN_8382; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8896 = unuse_way == 2'h2 ? _GEN_4659 : _GEN_8383; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8897 = unuse_way == 2'h2 ? _GEN_4660 : _GEN_8384; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8898 = unuse_way == 2'h2 ? _GEN_4661 : _GEN_8385; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8899 = unuse_way == 2'h2 ? _GEN_4662 : _GEN_8386; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8900 = unuse_way == 2'h2 ? _GEN_4663 : _GEN_8387; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8901 = unuse_way == 2'h2 ? _GEN_4664 : _GEN_8388; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8902 = unuse_way == 2'h2 ? _GEN_4665 : _GEN_8389; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8903 = unuse_way == 2'h2 ? _GEN_4666 : _GEN_8390; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8904 = unuse_way == 2'h2 ? _GEN_4667 : _GEN_8391; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8905 = unuse_way == 2'h2 ? _GEN_4668 : _GEN_8392; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8906 = unuse_way == 2'h2 ? _GEN_4669 : _GEN_8393; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8907 = unuse_way == 2'h2 ? _GEN_4670 : _GEN_8394; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8908 = unuse_way == 2'h2 ? _GEN_4671 : _GEN_8395; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8909 = unuse_way == 2'h2 ? _GEN_4672 : _GEN_8396; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8910 = unuse_way == 2'h2 ? _GEN_4673 : _GEN_8397; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8911 = unuse_way == 2'h2 ? _GEN_4674 : _GEN_8398; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8912 = unuse_way == 2'h2 ? _GEN_4675 : _GEN_8399; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8913 = unuse_way == 2'h2 ? _GEN_4676 : _GEN_8400; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8914 = unuse_way == 2'h2 ? _GEN_4677 : _GEN_8401; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8915 = unuse_way == 2'h2 ? _GEN_4678 : _GEN_8402; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8916 = unuse_way == 2'h2 ? _GEN_4679 : _GEN_8403; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8917 = unuse_way == 2'h2 ? _GEN_4680 : _GEN_8404; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8918 = unuse_way == 2'h2 ? _GEN_4681 : _GEN_8405; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8919 = unuse_way == 2'h2 ? _GEN_4682 : _GEN_8406; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8920 = unuse_way == 2'h2 ? _GEN_4683 : _GEN_8407; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8921 = unuse_way == 2'h2 ? _GEN_4684 : _GEN_8408; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8922 = unuse_way == 2'h2 ? _GEN_4685 : _GEN_8409; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8923 = unuse_way == 2'h2 ? _GEN_4686 : _GEN_8410; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8924 = unuse_way == 2'h2 ? _GEN_4687 : _GEN_8411; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8925 = unuse_way == 2'h2 ? _GEN_4688 : _GEN_8412; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8926 = unuse_way == 2'h2 ? _GEN_4689 : _GEN_8413; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8927 = unuse_way == 2'h2 ? _GEN_4690 : _GEN_8414; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8928 = unuse_way == 2'h2 ? _GEN_4691 : _GEN_8415; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8929 = unuse_way == 2'h2 ? _GEN_4692 : _GEN_8416; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8930 = unuse_way == 2'h2 ? _GEN_4693 : _GEN_8417; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8931 = unuse_way == 2'h2 ? _GEN_4694 : _GEN_8418; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8932 = unuse_way == 2'h2 ? _GEN_4695 : _GEN_8419; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8933 = unuse_way == 2'h2 ? _GEN_4696 : _GEN_8420; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8934 = unuse_way == 2'h2 ? _GEN_4697 : _GEN_8421; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8935 = unuse_way == 2'h2 ? _GEN_4698 : _GEN_8422; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8936 = unuse_way == 2'h2 ? _GEN_4699 : _GEN_8423; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8937 = unuse_way == 2'h2 ? _GEN_4700 : _GEN_8424; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8938 = unuse_way == 2'h2 ? _GEN_4701 : _GEN_8425; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8939 = unuse_way == 2'h2 ? _GEN_4702 : _GEN_8426; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8940 = unuse_way == 2'h2 ? _GEN_4703 : _GEN_8427; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8941 = unuse_way == 2'h2 ? _GEN_4704 : _GEN_8428; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8942 = unuse_way == 2'h2 ? _GEN_4705 : _GEN_8429; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8943 = unuse_way == 2'h2 ? _GEN_4706 : _GEN_8430; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8944 = unuse_way == 2'h2 ? _GEN_4707 : _GEN_8431; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8945 = unuse_way == 2'h2 ? _GEN_4708 : _GEN_8432; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8946 = unuse_way == 2'h2 ? _GEN_4709 : _GEN_8433; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8947 = unuse_way == 2'h2 ? _GEN_4710 : _GEN_8434; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8948 = unuse_way == 2'h2 ? _GEN_4711 : _GEN_8435; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8949 = unuse_way == 2'h2 ? _GEN_4712 : _GEN_8436; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8950 = unuse_way == 2'h2 ? _GEN_4713 : _GEN_8437; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8951 = unuse_way == 2'h2 ? _GEN_4714 : _GEN_8438; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8952 = unuse_way == 2'h2 ? _GEN_4715 : _GEN_8439; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8953 = unuse_way == 2'h2 ? _GEN_4716 : _GEN_8440; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8954 = unuse_way == 2'h2 ? _GEN_4717 : _GEN_8441; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8955 = unuse_way == 2'h2 ? _GEN_4718 : _GEN_8442; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8956 = unuse_way == 2'h2 ? _GEN_4719 : _GEN_8443; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8957 = unuse_way == 2'h2 ? _GEN_4720 : _GEN_8444; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8958 = unuse_way == 2'h2 ? _GEN_4721 : _GEN_8445; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8959 = unuse_way == 2'h2 ? _GEN_4722 : _GEN_8446; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8960 = unuse_way == 2'h2 ? _GEN_4723 : _GEN_8447; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8961 = unuse_way == 2'h2 ? _GEN_4724 : _GEN_8448; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8962 = unuse_way == 2'h2 ? _GEN_4725 : _GEN_8449; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8963 = unuse_way == 2'h2 ? _GEN_4726 : _GEN_8450; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8964 = unuse_way == 2'h2 ? _GEN_4727 : _GEN_8451; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8965 = unuse_way == 2'h2 ? _GEN_4728 : _GEN_8452; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8966 = unuse_way == 2'h2 ? _GEN_4729 : _GEN_8453; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8967 = unuse_way == 2'h2 ? _GEN_4730 : _GEN_8454; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8968 = unuse_way == 2'h2 ? _GEN_4731 : _GEN_8455; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8969 = unuse_way == 2'h2 ? _GEN_4732 : _GEN_8456; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8970 = unuse_way == 2'h2 ? _GEN_4733 : _GEN_8457; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8971 = unuse_way == 2'h2 ? _GEN_4734 : _GEN_8458; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8972 = unuse_way == 2'h2 ? _GEN_4735 : _GEN_8459; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8973 = unuse_way == 2'h2 ? _GEN_4736 : _GEN_8460; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8974 = unuse_way == 2'h2 ? _GEN_4737 : _GEN_8461; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8975 = unuse_way == 2'h2 ? _GEN_4738 : _GEN_8462; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8976 = unuse_way == 2'h2 ? _GEN_4739 : _GEN_8463; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8977 = unuse_way == 2'h2 ? _GEN_4740 : _GEN_8464; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8978 = unuse_way == 2'h2 ? _GEN_4741 : _GEN_8465; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8979 = unuse_way == 2'h2 ? _GEN_4742 : _GEN_8466; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8980 = unuse_way == 2'h2 ? _GEN_4743 : _GEN_8467; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8981 = unuse_way == 2'h2 ? _GEN_4744 : _GEN_8468; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8982 = unuse_way == 2'h2 ? _GEN_4745 : _GEN_8469; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8983 = unuse_way == 2'h2 ? _GEN_4746 : _GEN_8470; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8984 = unuse_way == 2'h2 ? _GEN_4747 : _GEN_8471; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8985 = unuse_way == 2'h2 ? _GEN_4748 : _GEN_8472; // @[d_cache.scala 156:40]
  wire [63:0] _GEN_8986 = unuse_way == 2'h2 ? _GEN_4749 : _GEN_8473; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8987 = unuse_way == 2'h2 ? _GEN_4750 : _GEN_8474; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8988 = unuse_way == 2'h2 ? _GEN_4751 : _GEN_8475; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8989 = unuse_way == 2'h2 ? _GEN_4752 : _GEN_8476; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8990 = unuse_way == 2'h2 ? _GEN_4753 : _GEN_8477; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8991 = unuse_way == 2'h2 ? _GEN_4754 : _GEN_8478; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8992 = unuse_way == 2'h2 ? _GEN_4755 : _GEN_8479; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8993 = unuse_way == 2'h2 ? _GEN_4756 : _GEN_8480; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8994 = unuse_way == 2'h2 ? _GEN_4757 : _GEN_8481; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8995 = unuse_way == 2'h2 ? _GEN_4758 : _GEN_8482; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8996 = unuse_way == 2'h2 ? _GEN_4759 : _GEN_8483; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8997 = unuse_way == 2'h2 ? _GEN_4760 : _GEN_8484; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8998 = unuse_way == 2'h2 ? _GEN_4761 : _GEN_8485; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_8999 = unuse_way == 2'h2 ? _GEN_4762 : _GEN_8486; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9000 = unuse_way == 2'h2 ? _GEN_4763 : _GEN_8487; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9001 = unuse_way == 2'h2 ? _GEN_4764 : _GEN_8488; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9002 = unuse_way == 2'h2 ? _GEN_4765 : _GEN_8489; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9003 = unuse_way == 2'h2 ? _GEN_4766 : _GEN_8490; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9004 = unuse_way == 2'h2 ? _GEN_4767 : _GEN_8491; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9005 = unuse_way == 2'h2 ? _GEN_4768 : _GEN_8492; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9006 = unuse_way == 2'h2 ? _GEN_4769 : _GEN_8493; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9007 = unuse_way == 2'h2 ? _GEN_4770 : _GEN_8494; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9008 = unuse_way == 2'h2 ? _GEN_4771 : _GEN_8495; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9009 = unuse_way == 2'h2 ? _GEN_4772 : _GEN_8496; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9010 = unuse_way == 2'h2 ? _GEN_4773 : _GEN_8497; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9011 = unuse_way == 2'h2 ? _GEN_4774 : _GEN_8498; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9012 = unuse_way == 2'h2 ? _GEN_4775 : _GEN_8499; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9013 = unuse_way == 2'h2 ? _GEN_4776 : _GEN_8500; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9014 = unuse_way == 2'h2 ? _GEN_4777 : _GEN_8501; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9015 = unuse_way == 2'h2 ? _GEN_4778 : _GEN_8502; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9016 = unuse_way == 2'h2 ? _GEN_4779 : _GEN_8503; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9017 = unuse_way == 2'h2 ? _GEN_4780 : _GEN_8504; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9018 = unuse_way == 2'h2 ? _GEN_4781 : _GEN_8505; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9019 = unuse_way == 2'h2 ? _GEN_4782 : _GEN_8506; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9020 = unuse_way == 2'h2 ? _GEN_4783 : _GEN_8507; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9021 = unuse_way == 2'h2 ? _GEN_4784 : _GEN_8508; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9022 = unuse_way == 2'h2 ? _GEN_4785 : _GEN_8509; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9023 = unuse_way == 2'h2 ? _GEN_4786 : _GEN_8510; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9024 = unuse_way == 2'h2 ? _GEN_4787 : _GEN_8511; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9025 = unuse_way == 2'h2 ? _GEN_4788 : _GEN_8512; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9026 = unuse_way == 2'h2 ? _GEN_4789 : _GEN_8513; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9027 = unuse_way == 2'h2 ? _GEN_4790 : _GEN_8514; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9028 = unuse_way == 2'h2 ? _GEN_4791 : _GEN_8515; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9029 = unuse_way == 2'h2 ? _GEN_4792 : _GEN_8516; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9030 = unuse_way == 2'h2 ? _GEN_4793 : _GEN_8517; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9031 = unuse_way == 2'h2 ? _GEN_4794 : _GEN_8518; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9032 = unuse_way == 2'h2 ? _GEN_4795 : _GEN_8519; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9033 = unuse_way == 2'h2 ? _GEN_4796 : _GEN_8520; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9034 = unuse_way == 2'h2 ? _GEN_4797 : _GEN_8521; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9035 = unuse_way == 2'h2 ? _GEN_4798 : _GEN_8522; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9036 = unuse_way == 2'h2 ? _GEN_4799 : _GEN_8523; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9037 = unuse_way == 2'h2 ? _GEN_4800 : _GEN_8524; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9038 = unuse_way == 2'h2 ? _GEN_4801 : _GEN_8525; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9039 = unuse_way == 2'h2 ? _GEN_4802 : _GEN_8526; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9040 = unuse_way == 2'h2 ? _GEN_4803 : _GEN_8527; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9041 = unuse_way == 2'h2 ? _GEN_4804 : _GEN_8528; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9042 = unuse_way == 2'h2 ? _GEN_4805 : _GEN_8529; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9043 = unuse_way == 2'h2 ? _GEN_4806 : _GEN_8530; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9044 = unuse_way == 2'h2 ? _GEN_4807 : _GEN_8531; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9045 = unuse_way == 2'h2 ? _GEN_4808 : _GEN_8532; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9046 = unuse_way == 2'h2 ? _GEN_4809 : _GEN_8533; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9047 = unuse_way == 2'h2 ? _GEN_4810 : _GEN_8534; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9048 = unuse_way == 2'h2 ? _GEN_4811 : _GEN_8535; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9049 = unuse_way == 2'h2 ? _GEN_4812 : _GEN_8536; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9050 = unuse_way == 2'h2 ? _GEN_4813 : _GEN_8537; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9051 = unuse_way == 2'h2 ? _GEN_4814 : _GEN_8538; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9052 = unuse_way == 2'h2 ? _GEN_4815 : _GEN_8539; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9053 = unuse_way == 2'h2 ? _GEN_4816 : _GEN_8540; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9054 = unuse_way == 2'h2 ? _GEN_4817 : _GEN_8541; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9055 = unuse_way == 2'h2 ? _GEN_4818 : _GEN_8542; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9056 = unuse_way == 2'h2 ? _GEN_4819 : _GEN_8543; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9057 = unuse_way == 2'h2 ? _GEN_4820 : _GEN_8544; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9058 = unuse_way == 2'h2 ? _GEN_4821 : _GEN_8545; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9059 = unuse_way == 2'h2 ? _GEN_4822 : _GEN_8546; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9060 = unuse_way == 2'h2 ? _GEN_4823 : _GEN_8547; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9061 = unuse_way == 2'h2 ? _GEN_4824 : _GEN_8548; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9062 = unuse_way == 2'h2 ? _GEN_4825 : _GEN_8549; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9063 = unuse_way == 2'h2 ? _GEN_4826 : _GEN_8550; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9064 = unuse_way == 2'h2 ? _GEN_4827 : _GEN_8551; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9065 = unuse_way == 2'h2 ? _GEN_4828 : _GEN_8552; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9066 = unuse_way == 2'h2 ? _GEN_4829 : _GEN_8553; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9067 = unuse_way == 2'h2 ? _GEN_4830 : _GEN_8554; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9068 = unuse_way == 2'h2 ? _GEN_4831 : _GEN_8555; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9069 = unuse_way == 2'h2 ? _GEN_4832 : _GEN_8556; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9070 = unuse_way == 2'h2 ? _GEN_4833 : _GEN_8557; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9071 = unuse_way == 2'h2 ? _GEN_4834 : _GEN_8558; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9072 = unuse_way == 2'h2 ? _GEN_4835 : _GEN_8559; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9073 = unuse_way == 2'h2 ? _GEN_4836 : _GEN_8560; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9074 = unuse_way == 2'h2 ? _GEN_4837 : _GEN_8561; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9075 = unuse_way == 2'h2 ? _GEN_4838 : _GEN_8562; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9076 = unuse_way == 2'h2 ? _GEN_4839 : _GEN_8563; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9077 = unuse_way == 2'h2 ? _GEN_4840 : _GEN_8564; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9078 = unuse_way == 2'h2 ? _GEN_4841 : _GEN_8565; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9079 = unuse_way == 2'h2 ? _GEN_4842 : _GEN_8566; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9080 = unuse_way == 2'h2 ? _GEN_4843 : _GEN_8567; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9081 = unuse_way == 2'h2 ? _GEN_4844 : _GEN_8568; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9082 = unuse_way == 2'h2 ? _GEN_4845 : _GEN_8569; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9083 = unuse_way == 2'h2 ? _GEN_4846 : _GEN_8570; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9084 = unuse_way == 2'h2 ? _GEN_4847 : _GEN_8571; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9085 = unuse_way == 2'h2 ? _GEN_4848 : _GEN_8572; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9086 = unuse_way == 2'h2 ? _GEN_4849 : _GEN_8573; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9087 = unuse_way == 2'h2 ? _GEN_4850 : _GEN_8574; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9088 = unuse_way == 2'h2 ? _GEN_4851 : _GEN_8575; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9089 = unuse_way == 2'h2 ? _GEN_4852 : _GEN_8576; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9090 = unuse_way == 2'h2 ? _GEN_4853 : _GEN_8577; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9091 = unuse_way == 2'h2 ? _GEN_4854 : _GEN_8578; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9092 = unuse_way == 2'h2 ? _GEN_4855 : _GEN_8579; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9093 = unuse_way == 2'h2 ? _GEN_4856 : _GEN_8580; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9094 = unuse_way == 2'h2 ? _GEN_4857 : _GEN_8581; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9095 = unuse_way == 2'h2 ? _GEN_4858 : _GEN_8582; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9096 = unuse_way == 2'h2 ? _GEN_4859 : _GEN_8583; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9097 = unuse_way == 2'h2 ? _GEN_4860 : _GEN_8584; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9098 = unuse_way == 2'h2 ? _GEN_4861 : _GEN_8585; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9099 = unuse_way == 2'h2 ? _GEN_4862 : _GEN_8586; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9100 = unuse_way == 2'h2 ? _GEN_4863 : _GEN_8587; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9101 = unuse_way == 2'h2 ? _GEN_4864 : _GEN_8588; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9102 = unuse_way == 2'h2 ? _GEN_4865 : _GEN_8589; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9103 = unuse_way == 2'h2 ? _GEN_4866 : _GEN_8590; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9104 = unuse_way == 2'h2 ? _GEN_4867 : _GEN_8591; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9105 = unuse_way == 2'h2 ? _GEN_4868 : _GEN_8592; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9106 = unuse_way == 2'h2 ? _GEN_4869 : _GEN_8593; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9107 = unuse_way == 2'h2 ? _GEN_4870 : _GEN_8594; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9108 = unuse_way == 2'h2 ? _GEN_4871 : _GEN_8595; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9109 = unuse_way == 2'h2 ? _GEN_4872 : _GEN_8596; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9110 = unuse_way == 2'h2 ? _GEN_4873 : _GEN_8597; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9111 = unuse_way == 2'h2 ? _GEN_4874 : _GEN_8598; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9112 = unuse_way == 2'h2 ? _GEN_4875 : _GEN_8599; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9113 = unuse_way == 2'h2 ? _GEN_4876 : _GEN_8600; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_9114 = unuse_way == 2'h2 ? _GEN_4877 : _GEN_8601; // @[d_cache.scala 156:40]
  wire  _GEN_9115 = unuse_way == 2'h2 ? _GEN_4878 : _GEN_8730; // @[d_cache.scala 156:40]
  wire  _GEN_9116 = unuse_way == 2'h2 ? _GEN_4879 : _GEN_8731; // @[d_cache.scala 156:40]
  wire  _GEN_9117 = unuse_way == 2'h2 ? _GEN_4880 : _GEN_8732; // @[d_cache.scala 156:40]
  wire  _GEN_9118 = unuse_way == 2'h2 ? _GEN_4881 : _GEN_8733; // @[d_cache.scala 156:40]
  wire  _GEN_9119 = unuse_way == 2'h2 ? _GEN_4882 : _GEN_8734; // @[d_cache.scala 156:40]
  wire  _GEN_9120 = unuse_way == 2'h2 ? _GEN_4883 : _GEN_8735; // @[d_cache.scala 156:40]
  wire  _GEN_9121 = unuse_way == 2'h2 ? _GEN_4884 : _GEN_8736; // @[d_cache.scala 156:40]
  wire  _GEN_9122 = unuse_way == 2'h2 ? _GEN_4885 : _GEN_8737; // @[d_cache.scala 156:40]
  wire  _GEN_9123 = unuse_way == 2'h2 ? _GEN_4886 : _GEN_8738; // @[d_cache.scala 156:40]
  wire  _GEN_9124 = unuse_way == 2'h2 ? _GEN_4887 : _GEN_8739; // @[d_cache.scala 156:40]
  wire  _GEN_9125 = unuse_way == 2'h2 ? _GEN_4888 : _GEN_8740; // @[d_cache.scala 156:40]
  wire  _GEN_9126 = unuse_way == 2'h2 ? _GEN_4889 : _GEN_8741; // @[d_cache.scala 156:40]
  wire  _GEN_9127 = unuse_way == 2'h2 ? _GEN_4890 : _GEN_8742; // @[d_cache.scala 156:40]
  wire  _GEN_9128 = unuse_way == 2'h2 ? _GEN_4891 : _GEN_8743; // @[d_cache.scala 156:40]
  wire  _GEN_9129 = unuse_way == 2'h2 ? _GEN_4892 : _GEN_8744; // @[d_cache.scala 156:40]
  wire  _GEN_9130 = unuse_way == 2'h2 ? _GEN_4893 : _GEN_8745; // @[d_cache.scala 156:40]
  wire  _GEN_9131 = unuse_way == 2'h2 ? _GEN_4894 : _GEN_8746; // @[d_cache.scala 156:40]
  wire  _GEN_9132 = unuse_way == 2'h2 ? _GEN_4895 : _GEN_8747; // @[d_cache.scala 156:40]
  wire  _GEN_9133 = unuse_way == 2'h2 ? _GEN_4896 : _GEN_8748; // @[d_cache.scala 156:40]
  wire  _GEN_9134 = unuse_way == 2'h2 ? _GEN_4897 : _GEN_8749; // @[d_cache.scala 156:40]
  wire  _GEN_9135 = unuse_way == 2'h2 ? _GEN_4898 : _GEN_8750; // @[d_cache.scala 156:40]
  wire  _GEN_9136 = unuse_way == 2'h2 ? _GEN_4899 : _GEN_8751; // @[d_cache.scala 156:40]
  wire  _GEN_9137 = unuse_way == 2'h2 ? _GEN_4900 : _GEN_8752; // @[d_cache.scala 156:40]
  wire  _GEN_9138 = unuse_way == 2'h2 ? _GEN_4901 : _GEN_8753; // @[d_cache.scala 156:40]
  wire  _GEN_9139 = unuse_way == 2'h2 ? _GEN_4902 : _GEN_8754; // @[d_cache.scala 156:40]
  wire  _GEN_9140 = unuse_way == 2'h2 ? _GEN_4903 : _GEN_8755; // @[d_cache.scala 156:40]
  wire  _GEN_9141 = unuse_way == 2'h2 ? _GEN_4904 : _GEN_8756; // @[d_cache.scala 156:40]
  wire  _GEN_9142 = unuse_way == 2'h2 ? _GEN_4905 : _GEN_8757; // @[d_cache.scala 156:40]
  wire  _GEN_9143 = unuse_way == 2'h2 ? _GEN_4906 : _GEN_8758; // @[d_cache.scala 156:40]
  wire  _GEN_9144 = unuse_way == 2'h2 ? _GEN_4907 : _GEN_8759; // @[d_cache.scala 156:40]
  wire  _GEN_9145 = unuse_way == 2'h2 ? _GEN_4908 : _GEN_8760; // @[d_cache.scala 156:40]
  wire  _GEN_9146 = unuse_way == 2'h2 ? _GEN_4909 : _GEN_8761; // @[d_cache.scala 156:40]
  wire  _GEN_9147 = unuse_way == 2'h2 ? _GEN_4910 : _GEN_8762; // @[d_cache.scala 156:40]
  wire  _GEN_9148 = unuse_way == 2'h2 ? _GEN_4911 : _GEN_8763; // @[d_cache.scala 156:40]
  wire  _GEN_9149 = unuse_way == 2'h2 ? _GEN_4912 : _GEN_8764; // @[d_cache.scala 156:40]
  wire  _GEN_9150 = unuse_way == 2'h2 ? _GEN_4913 : _GEN_8765; // @[d_cache.scala 156:40]
  wire  _GEN_9151 = unuse_way == 2'h2 ? _GEN_4914 : _GEN_8766; // @[d_cache.scala 156:40]
  wire  _GEN_9152 = unuse_way == 2'h2 ? _GEN_4915 : _GEN_8767; // @[d_cache.scala 156:40]
  wire  _GEN_9153 = unuse_way == 2'h2 ? _GEN_4916 : _GEN_8768; // @[d_cache.scala 156:40]
  wire  _GEN_9154 = unuse_way == 2'h2 ? _GEN_4917 : _GEN_8769; // @[d_cache.scala 156:40]
  wire  _GEN_9155 = unuse_way == 2'h2 ? _GEN_4918 : _GEN_8770; // @[d_cache.scala 156:40]
  wire  _GEN_9156 = unuse_way == 2'h2 ? _GEN_4919 : _GEN_8771; // @[d_cache.scala 156:40]
  wire  _GEN_9157 = unuse_way == 2'h2 ? _GEN_4920 : _GEN_8772; // @[d_cache.scala 156:40]
  wire  _GEN_9158 = unuse_way == 2'h2 ? _GEN_4921 : _GEN_8773; // @[d_cache.scala 156:40]
  wire  _GEN_9159 = unuse_way == 2'h2 ? _GEN_4922 : _GEN_8774; // @[d_cache.scala 156:40]
  wire  _GEN_9160 = unuse_way == 2'h2 ? _GEN_4923 : _GEN_8775; // @[d_cache.scala 156:40]
  wire  _GEN_9161 = unuse_way == 2'h2 ? _GEN_4924 : _GEN_8776; // @[d_cache.scala 156:40]
  wire  _GEN_9162 = unuse_way == 2'h2 ? _GEN_4925 : _GEN_8777; // @[d_cache.scala 156:40]
  wire  _GEN_9163 = unuse_way == 2'h2 ? _GEN_4926 : _GEN_8778; // @[d_cache.scala 156:40]
  wire  _GEN_9164 = unuse_way == 2'h2 ? _GEN_4927 : _GEN_8779; // @[d_cache.scala 156:40]
  wire  _GEN_9165 = unuse_way == 2'h2 ? _GEN_4928 : _GEN_8780; // @[d_cache.scala 156:40]
  wire  _GEN_9166 = unuse_way == 2'h2 ? _GEN_4929 : _GEN_8781; // @[d_cache.scala 156:40]
  wire  _GEN_9167 = unuse_way == 2'h2 ? _GEN_4930 : _GEN_8782; // @[d_cache.scala 156:40]
  wire  _GEN_9168 = unuse_way == 2'h2 ? _GEN_4931 : _GEN_8783; // @[d_cache.scala 156:40]
  wire  _GEN_9169 = unuse_way == 2'h2 ? _GEN_4932 : _GEN_8784; // @[d_cache.scala 156:40]
  wire  _GEN_9170 = unuse_way == 2'h2 ? _GEN_4933 : _GEN_8785; // @[d_cache.scala 156:40]
  wire  _GEN_9171 = unuse_way == 2'h2 ? _GEN_4934 : _GEN_8786; // @[d_cache.scala 156:40]
  wire  _GEN_9172 = unuse_way == 2'h2 ? _GEN_4935 : _GEN_8787; // @[d_cache.scala 156:40]
  wire  _GEN_9173 = unuse_way == 2'h2 ? _GEN_4936 : _GEN_8788; // @[d_cache.scala 156:40]
  wire  _GEN_9174 = unuse_way == 2'h2 ? _GEN_4937 : _GEN_8789; // @[d_cache.scala 156:40]
  wire  _GEN_9175 = unuse_way == 2'h2 ? _GEN_4938 : _GEN_8790; // @[d_cache.scala 156:40]
  wire  _GEN_9176 = unuse_way == 2'h2 ? _GEN_4939 : _GEN_8791; // @[d_cache.scala 156:40]
  wire  _GEN_9177 = unuse_way == 2'h2 ? _GEN_4940 : _GEN_8792; // @[d_cache.scala 156:40]
  wire  _GEN_9178 = unuse_way == 2'h2 ? _GEN_4941 : _GEN_8793; // @[d_cache.scala 156:40]
  wire  _GEN_9179 = unuse_way == 2'h2 ? _GEN_4942 : _GEN_8794; // @[d_cache.scala 156:40]
  wire  _GEN_9180 = unuse_way == 2'h2 ? _GEN_4943 : _GEN_8795; // @[d_cache.scala 156:40]
  wire  _GEN_9181 = unuse_way == 2'h2 ? _GEN_4944 : _GEN_8796; // @[d_cache.scala 156:40]
  wire  _GEN_9182 = unuse_way == 2'h2 ? _GEN_4945 : _GEN_8797; // @[d_cache.scala 156:40]
  wire  _GEN_9183 = unuse_way == 2'h2 ? _GEN_4946 : _GEN_8798; // @[d_cache.scala 156:40]
  wire  _GEN_9184 = unuse_way == 2'h2 ? _GEN_4947 : _GEN_8799; // @[d_cache.scala 156:40]
  wire  _GEN_9185 = unuse_way == 2'h2 ? _GEN_4948 : _GEN_8800; // @[d_cache.scala 156:40]
  wire  _GEN_9186 = unuse_way == 2'h2 ? _GEN_4949 : _GEN_8801; // @[d_cache.scala 156:40]
  wire  _GEN_9187 = unuse_way == 2'h2 ? _GEN_4950 : _GEN_8802; // @[d_cache.scala 156:40]
  wire  _GEN_9188 = unuse_way == 2'h2 ? _GEN_4951 : _GEN_8803; // @[d_cache.scala 156:40]
  wire  _GEN_9189 = unuse_way == 2'h2 ? _GEN_4952 : _GEN_8804; // @[d_cache.scala 156:40]
  wire  _GEN_9190 = unuse_way == 2'h2 ? _GEN_4953 : _GEN_8805; // @[d_cache.scala 156:40]
  wire  _GEN_9191 = unuse_way == 2'h2 ? _GEN_4954 : _GEN_8806; // @[d_cache.scala 156:40]
  wire  _GEN_9192 = unuse_way == 2'h2 ? _GEN_4955 : _GEN_8807; // @[d_cache.scala 156:40]
  wire  _GEN_9193 = unuse_way == 2'h2 ? _GEN_4956 : _GEN_8808; // @[d_cache.scala 156:40]
  wire  _GEN_9194 = unuse_way == 2'h2 ? _GEN_4957 : _GEN_8809; // @[d_cache.scala 156:40]
  wire  _GEN_9195 = unuse_way == 2'h2 ? _GEN_4958 : _GEN_8810; // @[d_cache.scala 156:40]
  wire  _GEN_9196 = unuse_way == 2'h2 ? _GEN_4959 : _GEN_8811; // @[d_cache.scala 156:40]
  wire  _GEN_9197 = unuse_way == 2'h2 ? _GEN_4960 : _GEN_8812; // @[d_cache.scala 156:40]
  wire  _GEN_9198 = unuse_way == 2'h2 ? _GEN_4961 : _GEN_8813; // @[d_cache.scala 156:40]
  wire  _GEN_9199 = unuse_way == 2'h2 ? _GEN_4962 : _GEN_8814; // @[d_cache.scala 156:40]
  wire  _GEN_9200 = unuse_way == 2'h2 ? _GEN_4963 : _GEN_8815; // @[d_cache.scala 156:40]
  wire  _GEN_9201 = unuse_way == 2'h2 ? _GEN_4964 : _GEN_8816; // @[d_cache.scala 156:40]
  wire  _GEN_9202 = unuse_way == 2'h2 ? _GEN_4965 : _GEN_8817; // @[d_cache.scala 156:40]
  wire  _GEN_9203 = unuse_way == 2'h2 ? _GEN_4966 : _GEN_8818; // @[d_cache.scala 156:40]
  wire  _GEN_9204 = unuse_way == 2'h2 ? _GEN_4967 : _GEN_8819; // @[d_cache.scala 156:40]
  wire  _GEN_9205 = unuse_way == 2'h2 ? _GEN_4968 : _GEN_8820; // @[d_cache.scala 156:40]
  wire  _GEN_9206 = unuse_way == 2'h2 ? _GEN_4969 : _GEN_8821; // @[d_cache.scala 156:40]
  wire  _GEN_9207 = unuse_way == 2'h2 ? _GEN_4970 : _GEN_8822; // @[d_cache.scala 156:40]
  wire  _GEN_9208 = unuse_way == 2'h2 ? _GEN_4971 : _GEN_8823; // @[d_cache.scala 156:40]
  wire  _GEN_9209 = unuse_way == 2'h2 ? _GEN_4972 : _GEN_8824; // @[d_cache.scala 156:40]
  wire  _GEN_9210 = unuse_way == 2'h2 ? _GEN_4973 : _GEN_8825; // @[d_cache.scala 156:40]
  wire  _GEN_9211 = unuse_way == 2'h2 ? _GEN_4974 : _GEN_8826; // @[d_cache.scala 156:40]
  wire  _GEN_9212 = unuse_way == 2'h2 ? _GEN_4975 : _GEN_8827; // @[d_cache.scala 156:40]
  wire  _GEN_9213 = unuse_way == 2'h2 ? _GEN_4976 : _GEN_8828; // @[d_cache.scala 156:40]
  wire  _GEN_9214 = unuse_way == 2'h2 ? _GEN_4977 : _GEN_8829; // @[d_cache.scala 156:40]
  wire  _GEN_9215 = unuse_way == 2'h2 ? _GEN_4978 : _GEN_8830; // @[d_cache.scala 156:40]
  wire  _GEN_9216 = unuse_way == 2'h2 ? _GEN_4979 : _GEN_8831; // @[d_cache.scala 156:40]
  wire  _GEN_9217 = unuse_way == 2'h2 ? _GEN_4980 : _GEN_8832; // @[d_cache.scala 156:40]
  wire  _GEN_9218 = unuse_way == 2'h2 ? _GEN_4981 : _GEN_8833; // @[d_cache.scala 156:40]
  wire  _GEN_9219 = unuse_way == 2'h2 ? _GEN_4982 : _GEN_8834; // @[d_cache.scala 156:40]
  wire  _GEN_9220 = unuse_way == 2'h2 ? _GEN_4983 : _GEN_8835; // @[d_cache.scala 156:40]
  wire  _GEN_9221 = unuse_way == 2'h2 ? _GEN_4984 : _GEN_8836; // @[d_cache.scala 156:40]
  wire  _GEN_9222 = unuse_way == 2'h2 ? _GEN_4985 : _GEN_8837; // @[d_cache.scala 156:40]
  wire  _GEN_9223 = unuse_way == 2'h2 ? _GEN_4986 : _GEN_8838; // @[d_cache.scala 156:40]
  wire  _GEN_9224 = unuse_way == 2'h2 ? _GEN_4987 : _GEN_8839; // @[d_cache.scala 156:40]
  wire  _GEN_9225 = unuse_way == 2'h2 ? _GEN_4988 : _GEN_8840; // @[d_cache.scala 156:40]
  wire  _GEN_9226 = unuse_way == 2'h2 ? _GEN_4989 : _GEN_8841; // @[d_cache.scala 156:40]
  wire  _GEN_9227 = unuse_way == 2'h2 ? _GEN_4990 : _GEN_8842; // @[d_cache.scala 156:40]
  wire  _GEN_9228 = unuse_way == 2'h2 ? _GEN_4991 : _GEN_8843; // @[d_cache.scala 156:40]
  wire  _GEN_9229 = unuse_way == 2'h2 ? _GEN_4992 : _GEN_8844; // @[d_cache.scala 156:40]
  wire  _GEN_9230 = unuse_way == 2'h2 ? _GEN_4993 : _GEN_8845; // @[d_cache.scala 156:40]
  wire  _GEN_9231 = unuse_way == 2'h2 ? _GEN_4994 : _GEN_8846; // @[d_cache.scala 156:40]
  wire  _GEN_9232 = unuse_way == 2'h2 ? _GEN_4995 : _GEN_8847; // @[d_cache.scala 156:40]
  wire  _GEN_9233 = unuse_way == 2'h2 ? _GEN_4996 : _GEN_8848; // @[d_cache.scala 156:40]
  wire  _GEN_9234 = unuse_way == 2'h2 ? _GEN_4997 : _GEN_8849; // @[d_cache.scala 156:40]
  wire  _GEN_9235 = unuse_way == 2'h2 ? _GEN_4998 : _GEN_8850; // @[d_cache.scala 156:40]
  wire  _GEN_9236 = unuse_way == 2'h2 ? _GEN_4999 : _GEN_8851; // @[d_cache.scala 156:40]
  wire  _GEN_9237 = unuse_way == 2'h2 ? _GEN_5000 : _GEN_8852; // @[d_cache.scala 156:40]
  wire  _GEN_9238 = unuse_way == 2'h2 ? _GEN_5001 : _GEN_8853; // @[d_cache.scala 156:40]
  wire  _GEN_9239 = unuse_way == 2'h2 ? _GEN_5002 : _GEN_8854; // @[d_cache.scala 156:40]
  wire  _GEN_9240 = unuse_way == 2'h2 ? _GEN_5003 : _GEN_8855; // @[d_cache.scala 156:40]
  wire  _GEN_9241 = unuse_way == 2'h2 ? _GEN_5004 : _GEN_8856; // @[d_cache.scala 156:40]
  wire  _GEN_9242 = unuse_way == 2'h2 ? _GEN_5005 : _GEN_8857; // @[d_cache.scala 156:40]
  wire  _GEN_9243 = unuse_way == 2'h2 ? 1'h0 : _T_26; // @[d_cache.scala 156:40 161:23]
  wire [63:0] _GEN_9244 = unuse_way == 2'h2 ? write_back_data : _GEN_7830; // @[d_cache.scala 156:40 37:34]
  wire [41:0] _GEN_9245 = unuse_way == 2'h2 ? {{10'd0}, write_back_addr} : _GEN_7831; // @[d_cache.scala 156:40 38:34]
  wire [63:0] _GEN_9246 = unuse_way == 2'h2 ? ram_0_0 : _GEN_7832; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9247 = unuse_way == 2'h2 ? ram_0_1 : _GEN_7833; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9248 = unuse_way == 2'h2 ? ram_0_2 : _GEN_7834; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9249 = unuse_way == 2'h2 ? ram_0_3 : _GEN_7835; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9250 = unuse_way == 2'h2 ? ram_0_4 : _GEN_7836; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9251 = unuse_way == 2'h2 ? ram_0_5 : _GEN_7837; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9252 = unuse_way == 2'h2 ? ram_0_6 : _GEN_7838; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9253 = unuse_way == 2'h2 ? ram_0_7 : _GEN_7839; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9254 = unuse_way == 2'h2 ? ram_0_8 : _GEN_7840; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9255 = unuse_way == 2'h2 ? ram_0_9 : _GEN_7841; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9256 = unuse_way == 2'h2 ? ram_0_10 : _GEN_7842; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9257 = unuse_way == 2'h2 ? ram_0_11 : _GEN_7843; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9258 = unuse_way == 2'h2 ? ram_0_12 : _GEN_7844; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9259 = unuse_way == 2'h2 ? ram_0_13 : _GEN_7845; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9260 = unuse_way == 2'h2 ? ram_0_14 : _GEN_7846; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9261 = unuse_way == 2'h2 ? ram_0_15 : _GEN_7847; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9262 = unuse_way == 2'h2 ? ram_0_16 : _GEN_7848; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9263 = unuse_way == 2'h2 ? ram_0_17 : _GEN_7849; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9264 = unuse_way == 2'h2 ? ram_0_18 : _GEN_7850; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9265 = unuse_way == 2'h2 ? ram_0_19 : _GEN_7851; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9266 = unuse_way == 2'h2 ? ram_0_20 : _GEN_7852; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9267 = unuse_way == 2'h2 ? ram_0_21 : _GEN_7853; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9268 = unuse_way == 2'h2 ? ram_0_22 : _GEN_7854; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9269 = unuse_way == 2'h2 ? ram_0_23 : _GEN_7855; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9270 = unuse_way == 2'h2 ? ram_0_24 : _GEN_7856; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9271 = unuse_way == 2'h2 ? ram_0_25 : _GEN_7857; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9272 = unuse_way == 2'h2 ? ram_0_26 : _GEN_7858; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9273 = unuse_way == 2'h2 ? ram_0_27 : _GEN_7859; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9274 = unuse_way == 2'h2 ? ram_0_28 : _GEN_7860; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9275 = unuse_way == 2'h2 ? ram_0_29 : _GEN_7861; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9276 = unuse_way == 2'h2 ? ram_0_30 : _GEN_7862; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9277 = unuse_way == 2'h2 ? ram_0_31 : _GEN_7863; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9278 = unuse_way == 2'h2 ? ram_0_32 : _GEN_7864; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9279 = unuse_way == 2'h2 ? ram_0_33 : _GEN_7865; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9280 = unuse_way == 2'h2 ? ram_0_34 : _GEN_7866; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9281 = unuse_way == 2'h2 ? ram_0_35 : _GEN_7867; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9282 = unuse_way == 2'h2 ? ram_0_36 : _GEN_7868; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9283 = unuse_way == 2'h2 ? ram_0_37 : _GEN_7869; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9284 = unuse_way == 2'h2 ? ram_0_38 : _GEN_7870; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9285 = unuse_way == 2'h2 ? ram_0_39 : _GEN_7871; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9286 = unuse_way == 2'h2 ? ram_0_40 : _GEN_7872; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9287 = unuse_way == 2'h2 ? ram_0_41 : _GEN_7873; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9288 = unuse_way == 2'h2 ? ram_0_42 : _GEN_7874; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9289 = unuse_way == 2'h2 ? ram_0_43 : _GEN_7875; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9290 = unuse_way == 2'h2 ? ram_0_44 : _GEN_7876; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9291 = unuse_way == 2'h2 ? ram_0_45 : _GEN_7877; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9292 = unuse_way == 2'h2 ? ram_0_46 : _GEN_7878; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9293 = unuse_way == 2'h2 ? ram_0_47 : _GEN_7879; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9294 = unuse_way == 2'h2 ? ram_0_48 : _GEN_7880; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9295 = unuse_way == 2'h2 ? ram_0_49 : _GEN_7881; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9296 = unuse_way == 2'h2 ? ram_0_50 : _GEN_7882; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9297 = unuse_way == 2'h2 ? ram_0_51 : _GEN_7883; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9298 = unuse_way == 2'h2 ? ram_0_52 : _GEN_7884; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9299 = unuse_way == 2'h2 ? ram_0_53 : _GEN_7885; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9300 = unuse_way == 2'h2 ? ram_0_54 : _GEN_7886; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9301 = unuse_way == 2'h2 ? ram_0_55 : _GEN_7887; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9302 = unuse_way == 2'h2 ? ram_0_56 : _GEN_7888; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9303 = unuse_way == 2'h2 ? ram_0_57 : _GEN_7889; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9304 = unuse_way == 2'h2 ? ram_0_58 : _GEN_7890; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9305 = unuse_way == 2'h2 ? ram_0_59 : _GEN_7891; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9306 = unuse_way == 2'h2 ? ram_0_60 : _GEN_7892; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9307 = unuse_way == 2'h2 ? ram_0_61 : _GEN_7893; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9308 = unuse_way == 2'h2 ? ram_0_62 : _GEN_7894; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9309 = unuse_way == 2'h2 ? ram_0_63 : _GEN_7895; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9310 = unuse_way == 2'h2 ? ram_0_64 : _GEN_7896; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9311 = unuse_way == 2'h2 ? ram_0_65 : _GEN_7897; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9312 = unuse_way == 2'h2 ? ram_0_66 : _GEN_7898; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9313 = unuse_way == 2'h2 ? ram_0_67 : _GEN_7899; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9314 = unuse_way == 2'h2 ? ram_0_68 : _GEN_7900; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9315 = unuse_way == 2'h2 ? ram_0_69 : _GEN_7901; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9316 = unuse_way == 2'h2 ? ram_0_70 : _GEN_7902; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9317 = unuse_way == 2'h2 ? ram_0_71 : _GEN_7903; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9318 = unuse_way == 2'h2 ? ram_0_72 : _GEN_7904; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9319 = unuse_way == 2'h2 ? ram_0_73 : _GEN_7905; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9320 = unuse_way == 2'h2 ? ram_0_74 : _GEN_7906; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9321 = unuse_way == 2'h2 ? ram_0_75 : _GEN_7907; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9322 = unuse_way == 2'h2 ? ram_0_76 : _GEN_7908; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9323 = unuse_way == 2'h2 ? ram_0_77 : _GEN_7909; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9324 = unuse_way == 2'h2 ? ram_0_78 : _GEN_7910; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9325 = unuse_way == 2'h2 ? ram_0_79 : _GEN_7911; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9326 = unuse_way == 2'h2 ? ram_0_80 : _GEN_7912; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9327 = unuse_way == 2'h2 ? ram_0_81 : _GEN_7913; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9328 = unuse_way == 2'h2 ? ram_0_82 : _GEN_7914; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9329 = unuse_way == 2'h2 ? ram_0_83 : _GEN_7915; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9330 = unuse_way == 2'h2 ? ram_0_84 : _GEN_7916; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9331 = unuse_way == 2'h2 ? ram_0_85 : _GEN_7917; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9332 = unuse_way == 2'h2 ? ram_0_86 : _GEN_7918; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9333 = unuse_way == 2'h2 ? ram_0_87 : _GEN_7919; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9334 = unuse_way == 2'h2 ? ram_0_88 : _GEN_7920; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9335 = unuse_way == 2'h2 ? ram_0_89 : _GEN_7921; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9336 = unuse_way == 2'h2 ? ram_0_90 : _GEN_7922; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9337 = unuse_way == 2'h2 ? ram_0_91 : _GEN_7923; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9338 = unuse_way == 2'h2 ? ram_0_92 : _GEN_7924; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9339 = unuse_way == 2'h2 ? ram_0_93 : _GEN_7925; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9340 = unuse_way == 2'h2 ? ram_0_94 : _GEN_7926; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9341 = unuse_way == 2'h2 ? ram_0_95 : _GEN_7927; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9342 = unuse_way == 2'h2 ? ram_0_96 : _GEN_7928; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9343 = unuse_way == 2'h2 ? ram_0_97 : _GEN_7929; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9344 = unuse_way == 2'h2 ? ram_0_98 : _GEN_7930; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9345 = unuse_way == 2'h2 ? ram_0_99 : _GEN_7931; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9346 = unuse_way == 2'h2 ? ram_0_100 : _GEN_7932; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9347 = unuse_way == 2'h2 ? ram_0_101 : _GEN_7933; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9348 = unuse_way == 2'h2 ? ram_0_102 : _GEN_7934; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9349 = unuse_way == 2'h2 ? ram_0_103 : _GEN_7935; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9350 = unuse_way == 2'h2 ? ram_0_104 : _GEN_7936; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9351 = unuse_way == 2'h2 ? ram_0_105 : _GEN_7937; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9352 = unuse_way == 2'h2 ? ram_0_106 : _GEN_7938; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9353 = unuse_way == 2'h2 ? ram_0_107 : _GEN_7939; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9354 = unuse_way == 2'h2 ? ram_0_108 : _GEN_7940; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9355 = unuse_way == 2'h2 ? ram_0_109 : _GEN_7941; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9356 = unuse_way == 2'h2 ? ram_0_110 : _GEN_7942; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9357 = unuse_way == 2'h2 ? ram_0_111 : _GEN_7943; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9358 = unuse_way == 2'h2 ? ram_0_112 : _GEN_7944; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9359 = unuse_way == 2'h2 ? ram_0_113 : _GEN_7945; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9360 = unuse_way == 2'h2 ? ram_0_114 : _GEN_7946; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9361 = unuse_way == 2'h2 ? ram_0_115 : _GEN_7947; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9362 = unuse_way == 2'h2 ? ram_0_116 : _GEN_7948; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9363 = unuse_way == 2'h2 ? ram_0_117 : _GEN_7949; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9364 = unuse_way == 2'h2 ? ram_0_118 : _GEN_7950; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9365 = unuse_way == 2'h2 ? ram_0_119 : _GEN_7951; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9366 = unuse_way == 2'h2 ? ram_0_120 : _GEN_7952; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9367 = unuse_way == 2'h2 ? ram_0_121 : _GEN_7953; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9368 = unuse_way == 2'h2 ? ram_0_122 : _GEN_7954; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9369 = unuse_way == 2'h2 ? ram_0_123 : _GEN_7955; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9370 = unuse_way == 2'h2 ? ram_0_124 : _GEN_7956; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9371 = unuse_way == 2'h2 ? ram_0_125 : _GEN_7957; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9372 = unuse_way == 2'h2 ? ram_0_126 : _GEN_7958; // @[d_cache.scala 156:40 19:24]
  wire [63:0] _GEN_9373 = unuse_way == 2'h2 ? ram_0_127 : _GEN_7959; // @[d_cache.scala 156:40 19:24]
  wire [31:0] _GEN_9374 = unuse_way == 2'h2 ? tag_0_0 : _GEN_7960; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9375 = unuse_way == 2'h2 ? tag_0_1 : _GEN_7961; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9376 = unuse_way == 2'h2 ? tag_0_2 : _GEN_7962; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9377 = unuse_way == 2'h2 ? tag_0_3 : _GEN_7963; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9378 = unuse_way == 2'h2 ? tag_0_4 : _GEN_7964; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9379 = unuse_way == 2'h2 ? tag_0_5 : _GEN_7965; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9380 = unuse_way == 2'h2 ? tag_0_6 : _GEN_7966; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9381 = unuse_way == 2'h2 ? tag_0_7 : _GEN_7967; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9382 = unuse_way == 2'h2 ? tag_0_8 : _GEN_7968; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9383 = unuse_way == 2'h2 ? tag_0_9 : _GEN_7969; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9384 = unuse_way == 2'h2 ? tag_0_10 : _GEN_7970; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9385 = unuse_way == 2'h2 ? tag_0_11 : _GEN_7971; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9386 = unuse_way == 2'h2 ? tag_0_12 : _GEN_7972; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9387 = unuse_way == 2'h2 ? tag_0_13 : _GEN_7973; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9388 = unuse_way == 2'h2 ? tag_0_14 : _GEN_7974; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9389 = unuse_way == 2'h2 ? tag_0_15 : _GEN_7975; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9390 = unuse_way == 2'h2 ? tag_0_16 : _GEN_7976; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9391 = unuse_way == 2'h2 ? tag_0_17 : _GEN_7977; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9392 = unuse_way == 2'h2 ? tag_0_18 : _GEN_7978; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9393 = unuse_way == 2'h2 ? tag_0_19 : _GEN_7979; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9394 = unuse_way == 2'h2 ? tag_0_20 : _GEN_7980; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9395 = unuse_way == 2'h2 ? tag_0_21 : _GEN_7981; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9396 = unuse_way == 2'h2 ? tag_0_22 : _GEN_7982; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9397 = unuse_way == 2'h2 ? tag_0_23 : _GEN_7983; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9398 = unuse_way == 2'h2 ? tag_0_24 : _GEN_7984; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9399 = unuse_way == 2'h2 ? tag_0_25 : _GEN_7985; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9400 = unuse_way == 2'h2 ? tag_0_26 : _GEN_7986; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9401 = unuse_way == 2'h2 ? tag_0_27 : _GEN_7987; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9402 = unuse_way == 2'h2 ? tag_0_28 : _GEN_7988; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9403 = unuse_way == 2'h2 ? tag_0_29 : _GEN_7989; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9404 = unuse_way == 2'h2 ? tag_0_30 : _GEN_7990; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9405 = unuse_way == 2'h2 ? tag_0_31 : _GEN_7991; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9406 = unuse_way == 2'h2 ? tag_0_32 : _GEN_7992; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9407 = unuse_way == 2'h2 ? tag_0_33 : _GEN_7993; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9408 = unuse_way == 2'h2 ? tag_0_34 : _GEN_7994; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9409 = unuse_way == 2'h2 ? tag_0_35 : _GEN_7995; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9410 = unuse_way == 2'h2 ? tag_0_36 : _GEN_7996; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9411 = unuse_way == 2'h2 ? tag_0_37 : _GEN_7997; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9412 = unuse_way == 2'h2 ? tag_0_38 : _GEN_7998; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9413 = unuse_way == 2'h2 ? tag_0_39 : _GEN_7999; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9414 = unuse_way == 2'h2 ? tag_0_40 : _GEN_8000; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9415 = unuse_way == 2'h2 ? tag_0_41 : _GEN_8001; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9416 = unuse_way == 2'h2 ? tag_0_42 : _GEN_8002; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9417 = unuse_way == 2'h2 ? tag_0_43 : _GEN_8003; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9418 = unuse_way == 2'h2 ? tag_0_44 : _GEN_8004; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9419 = unuse_way == 2'h2 ? tag_0_45 : _GEN_8005; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9420 = unuse_way == 2'h2 ? tag_0_46 : _GEN_8006; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9421 = unuse_way == 2'h2 ? tag_0_47 : _GEN_8007; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9422 = unuse_way == 2'h2 ? tag_0_48 : _GEN_8008; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9423 = unuse_way == 2'h2 ? tag_0_49 : _GEN_8009; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9424 = unuse_way == 2'h2 ? tag_0_50 : _GEN_8010; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9425 = unuse_way == 2'h2 ? tag_0_51 : _GEN_8011; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9426 = unuse_way == 2'h2 ? tag_0_52 : _GEN_8012; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9427 = unuse_way == 2'h2 ? tag_0_53 : _GEN_8013; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9428 = unuse_way == 2'h2 ? tag_0_54 : _GEN_8014; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9429 = unuse_way == 2'h2 ? tag_0_55 : _GEN_8015; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9430 = unuse_way == 2'h2 ? tag_0_56 : _GEN_8016; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9431 = unuse_way == 2'h2 ? tag_0_57 : _GEN_8017; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9432 = unuse_way == 2'h2 ? tag_0_58 : _GEN_8018; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9433 = unuse_way == 2'h2 ? tag_0_59 : _GEN_8019; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9434 = unuse_way == 2'h2 ? tag_0_60 : _GEN_8020; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9435 = unuse_way == 2'h2 ? tag_0_61 : _GEN_8021; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9436 = unuse_way == 2'h2 ? tag_0_62 : _GEN_8022; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9437 = unuse_way == 2'h2 ? tag_0_63 : _GEN_8023; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9438 = unuse_way == 2'h2 ? tag_0_64 : _GEN_8024; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9439 = unuse_way == 2'h2 ? tag_0_65 : _GEN_8025; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9440 = unuse_way == 2'h2 ? tag_0_66 : _GEN_8026; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9441 = unuse_way == 2'h2 ? tag_0_67 : _GEN_8027; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9442 = unuse_way == 2'h2 ? tag_0_68 : _GEN_8028; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9443 = unuse_way == 2'h2 ? tag_0_69 : _GEN_8029; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9444 = unuse_way == 2'h2 ? tag_0_70 : _GEN_8030; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9445 = unuse_way == 2'h2 ? tag_0_71 : _GEN_8031; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9446 = unuse_way == 2'h2 ? tag_0_72 : _GEN_8032; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9447 = unuse_way == 2'h2 ? tag_0_73 : _GEN_8033; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9448 = unuse_way == 2'h2 ? tag_0_74 : _GEN_8034; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9449 = unuse_way == 2'h2 ? tag_0_75 : _GEN_8035; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9450 = unuse_way == 2'h2 ? tag_0_76 : _GEN_8036; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9451 = unuse_way == 2'h2 ? tag_0_77 : _GEN_8037; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9452 = unuse_way == 2'h2 ? tag_0_78 : _GEN_8038; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9453 = unuse_way == 2'h2 ? tag_0_79 : _GEN_8039; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9454 = unuse_way == 2'h2 ? tag_0_80 : _GEN_8040; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9455 = unuse_way == 2'h2 ? tag_0_81 : _GEN_8041; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9456 = unuse_way == 2'h2 ? tag_0_82 : _GEN_8042; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9457 = unuse_way == 2'h2 ? tag_0_83 : _GEN_8043; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9458 = unuse_way == 2'h2 ? tag_0_84 : _GEN_8044; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9459 = unuse_way == 2'h2 ? tag_0_85 : _GEN_8045; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9460 = unuse_way == 2'h2 ? tag_0_86 : _GEN_8046; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9461 = unuse_way == 2'h2 ? tag_0_87 : _GEN_8047; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9462 = unuse_way == 2'h2 ? tag_0_88 : _GEN_8048; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9463 = unuse_way == 2'h2 ? tag_0_89 : _GEN_8049; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9464 = unuse_way == 2'h2 ? tag_0_90 : _GEN_8050; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9465 = unuse_way == 2'h2 ? tag_0_91 : _GEN_8051; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9466 = unuse_way == 2'h2 ? tag_0_92 : _GEN_8052; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9467 = unuse_way == 2'h2 ? tag_0_93 : _GEN_8053; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9468 = unuse_way == 2'h2 ? tag_0_94 : _GEN_8054; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9469 = unuse_way == 2'h2 ? tag_0_95 : _GEN_8055; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9470 = unuse_way == 2'h2 ? tag_0_96 : _GEN_8056; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9471 = unuse_way == 2'h2 ? tag_0_97 : _GEN_8057; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9472 = unuse_way == 2'h2 ? tag_0_98 : _GEN_8058; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9473 = unuse_way == 2'h2 ? tag_0_99 : _GEN_8059; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9474 = unuse_way == 2'h2 ? tag_0_100 : _GEN_8060; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9475 = unuse_way == 2'h2 ? tag_0_101 : _GEN_8061; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9476 = unuse_way == 2'h2 ? tag_0_102 : _GEN_8062; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9477 = unuse_way == 2'h2 ? tag_0_103 : _GEN_8063; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9478 = unuse_way == 2'h2 ? tag_0_104 : _GEN_8064; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9479 = unuse_way == 2'h2 ? tag_0_105 : _GEN_8065; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9480 = unuse_way == 2'h2 ? tag_0_106 : _GEN_8066; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9481 = unuse_way == 2'h2 ? tag_0_107 : _GEN_8067; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9482 = unuse_way == 2'h2 ? tag_0_108 : _GEN_8068; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9483 = unuse_way == 2'h2 ? tag_0_109 : _GEN_8069; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9484 = unuse_way == 2'h2 ? tag_0_110 : _GEN_8070; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9485 = unuse_way == 2'h2 ? tag_0_111 : _GEN_8071; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9486 = unuse_way == 2'h2 ? tag_0_112 : _GEN_8072; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9487 = unuse_way == 2'h2 ? tag_0_113 : _GEN_8073; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9488 = unuse_way == 2'h2 ? tag_0_114 : _GEN_8074; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9489 = unuse_way == 2'h2 ? tag_0_115 : _GEN_8075; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9490 = unuse_way == 2'h2 ? tag_0_116 : _GEN_8076; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9491 = unuse_way == 2'h2 ? tag_0_117 : _GEN_8077; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9492 = unuse_way == 2'h2 ? tag_0_118 : _GEN_8078; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9493 = unuse_way == 2'h2 ? tag_0_119 : _GEN_8079; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9494 = unuse_way == 2'h2 ? tag_0_120 : _GEN_8080; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9495 = unuse_way == 2'h2 ? tag_0_121 : _GEN_8081; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9496 = unuse_way == 2'h2 ? tag_0_122 : _GEN_8082; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9497 = unuse_way == 2'h2 ? tag_0_123 : _GEN_8083; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9498 = unuse_way == 2'h2 ? tag_0_124 : _GEN_8084; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9499 = unuse_way == 2'h2 ? tag_0_125 : _GEN_8085; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9500 = unuse_way == 2'h2 ? tag_0_126 : _GEN_8086; // @[d_cache.scala 156:40 28:24]
  wire [31:0] _GEN_9501 = unuse_way == 2'h2 ? tag_0_127 : _GEN_8087; // @[d_cache.scala 156:40 28:24]
  wire  _GEN_9502 = unuse_way == 2'h2 ? dirty_0_0 : _GEN_8088; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9503 = unuse_way == 2'h2 ? dirty_0_1 : _GEN_8089; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9504 = unuse_way == 2'h2 ? dirty_0_2 : _GEN_8090; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9505 = unuse_way == 2'h2 ? dirty_0_3 : _GEN_8091; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9506 = unuse_way == 2'h2 ? dirty_0_4 : _GEN_8092; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9507 = unuse_way == 2'h2 ? dirty_0_5 : _GEN_8093; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9508 = unuse_way == 2'h2 ? dirty_0_6 : _GEN_8094; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9509 = unuse_way == 2'h2 ? dirty_0_7 : _GEN_8095; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9510 = unuse_way == 2'h2 ? dirty_0_8 : _GEN_8096; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9511 = unuse_way == 2'h2 ? dirty_0_9 : _GEN_8097; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9512 = unuse_way == 2'h2 ? dirty_0_10 : _GEN_8098; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9513 = unuse_way == 2'h2 ? dirty_0_11 : _GEN_8099; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9514 = unuse_way == 2'h2 ? dirty_0_12 : _GEN_8100; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9515 = unuse_way == 2'h2 ? dirty_0_13 : _GEN_8101; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9516 = unuse_way == 2'h2 ? dirty_0_14 : _GEN_8102; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9517 = unuse_way == 2'h2 ? dirty_0_15 : _GEN_8103; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9518 = unuse_way == 2'h2 ? dirty_0_16 : _GEN_8104; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9519 = unuse_way == 2'h2 ? dirty_0_17 : _GEN_8105; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9520 = unuse_way == 2'h2 ? dirty_0_18 : _GEN_8106; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9521 = unuse_way == 2'h2 ? dirty_0_19 : _GEN_8107; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9522 = unuse_way == 2'h2 ? dirty_0_20 : _GEN_8108; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9523 = unuse_way == 2'h2 ? dirty_0_21 : _GEN_8109; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9524 = unuse_way == 2'h2 ? dirty_0_22 : _GEN_8110; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9525 = unuse_way == 2'h2 ? dirty_0_23 : _GEN_8111; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9526 = unuse_way == 2'h2 ? dirty_0_24 : _GEN_8112; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9527 = unuse_way == 2'h2 ? dirty_0_25 : _GEN_8113; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9528 = unuse_way == 2'h2 ? dirty_0_26 : _GEN_8114; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9529 = unuse_way == 2'h2 ? dirty_0_27 : _GEN_8115; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9530 = unuse_way == 2'h2 ? dirty_0_28 : _GEN_8116; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9531 = unuse_way == 2'h2 ? dirty_0_29 : _GEN_8117; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9532 = unuse_way == 2'h2 ? dirty_0_30 : _GEN_8118; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9533 = unuse_way == 2'h2 ? dirty_0_31 : _GEN_8119; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9534 = unuse_way == 2'h2 ? dirty_0_32 : _GEN_8120; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9535 = unuse_way == 2'h2 ? dirty_0_33 : _GEN_8121; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9536 = unuse_way == 2'h2 ? dirty_0_34 : _GEN_8122; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9537 = unuse_way == 2'h2 ? dirty_0_35 : _GEN_8123; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9538 = unuse_way == 2'h2 ? dirty_0_36 : _GEN_8124; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9539 = unuse_way == 2'h2 ? dirty_0_37 : _GEN_8125; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9540 = unuse_way == 2'h2 ? dirty_0_38 : _GEN_8126; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9541 = unuse_way == 2'h2 ? dirty_0_39 : _GEN_8127; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9542 = unuse_way == 2'h2 ? dirty_0_40 : _GEN_8128; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9543 = unuse_way == 2'h2 ? dirty_0_41 : _GEN_8129; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9544 = unuse_way == 2'h2 ? dirty_0_42 : _GEN_8130; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9545 = unuse_way == 2'h2 ? dirty_0_43 : _GEN_8131; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9546 = unuse_way == 2'h2 ? dirty_0_44 : _GEN_8132; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9547 = unuse_way == 2'h2 ? dirty_0_45 : _GEN_8133; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9548 = unuse_way == 2'h2 ? dirty_0_46 : _GEN_8134; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9549 = unuse_way == 2'h2 ? dirty_0_47 : _GEN_8135; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9550 = unuse_way == 2'h2 ? dirty_0_48 : _GEN_8136; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9551 = unuse_way == 2'h2 ? dirty_0_49 : _GEN_8137; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9552 = unuse_way == 2'h2 ? dirty_0_50 : _GEN_8138; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9553 = unuse_way == 2'h2 ? dirty_0_51 : _GEN_8139; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9554 = unuse_way == 2'h2 ? dirty_0_52 : _GEN_8140; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9555 = unuse_way == 2'h2 ? dirty_0_53 : _GEN_8141; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9556 = unuse_way == 2'h2 ? dirty_0_54 : _GEN_8142; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9557 = unuse_way == 2'h2 ? dirty_0_55 : _GEN_8143; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9558 = unuse_way == 2'h2 ? dirty_0_56 : _GEN_8144; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9559 = unuse_way == 2'h2 ? dirty_0_57 : _GEN_8145; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9560 = unuse_way == 2'h2 ? dirty_0_58 : _GEN_8146; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9561 = unuse_way == 2'h2 ? dirty_0_59 : _GEN_8147; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9562 = unuse_way == 2'h2 ? dirty_0_60 : _GEN_8148; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9563 = unuse_way == 2'h2 ? dirty_0_61 : _GEN_8149; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9564 = unuse_way == 2'h2 ? dirty_0_62 : _GEN_8150; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9565 = unuse_way == 2'h2 ? dirty_0_63 : _GEN_8151; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9566 = unuse_way == 2'h2 ? dirty_0_64 : _GEN_8152; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9567 = unuse_way == 2'h2 ? dirty_0_65 : _GEN_8153; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9568 = unuse_way == 2'h2 ? dirty_0_66 : _GEN_8154; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9569 = unuse_way == 2'h2 ? dirty_0_67 : _GEN_8155; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9570 = unuse_way == 2'h2 ? dirty_0_68 : _GEN_8156; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9571 = unuse_way == 2'h2 ? dirty_0_69 : _GEN_8157; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9572 = unuse_way == 2'h2 ? dirty_0_70 : _GEN_8158; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9573 = unuse_way == 2'h2 ? dirty_0_71 : _GEN_8159; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9574 = unuse_way == 2'h2 ? dirty_0_72 : _GEN_8160; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9575 = unuse_way == 2'h2 ? dirty_0_73 : _GEN_8161; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9576 = unuse_way == 2'h2 ? dirty_0_74 : _GEN_8162; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9577 = unuse_way == 2'h2 ? dirty_0_75 : _GEN_8163; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9578 = unuse_way == 2'h2 ? dirty_0_76 : _GEN_8164; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9579 = unuse_way == 2'h2 ? dirty_0_77 : _GEN_8165; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9580 = unuse_way == 2'h2 ? dirty_0_78 : _GEN_8166; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9581 = unuse_way == 2'h2 ? dirty_0_79 : _GEN_8167; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9582 = unuse_way == 2'h2 ? dirty_0_80 : _GEN_8168; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9583 = unuse_way == 2'h2 ? dirty_0_81 : _GEN_8169; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9584 = unuse_way == 2'h2 ? dirty_0_82 : _GEN_8170; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9585 = unuse_way == 2'h2 ? dirty_0_83 : _GEN_8171; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9586 = unuse_way == 2'h2 ? dirty_0_84 : _GEN_8172; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9587 = unuse_way == 2'h2 ? dirty_0_85 : _GEN_8173; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9588 = unuse_way == 2'h2 ? dirty_0_86 : _GEN_8174; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9589 = unuse_way == 2'h2 ? dirty_0_87 : _GEN_8175; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9590 = unuse_way == 2'h2 ? dirty_0_88 : _GEN_8176; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9591 = unuse_way == 2'h2 ? dirty_0_89 : _GEN_8177; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9592 = unuse_way == 2'h2 ? dirty_0_90 : _GEN_8178; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9593 = unuse_way == 2'h2 ? dirty_0_91 : _GEN_8179; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9594 = unuse_way == 2'h2 ? dirty_0_92 : _GEN_8180; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9595 = unuse_way == 2'h2 ? dirty_0_93 : _GEN_8181; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9596 = unuse_way == 2'h2 ? dirty_0_94 : _GEN_8182; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9597 = unuse_way == 2'h2 ? dirty_0_95 : _GEN_8183; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9598 = unuse_way == 2'h2 ? dirty_0_96 : _GEN_8184; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9599 = unuse_way == 2'h2 ? dirty_0_97 : _GEN_8185; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9600 = unuse_way == 2'h2 ? dirty_0_98 : _GEN_8186; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9601 = unuse_way == 2'h2 ? dirty_0_99 : _GEN_8187; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9602 = unuse_way == 2'h2 ? dirty_0_100 : _GEN_8188; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9603 = unuse_way == 2'h2 ? dirty_0_101 : _GEN_8189; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9604 = unuse_way == 2'h2 ? dirty_0_102 : _GEN_8190; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9605 = unuse_way == 2'h2 ? dirty_0_103 : _GEN_8191; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9606 = unuse_way == 2'h2 ? dirty_0_104 : _GEN_8192; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9607 = unuse_way == 2'h2 ? dirty_0_105 : _GEN_8193; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9608 = unuse_way == 2'h2 ? dirty_0_106 : _GEN_8194; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9609 = unuse_way == 2'h2 ? dirty_0_107 : _GEN_8195; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9610 = unuse_way == 2'h2 ? dirty_0_108 : _GEN_8196; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9611 = unuse_way == 2'h2 ? dirty_0_109 : _GEN_8197; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9612 = unuse_way == 2'h2 ? dirty_0_110 : _GEN_8198; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9613 = unuse_way == 2'h2 ? dirty_0_111 : _GEN_8199; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9614 = unuse_way == 2'h2 ? dirty_0_112 : _GEN_8200; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9615 = unuse_way == 2'h2 ? dirty_0_113 : _GEN_8201; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9616 = unuse_way == 2'h2 ? dirty_0_114 : _GEN_8202; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9617 = unuse_way == 2'h2 ? dirty_0_115 : _GEN_8203; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9618 = unuse_way == 2'h2 ? dirty_0_116 : _GEN_8204; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9619 = unuse_way == 2'h2 ? dirty_0_117 : _GEN_8205; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9620 = unuse_way == 2'h2 ? dirty_0_118 : _GEN_8206; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9621 = unuse_way == 2'h2 ? dirty_0_119 : _GEN_8207; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9622 = unuse_way == 2'h2 ? dirty_0_120 : _GEN_8208; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9623 = unuse_way == 2'h2 ? dirty_0_121 : _GEN_8209; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9624 = unuse_way == 2'h2 ? dirty_0_122 : _GEN_8210; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9625 = unuse_way == 2'h2 ? dirty_0_123 : _GEN_8211; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9626 = unuse_way == 2'h2 ? dirty_0_124 : _GEN_8212; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9627 = unuse_way == 2'h2 ? dirty_0_125 : _GEN_8213; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9628 = unuse_way == 2'h2 ? dirty_0_126 : _GEN_8214; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9629 = unuse_way == 2'h2 ? dirty_0_127 : _GEN_8215; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_9630 = unuse_way == 2'h2 ? valid_0_0 : _GEN_8216; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9631 = unuse_way == 2'h2 ? valid_0_1 : _GEN_8217; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9632 = unuse_way == 2'h2 ? valid_0_2 : _GEN_8218; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9633 = unuse_way == 2'h2 ? valid_0_3 : _GEN_8219; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9634 = unuse_way == 2'h2 ? valid_0_4 : _GEN_8220; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9635 = unuse_way == 2'h2 ? valid_0_5 : _GEN_8221; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9636 = unuse_way == 2'h2 ? valid_0_6 : _GEN_8222; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9637 = unuse_way == 2'h2 ? valid_0_7 : _GEN_8223; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9638 = unuse_way == 2'h2 ? valid_0_8 : _GEN_8224; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9639 = unuse_way == 2'h2 ? valid_0_9 : _GEN_8225; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9640 = unuse_way == 2'h2 ? valid_0_10 : _GEN_8226; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9641 = unuse_way == 2'h2 ? valid_0_11 : _GEN_8227; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9642 = unuse_way == 2'h2 ? valid_0_12 : _GEN_8228; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9643 = unuse_way == 2'h2 ? valid_0_13 : _GEN_8229; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9644 = unuse_way == 2'h2 ? valid_0_14 : _GEN_8230; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9645 = unuse_way == 2'h2 ? valid_0_15 : _GEN_8231; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9646 = unuse_way == 2'h2 ? valid_0_16 : _GEN_8232; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9647 = unuse_way == 2'h2 ? valid_0_17 : _GEN_8233; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9648 = unuse_way == 2'h2 ? valid_0_18 : _GEN_8234; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9649 = unuse_way == 2'h2 ? valid_0_19 : _GEN_8235; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9650 = unuse_way == 2'h2 ? valid_0_20 : _GEN_8236; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9651 = unuse_way == 2'h2 ? valid_0_21 : _GEN_8237; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9652 = unuse_way == 2'h2 ? valid_0_22 : _GEN_8238; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9653 = unuse_way == 2'h2 ? valid_0_23 : _GEN_8239; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9654 = unuse_way == 2'h2 ? valid_0_24 : _GEN_8240; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9655 = unuse_way == 2'h2 ? valid_0_25 : _GEN_8241; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9656 = unuse_way == 2'h2 ? valid_0_26 : _GEN_8242; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9657 = unuse_way == 2'h2 ? valid_0_27 : _GEN_8243; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9658 = unuse_way == 2'h2 ? valid_0_28 : _GEN_8244; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9659 = unuse_way == 2'h2 ? valid_0_29 : _GEN_8245; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9660 = unuse_way == 2'h2 ? valid_0_30 : _GEN_8246; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9661 = unuse_way == 2'h2 ? valid_0_31 : _GEN_8247; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9662 = unuse_way == 2'h2 ? valid_0_32 : _GEN_8248; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9663 = unuse_way == 2'h2 ? valid_0_33 : _GEN_8249; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9664 = unuse_way == 2'h2 ? valid_0_34 : _GEN_8250; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9665 = unuse_way == 2'h2 ? valid_0_35 : _GEN_8251; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9666 = unuse_way == 2'h2 ? valid_0_36 : _GEN_8252; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9667 = unuse_way == 2'h2 ? valid_0_37 : _GEN_8253; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9668 = unuse_way == 2'h2 ? valid_0_38 : _GEN_8254; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9669 = unuse_way == 2'h2 ? valid_0_39 : _GEN_8255; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9670 = unuse_way == 2'h2 ? valid_0_40 : _GEN_8256; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9671 = unuse_way == 2'h2 ? valid_0_41 : _GEN_8257; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9672 = unuse_way == 2'h2 ? valid_0_42 : _GEN_8258; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9673 = unuse_way == 2'h2 ? valid_0_43 : _GEN_8259; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9674 = unuse_way == 2'h2 ? valid_0_44 : _GEN_8260; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9675 = unuse_way == 2'h2 ? valid_0_45 : _GEN_8261; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9676 = unuse_way == 2'h2 ? valid_0_46 : _GEN_8262; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9677 = unuse_way == 2'h2 ? valid_0_47 : _GEN_8263; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9678 = unuse_way == 2'h2 ? valid_0_48 : _GEN_8264; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9679 = unuse_way == 2'h2 ? valid_0_49 : _GEN_8265; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9680 = unuse_way == 2'h2 ? valid_0_50 : _GEN_8266; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9681 = unuse_way == 2'h2 ? valid_0_51 : _GEN_8267; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9682 = unuse_way == 2'h2 ? valid_0_52 : _GEN_8268; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9683 = unuse_way == 2'h2 ? valid_0_53 : _GEN_8269; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9684 = unuse_way == 2'h2 ? valid_0_54 : _GEN_8270; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9685 = unuse_way == 2'h2 ? valid_0_55 : _GEN_8271; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9686 = unuse_way == 2'h2 ? valid_0_56 : _GEN_8272; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9687 = unuse_way == 2'h2 ? valid_0_57 : _GEN_8273; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9688 = unuse_way == 2'h2 ? valid_0_58 : _GEN_8274; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9689 = unuse_way == 2'h2 ? valid_0_59 : _GEN_8275; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9690 = unuse_way == 2'h2 ? valid_0_60 : _GEN_8276; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9691 = unuse_way == 2'h2 ? valid_0_61 : _GEN_8277; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9692 = unuse_way == 2'h2 ? valid_0_62 : _GEN_8278; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9693 = unuse_way == 2'h2 ? valid_0_63 : _GEN_8279; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9694 = unuse_way == 2'h2 ? valid_0_64 : _GEN_8280; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9695 = unuse_way == 2'h2 ? valid_0_65 : _GEN_8281; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9696 = unuse_way == 2'h2 ? valid_0_66 : _GEN_8282; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9697 = unuse_way == 2'h2 ? valid_0_67 : _GEN_8283; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9698 = unuse_way == 2'h2 ? valid_0_68 : _GEN_8284; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9699 = unuse_way == 2'h2 ? valid_0_69 : _GEN_8285; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9700 = unuse_way == 2'h2 ? valid_0_70 : _GEN_8286; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9701 = unuse_way == 2'h2 ? valid_0_71 : _GEN_8287; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9702 = unuse_way == 2'h2 ? valid_0_72 : _GEN_8288; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9703 = unuse_way == 2'h2 ? valid_0_73 : _GEN_8289; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9704 = unuse_way == 2'h2 ? valid_0_74 : _GEN_8290; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9705 = unuse_way == 2'h2 ? valid_0_75 : _GEN_8291; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9706 = unuse_way == 2'h2 ? valid_0_76 : _GEN_8292; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9707 = unuse_way == 2'h2 ? valid_0_77 : _GEN_8293; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9708 = unuse_way == 2'h2 ? valid_0_78 : _GEN_8294; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9709 = unuse_way == 2'h2 ? valid_0_79 : _GEN_8295; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9710 = unuse_way == 2'h2 ? valid_0_80 : _GEN_8296; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9711 = unuse_way == 2'h2 ? valid_0_81 : _GEN_8297; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9712 = unuse_way == 2'h2 ? valid_0_82 : _GEN_8298; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9713 = unuse_way == 2'h2 ? valid_0_83 : _GEN_8299; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9714 = unuse_way == 2'h2 ? valid_0_84 : _GEN_8300; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9715 = unuse_way == 2'h2 ? valid_0_85 : _GEN_8301; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9716 = unuse_way == 2'h2 ? valid_0_86 : _GEN_8302; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9717 = unuse_way == 2'h2 ? valid_0_87 : _GEN_8303; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9718 = unuse_way == 2'h2 ? valid_0_88 : _GEN_8304; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9719 = unuse_way == 2'h2 ? valid_0_89 : _GEN_8305; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9720 = unuse_way == 2'h2 ? valid_0_90 : _GEN_8306; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9721 = unuse_way == 2'h2 ? valid_0_91 : _GEN_8307; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9722 = unuse_way == 2'h2 ? valid_0_92 : _GEN_8308; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9723 = unuse_way == 2'h2 ? valid_0_93 : _GEN_8309; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9724 = unuse_way == 2'h2 ? valid_0_94 : _GEN_8310; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9725 = unuse_way == 2'h2 ? valid_0_95 : _GEN_8311; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9726 = unuse_way == 2'h2 ? valid_0_96 : _GEN_8312; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9727 = unuse_way == 2'h2 ? valid_0_97 : _GEN_8313; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9728 = unuse_way == 2'h2 ? valid_0_98 : _GEN_8314; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9729 = unuse_way == 2'h2 ? valid_0_99 : _GEN_8315; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9730 = unuse_way == 2'h2 ? valid_0_100 : _GEN_8316; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9731 = unuse_way == 2'h2 ? valid_0_101 : _GEN_8317; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9732 = unuse_way == 2'h2 ? valid_0_102 : _GEN_8318; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9733 = unuse_way == 2'h2 ? valid_0_103 : _GEN_8319; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9734 = unuse_way == 2'h2 ? valid_0_104 : _GEN_8320; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9735 = unuse_way == 2'h2 ? valid_0_105 : _GEN_8321; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9736 = unuse_way == 2'h2 ? valid_0_106 : _GEN_8322; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9737 = unuse_way == 2'h2 ? valid_0_107 : _GEN_8323; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9738 = unuse_way == 2'h2 ? valid_0_108 : _GEN_8324; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9739 = unuse_way == 2'h2 ? valid_0_109 : _GEN_8325; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9740 = unuse_way == 2'h2 ? valid_0_110 : _GEN_8326; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9741 = unuse_way == 2'h2 ? valid_0_111 : _GEN_8327; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9742 = unuse_way == 2'h2 ? valid_0_112 : _GEN_8328; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9743 = unuse_way == 2'h2 ? valid_0_113 : _GEN_8329; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9744 = unuse_way == 2'h2 ? valid_0_114 : _GEN_8330; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9745 = unuse_way == 2'h2 ? valid_0_115 : _GEN_8331; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9746 = unuse_way == 2'h2 ? valid_0_116 : _GEN_8332; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9747 = unuse_way == 2'h2 ? valid_0_117 : _GEN_8333; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9748 = unuse_way == 2'h2 ? valid_0_118 : _GEN_8334; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9749 = unuse_way == 2'h2 ? valid_0_119 : _GEN_8335; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9750 = unuse_way == 2'h2 ? valid_0_120 : _GEN_8336; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9751 = unuse_way == 2'h2 ? valid_0_121 : _GEN_8337; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9752 = unuse_way == 2'h2 ? valid_0_122 : _GEN_8338; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9753 = unuse_way == 2'h2 ? valid_0_123 : _GEN_8339; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9754 = unuse_way == 2'h2 ? valid_0_124 : _GEN_8340; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9755 = unuse_way == 2'h2 ? valid_0_125 : _GEN_8341; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9756 = unuse_way == 2'h2 ? valid_0_126 : _GEN_8342; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9757 = unuse_way == 2'h2 ? valid_0_127 : _GEN_8343; // @[d_cache.scala 156:40 30:26]
  wire  _GEN_9758 = unuse_way == 2'h2 ? dirty_1_0 : _GEN_8602; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9759 = unuse_way == 2'h2 ? dirty_1_1 : _GEN_8603; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9760 = unuse_way == 2'h2 ? dirty_1_2 : _GEN_8604; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9761 = unuse_way == 2'h2 ? dirty_1_3 : _GEN_8605; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9762 = unuse_way == 2'h2 ? dirty_1_4 : _GEN_8606; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9763 = unuse_way == 2'h2 ? dirty_1_5 : _GEN_8607; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9764 = unuse_way == 2'h2 ? dirty_1_6 : _GEN_8608; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9765 = unuse_way == 2'h2 ? dirty_1_7 : _GEN_8609; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9766 = unuse_way == 2'h2 ? dirty_1_8 : _GEN_8610; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9767 = unuse_way == 2'h2 ? dirty_1_9 : _GEN_8611; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9768 = unuse_way == 2'h2 ? dirty_1_10 : _GEN_8612; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9769 = unuse_way == 2'h2 ? dirty_1_11 : _GEN_8613; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9770 = unuse_way == 2'h2 ? dirty_1_12 : _GEN_8614; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9771 = unuse_way == 2'h2 ? dirty_1_13 : _GEN_8615; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9772 = unuse_way == 2'h2 ? dirty_1_14 : _GEN_8616; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9773 = unuse_way == 2'h2 ? dirty_1_15 : _GEN_8617; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9774 = unuse_way == 2'h2 ? dirty_1_16 : _GEN_8618; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9775 = unuse_way == 2'h2 ? dirty_1_17 : _GEN_8619; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9776 = unuse_way == 2'h2 ? dirty_1_18 : _GEN_8620; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9777 = unuse_way == 2'h2 ? dirty_1_19 : _GEN_8621; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9778 = unuse_way == 2'h2 ? dirty_1_20 : _GEN_8622; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9779 = unuse_way == 2'h2 ? dirty_1_21 : _GEN_8623; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9780 = unuse_way == 2'h2 ? dirty_1_22 : _GEN_8624; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9781 = unuse_way == 2'h2 ? dirty_1_23 : _GEN_8625; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9782 = unuse_way == 2'h2 ? dirty_1_24 : _GEN_8626; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9783 = unuse_way == 2'h2 ? dirty_1_25 : _GEN_8627; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9784 = unuse_way == 2'h2 ? dirty_1_26 : _GEN_8628; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9785 = unuse_way == 2'h2 ? dirty_1_27 : _GEN_8629; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9786 = unuse_way == 2'h2 ? dirty_1_28 : _GEN_8630; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9787 = unuse_way == 2'h2 ? dirty_1_29 : _GEN_8631; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9788 = unuse_way == 2'h2 ? dirty_1_30 : _GEN_8632; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9789 = unuse_way == 2'h2 ? dirty_1_31 : _GEN_8633; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9790 = unuse_way == 2'h2 ? dirty_1_32 : _GEN_8634; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9791 = unuse_way == 2'h2 ? dirty_1_33 : _GEN_8635; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9792 = unuse_way == 2'h2 ? dirty_1_34 : _GEN_8636; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9793 = unuse_way == 2'h2 ? dirty_1_35 : _GEN_8637; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9794 = unuse_way == 2'h2 ? dirty_1_36 : _GEN_8638; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9795 = unuse_way == 2'h2 ? dirty_1_37 : _GEN_8639; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9796 = unuse_way == 2'h2 ? dirty_1_38 : _GEN_8640; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9797 = unuse_way == 2'h2 ? dirty_1_39 : _GEN_8641; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9798 = unuse_way == 2'h2 ? dirty_1_40 : _GEN_8642; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9799 = unuse_way == 2'h2 ? dirty_1_41 : _GEN_8643; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9800 = unuse_way == 2'h2 ? dirty_1_42 : _GEN_8644; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9801 = unuse_way == 2'h2 ? dirty_1_43 : _GEN_8645; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9802 = unuse_way == 2'h2 ? dirty_1_44 : _GEN_8646; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9803 = unuse_way == 2'h2 ? dirty_1_45 : _GEN_8647; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9804 = unuse_way == 2'h2 ? dirty_1_46 : _GEN_8648; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9805 = unuse_way == 2'h2 ? dirty_1_47 : _GEN_8649; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9806 = unuse_way == 2'h2 ? dirty_1_48 : _GEN_8650; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9807 = unuse_way == 2'h2 ? dirty_1_49 : _GEN_8651; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9808 = unuse_way == 2'h2 ? dirty_1_50 : _GEN_8652; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9809 = unuse_way == 2'h2 ? dirty_1_51 : _GEN_8653; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9810 = unuse_way == 2'h2 ? dirty_1_52 : _GEN_8654; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9811 = unuse_way == 2'h2 ? dirty_1_53 : _GEN_8655; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9812 = unuse_way == 2'h2 ? dirty_1_54 : _GEN_8656; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9813 = unuse_way == 2'h2 ? dirty_1_55 : _GEN_8657; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9814 = unuse_way == 2'h2 ? dirty_1_56 : _GEN_8658; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9815 = unuse_way == 2'h2 ? dirty_1_57 : _GEN_8659; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9816 = unuse_way == 2'h2 ? dirty_1_58 : _GEN_8660; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9817 = unuse_way == 2'h2 ? dirty_1_59 : _GEN_8661; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9818 = unuse_way == 2'h2 ? dirty_1_60 : _GEN_8662; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9819 = unuse_way == 2'h2 ? dirty_1_61 : _GEN_8663; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9820 = unuse_way == 2'h2 ? dirty_1_62 : _GEN_8664; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9821 = unuse_way == 2'h2 ? dirty_1_63 : _GEN_8665; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9822 = unuse_way == 2'h2 ? dirty_1_64 : _GEN_8666; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9823 = unuse_way == 2'h2 ? dirty_1_65 : _GEN_8667; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9824 = unuse_way == 2'h2 ? dirty_1_66 : _GEN_8668; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9825 = unuse_way == 2'h2 ? dirty_1_67 : _GEN_8669; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9826 = unuse_way == 2'h2 ? dirty_1_68 : _GEN_8670; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9827 = unuse_way == 2'h2 ? dirty_1_69 : _GEN_8671; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9828 = unuse_way == 2'h2 ? dirty_1_70 : _GEN_8672; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9829 = unuse_way == 2'h2 ? dirty_1_71 : _GEN_8673; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9830 = unuse_way == 2'h2 ? dirty_1_72 : _GEN_8674; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9831 = unuse_way == 2'h2 ? dirty_1_73 : _GEN_8675; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9832 = unuse_way == 2'h2 ? dirty_1_74 : _GEN_8676; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9833 = unuse_way == 2'h2 ? dirty_1_75 : _GEN_8677; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9834 = unuse_way == 2'h2 ? dirty_1_76 : _GEN_8678; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9835 = unuse_way == 2'h2 ? dirty_1_77 : _GEN_8679; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9836 = unuse_way == 2'h2 ? dirty_1_78 : _GEN_8680; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9837 = unuse_way == 2'h2 ? dirty_1_79 : _GEN_8681; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9838 = unuse_way == 2'h2 ? dirty_1_80 : _GEN_8682; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9839 = unuse_way == 2'h2 ? dirty_1_81 : _GEN_8683; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9840 = unuse_way == 2'h2 ? dirty_1_82 : _GEN_8684; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9841 = unuse_way == 2'h2 ? dirty_1_83 : _GEN_8685; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9842 = unuse_way == 2'h2 ? dirty_1_84 : _GEN_8686; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9843 = unuse_way == 2'h2 ? dirty_1_85 : _GEN_8687; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9844 = unuse_way == 2'h2 ? dirty_1_86 : _GEN_8688; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9845 = unuse_way == 2'h2 ? dirty_1_87 : _GEN_8689; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9846 = unuse_way == 2'h2 ? dirty_1_88 : _GEN_8690; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9847 = unuse_way == 2'h2 ? dirty_1_89 : _GEN_8691; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9848 = unuse_way == 2'h2 ? dirty_1_90 : _GEN_8692; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9849 = unuse_way == 2'h2 ? dirty_1_91 : _GEN_8693; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9850 = unuse_way == 2'h2 ? dirty_1_92 : _GEN_8694; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9851 = unuse_way == 2'h2 ? dirty_1_93 : _GEN_8695; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9852 = unuse_way == 2'h2 ? dirty_1_94 : _GEN_8696; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9853 = unuse_way == 2'h2 ? dirty_1_95 : _GEN_8697; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9854 = unuse_way == 2'h2 ? dirty_1_96 : _GEN_8698; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9855 = unuse_way == 2'h2 ? dirty_1_97 : _GEN_8699; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9856 = unuse_way == 2'h2 ? dirty_1_98 : _GEN_8700; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9857 = unuse_way == 2'h2 ? dirty_1_99 : _GEN_8701; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9858 = unuse_way == 2'h2 ? dirty_1_100 : _GEN_8702; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9859 = unuse_way == 2'h2 ? dirty_1_101 : _GEN_8703; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9860 = unuse_way == 2'h2 ? dirty_1_102 : _GEN_8704; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9861 = unuse_way == 2'h2 ? dirty_1_103 : _GEN_8705; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9862 = unuse_way == 2'h2 ? dirty_1_104 : _GEN_8706; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9863 = unuse_way == 2'h2 ? dirty_1_105 : _GEN_8707; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9864 = unuse_way == 2'h2 ? dirty_1_106 : _GEN_8708; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9865 = unuse_way == 2'h2 ? dirty_1_107 : _GEN_8709; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9866 = unuse_way == 2'h2 ? dirty_1_108 : _GEN_8710; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9867 = unuse_way == 2'h2 ? dirty_1_109 : _GEN_8711; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9868 = unuse_way == 2'h2 ? dirty_1_110 : _GEN_8712; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9869 = unuse_way == 2'h2 ? dirty_1_111 : _GEN_8713; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9870 = unuse_way == 2'h2 ? dirty_1_112 : _GEN_8714; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9871 = unuse_way == 2'h2 ? dirty_1_113 : _GEN_8715; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9872 = unuse_way == 2'h2 ? dirty_1_114 : _GEN_8716; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9873 = unuse_way == 2'h2 ? dirty_1_115 : _GEN_8717; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9874 = unuse_way == 2'h2 ? dirty_1_116 : _GEN_8718; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9875 = unuse_way == 2'h2 ? dirty_1_117 : _GEN_8719; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9876 = unuse_way == 2'h2 ? dirty_1_118 : _GEN_8720; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9877 = unuse_way == 2'h2 ? dirty_1_119 : _GEN_8721; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9878 = unuse_way == 2'h2 ? dirty_1_120 : _GEN_8722; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9879 = unuse_way == 2'h2 ? dirty_1_121 : _GEN_8723; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9880 = unuse_way == 2'h2 ? dirty_1_122 : _GEN_8724; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9881 = unuse_way == 2'h2 ? dirty_1_123 : _GEN_8725; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9882 = unuse_way == 2'h2 ? dirty_1_124 : _GEN_8726; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9883 = unuse_way == 2'h2 ? dirty_1_125 : _GEN_8727; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9884 = unuse_way == 2'h2 ? dirty_1_126 : _GEN_8728; // @[d_cache.scala 156:40 33:26]
  wire  _GEN_9885 = unuse_way == 2'h2 ? dirty_1_127 : _GEN_8729; // @[d_cache.scala 156:40 33:26]
  wire [2:0] _GEN_9886 = unuse_way == 2'h1 ? 3'h7 : _GEN_8858; // @[d_cache.scala 150:34 151:23]
  wire [63:0] _GEN_9887 = unuse_way == 2'h1 ? _GEN_4238 : _GEN_9246; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9888 = unuse_way == 2'h1 ? _GEN_4239 : _GEN_9247; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9889 = unuse_way == 2'h1 ? _GEN_4240 : _GEN_9248; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9890 = unuse_way == 2'h1 ? _GEN_4241 : _GEN_9249; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9891 = unuse_way == 2'h1 ? _GEN_4242 : _GEN_9250; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9892 = unuse_way == 2'h1 ? _GEN_4243 : _GEN_9251; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9893 = unuse_way == 2'h1 ? _GEN_4244 : _GEN_9252; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9894 = unuse_way == 2'h1 ? _GEN_4245 : _GEN_9253; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9895 = unuse_way == 2'h1 ? _GEN_4246 : _GEN_9254; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9896 = unuse_way == 2'h1 ? _GEN_4247 : _GEN_9255; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9897 = unuse_way == 2'h1 ? _GEN_4248 : _GEN_9256; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9898 = unuse_way == 2'h1 ? _GEN_4249 : _GEN_9257; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9899 = unuse_way == 2'h1 ? _GEN_4250 : _GEN_9258; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9900 = unuse_way == 2'h1 ? _GEN_4251 : _GEN_9259; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9901 = unuse_way == 2'h1 ? _GEN_4252 : _GEN_9260; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9902 = unuse_way == 2'h1 ? _GEN_4253 : _GEN_9261; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9903 = unuse_way == 2'h1 ? _GEN_4254 : _GEN_9262; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9904 = unuse_way == 2'h1 ? _GEN_4255 : _GEN_9263; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9905 = unuse_way == 2'h1 ? _GEN_4256 : _GEN_9264; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9906 = unuse_way == 2'h1 ? _GEN_4257 : _GEN_9265; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9907 = unuse_way == 2'h1 ? _GEN_4258 : _GEN_9266; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9908 = unuse_way == 2'h1 ? _GEN_4259 : _GEN_9267; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9909 = unuse_way == 2'h1 ? _GEN_4260 : _GEN_9268; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9910 = unuse_way == 2'h1 ? _GEN_4261 : _GEN_9269; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9911 = unuse_way == 2'h1 ? _GEN_4262 : _GEN_9270; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9912 = unuse_way == 2'h1 ? _GEN_4263 : _GEN_9271; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9913 = unuse_way == 2'h1 ? _GEN_4264 : _GEN_9272; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9914 = unuse_way == 2'h1 ? _GEN_4265 : _GEN_9273; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9915 = unuse_way == 2'h1 ? _GEN_4266 : _GEN_9274; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9916 = unuse_way == 2'h1 ? _GEN_4267 : _GEN_9275; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9917 = unuse_way == 2'h1 ? _GEN_4268 : _GEN_9276; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9918 = unuse_way == 2'h1 ? _GEN_4269 : _GEN_9277; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9919 = unuse_way == 2'h1 ? _GEN_4270 : _GEN_9278; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9920 = unuse_way == 2'h1 ? _GEN_4271 : _GEN_9279; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9921 = unuse_way == 2'h1 ? _GEN_4272 : _GEN_9280; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9922 = unuse_way == 2'h1 ? _GEN_4273 : _GEN_9281; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9923 = unuse_way == 2'h1 ? _GEN_4274 : _GEN_9282; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9924 = unuse_way == 2'h1 ? _GEN_4275 : _GEN_9283; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9925 = unuse_way == 2'h1 ? _GEN_4276 : _GEN_9284; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9926 = unuse_way == 2'h1 ? _GEN_4277 : _GEN_9285; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9927 = unuse_way == 2'h1 ? _GEN_4278 : _GEN_9286; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9928 = unuse_way == 2'h1 ? _GEN_4279 : _GEN_9287; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9929 = unuse_way == 2'h1 ? _GEN_4280 : _GEN_9288; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9930 = unuse_way == 2'h1 ? _GEN_4281 : _GEN_9289; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9931 = unuse_way == 2'h1 ? _GEN_4282 : _GEN_9290; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9932 = unuse_way == 2'h1 ? _GEN_4283 : _GEN_9291; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9933 = unuse_way == 2'h1 ? _GEN_4284 : _GEN_9292; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9934 = unuse_way == 2'h1 ? _GEN_4285 : _GEN_9293; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9935 = unuse_way == 2'h1 ? _GEN_4286 : _GEN_9294; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9936 = unuse_way == 2'h1 ? _GEN_4287 : _GEN_9295; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9937 = unuse_way == 2'h1 ? _GEN_4288 : _GEN_9296; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9938 = unuse_way == 2'h1 ? _GEN_4289 : _GEN_9297; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9939 = unuse_way == 2'h1 ? _GEN_4290 : _GEN_9298; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9940 = unuse_way == 2'h1 ? _GEN_4291 : _GEN_9299; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9941 = unuse_way == 2'h1 ? _GEN_4292 : _GEN_9300; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9942 = unuse_way == 2'h1 ? _GEN_4293 : _GEN_9301; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9943 = unuse_way == 2'h1 ? _GEN_4294 : _GEN_9302; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9944 = unuse_way == 2'h1 ? _GEN_4295 : _GEN_9303; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9945 = unuse_way == 2'h1 ? _GEN_4296 : _GEN_9304; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9946 = unuse_way == 2'h1 ? _GEN_4297 : _GEN_9305; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9947 = unuse_way == 2'h1 ? _GEN_4298 : _GEN_9306; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9948 = unuse_way == 2'h1 ? _GEN_4299 : _GEN_9307; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9949 = unuse_way == 2'h1 ? _GEN_4300 : _GEN_9308; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9950 = unuse_way == 2'h1 ? _GEN_4301 : _GEN_9309; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9951 = unuse_way == 2'h1 ? _GEN_4302 : _GEN_9310; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9952 = unuse_way == 2'h1 ? _GEN_4303 : _GEN_9311; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9953 = unuse_way == 2'h1 ? _GEN_4304 : _GEN_9312; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9954 = unuse_way == 2'h1 ? _GEN_4305 : _GEN_9313; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9955 = unuse_way == 2'h1 ? _GEN_4306 : _GEN_9314; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9956 = unuse_way == 2'h1 ? _GEN_4307 : _GEN_9315; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9957 = unuse_way == 2'h1 ? _GEN_4308 : _GEN_9316; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9958 = unuse_way == 2'h1 ? _GEN_4309 : _GEN_9317; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9959 = unuse_way == 2'h1 ? _GEN_4310 : _GEN_9318; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9960 = unuse_way == 2'h1 ? _GEN_4311 : _GEN_9319; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9961 = unuse_way == 2'h1 ? _GEN_4312 : _GEN_9320; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9962 = unuse_way == 2'h1 ? _GEN_4313 : _GEN_9321; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9963 = unuse_way == 2'h1 ? _GEN_4314 : _GEN_9322; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9964 = unuse_way == 2'h1 ? _GEN_4315 : _GEN_9323; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9965 = unuse_way == 2'h1 ? _GEN_4316 : _GEN_9324; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9966 = unuse_way == 2'h1 ? _GEN_4317 : _GEN_9325; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9967 = unuse_way == 2'h1 ? _GEN_4318 : _GEN_9326; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9968 = unuse_way == 2'h1 ? _GEN_4319 : _GEN_9327; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9969 = unuse_way == 2'h1 ? _GEN_4320 : _GEN_9328; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9970 = unuse_way == 2'h1 ? _GEN_4321 : _GEN_9329; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9971 = unuse_way == 2'h1 ? _GEN_4322 : _GEN_9330; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9972 = unuse_way == 2'h1 ? _GEN_4323 : _GEN_9331; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9973 = unuse_way == 2'h1 ? _GEN_4324 : _GEN_9332; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9974 = unuse_way == 2'h1 ? _GEN_4325 : _GEN_9333; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9975 = unuse_way == 2'h1 ? _GEN_4326 : _GEN_9334; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9976 = unuse_way == 2'h1 ? _GEN_4327 : _GEN_9335; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9977 = unuse_way == 2'h1 ? _GEN_4328 : _GEN_9336; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9978 = unuse_way == 2'h1 ? _GEN_4329 : _GEN_9337; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9979 = unuse_way == 2'h1 ? _GEN_4330 : _GEN_9338; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9980 = unuse_way == 2'h1 ? _GEN_4331 : _GEN_9339; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9981 = unuse_way == 2'h1 ? _GEN_4332 : _GEN_9340; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9982 = unuse_way == 2'h1 ? _GEN_4333 : _GEN_9341; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9983 = unuse_way == 2'h1 ? _GEN_4334 : _GEN_9342; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9984 = unuse_way == 2'h1 ? _GEN_4335 : _GEN_9343; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9985 = unuse_way == 2'h1 ? _GEN_4336 : _GEN_9344; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9986 = unuse_way == 2'h1 ? _GEN_4337 : _GEN_9345; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9987 = unuse_way == 2'h1 ? _GEN_4338 : _GEN_9346; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9988 = unuse_way == 2'h1 ? _GEN_4339 : _GEN_9347; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9989 = unuse_way == 2'h1 ? _GEN_4340 : _GEN_9348; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9990 = unuse_way == 2'h1 ? _GEN_4341 : _GEN_9349; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9991 = unuse_way == 2'h1 ? _GEN_4342 : _GEN_9350; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9992 = unuse_way == 2'h1 ? _GEN_4343 : _GEN_9351; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9993 = unuse_way == 2'h1 ? _GEN_4344 : _GEN_9352; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9994 = unuse_way == 2'h1 ? _GEN_4345 : _GEN_9353; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9995 = unuse_way == 2'h1 ? _GEN_4346 : _GEN_9354; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9996 = unuse_way == 2'h1 ? _GEN_4347 : _GEN_9355; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9997 = unuse_way == 2'h1 ? _GEN_4348 : _GEN_9356; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9998 = unuse_way == 2'h1 ? _GEN_4349 : _GEN_9357; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_9999 = unuse_way == 2'h1 ? _GEN_4350 : _GEN_9358; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10000 = unuse_way == 2'h1 ? _GEN_4351 : _GEN_9359; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10001 = unuse_way == 2'h1 ? _GEN_4352 : _GEN_9360; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10002 = unuse_way == 2'h1 ? _GEN_4353 : _GEN_9361; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10003 = unuse_way == 2'h1 ? _GEN_4354 : _GEN_9362; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10004 = unuse_way == 2'h1 ? _GEN_4355 : _GEN_9363; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10005 = unuse_way == 2'h1 ? _GEN_4356 : _GEN_9364; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10006 = unuse_way == 2'h1 ? _GEN_4357 : _GEN_9365; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10007 = unuse_way == 2'h1 ? _GEN_4358 : _GEN_9366; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10008 = unuse_way == 2'h1 ? _GEN_4359 : _GEN_9367; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10009 = unuse_way == 2'h1 ? _GEN_4360 : _GEN_9368; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10010 = unuse_way == 2'h1 ? _GEN_4361 : _GEN_9369; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10011 = unuse_way == 2'h1 ? _GEN_4362 : _GEN_9370; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10012 = unuse_way == 2'h1 ? _GEN_4363 : _GEN_9371; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10013 = unuse_way == 2'h1 ? _GEN_4364 : _GEN_9372; // @[d_cache.scala 150:34]
  wire [63:0] _GEN_10014 = unuse_way == 2'h1 ? _GEN_4365 : _GEN_9373; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10015 = unuse_way == 2'h1 ? _GEN_4366 : _GEN_9374; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10016 = unuse_way == 2'h1 ? _GEN_4367 : _GEN_9375; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10017 = unuse_way == 2'h1 ? _GEN_4368 : _GEN_9376; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10018 = unuse_way == 2'h1 ? _GEN_4369 : _GEN_9377; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10019 = unuse_way == 2'h1 ? _GEN_4370 : _GEN_9378; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10020 = unuse_way == 2'h1 ? _GEN_4371 : _GEN_9379; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10021 = unuse_way == 2'h1 ? _GEN_4372 : _GEN_9380; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10022 = unuse_way == 2'h1 ? _GEN_4373 : _GEN_9381; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10023 = unuse_way == 2'h1 ? _GEN_4374 : _GEN_9382; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10024 = unuse_way == 2'h1 ? _GEN_4375 : _GEN_9383; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10025 = unuse_way == 2'h1 ? _GEN_4376 : _GEN_9384; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10026 = unuse_way == 2'h1 ? _GEN_4377 : _GEN_9385; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10027 = unuse_way == 2'h1 ? _GEN_4378 : _GEN_9386; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10028 = unuse_way == 2'h1 ? _GEN_4379 : _GEN_9387; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10029 = unuse_way == 2'h1 ? _GEN_4380 : _GEN_9388; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10030 = unuse_way == 2'h1 ? _GEN_4381 : _GEN_9389; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10031 = unuse_way == 2'h1 ? _GEN_4382 : _GEN_9390; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10032 = unuse_way == 2'h1 ? _GEN_4383 : _GEN_9391; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10033 = unuse_way == 2'h1 ? _GEN_4384 : _GEN_9392; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10034 = unuse_way == 2'h1 ? _GEN_4385 : _GEN_9393; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10035 = unuse_way == 2'h1 ? _GEN_4386 : _GEN_9394; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10036 = unuse_way == 2'h1 ? _GEN_4387 : _GEN_9395; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10037 = unuse_way == 2'h1 ? _GEN_4388 : _GEN_9396; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10038 = unuse_way == 2'h1 ? _GEN_4389 : _GEN_9397; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10039 = unuse_way == 2'h1 ? _GEN_4390 : _GEN_9398; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10040 = unuse_way == 2'h1 ? _GEN_4391 : _GEN_9399; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10041 = unuse_way == 2'h1 ? _GEN_4392 : _GEN_9400; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10042 = unuse_way == 2'h1 ? _GEN_4393 : _GEN_9401; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10043 = unuse_way == 2'h1 ? _GEN_4394 : _GEN_9402; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10044 = unuse_way == 2'h1 ? _GEN_4395 : _GEN_9403; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10045 = unuse_way == 2'h1 ? _GEN_4396 : _GEN_9404; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10046 = unuse_way == 2'h1 ? _GEN_4397 : _GEN_9405; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10047 = unuse_way == 2'h1 ? _GEN_4398 : _GEN_9406; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10048 = unuse_way == 2'h1 ? _GEN_4399 : _GEN_9407; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10049 = unuse_way == 2'h1 ? _GEN_4400 : _GEN_9408; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10050 = unuse_way == 2'h1 ? _GEN_4401 : _GEN_9409; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10051 = unuse_way == 2'h1 ? _GEN_4402 : _GEN_9410; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10052 = unuse_way == 2'h1 ? _GEN_4403 : _GEN_9411; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10053 = unuse_way == 2'h1 ? _GEN_4404 : _GEN_9412; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10054 = unuse_way == 2'h1 ? _GEN_4405 : _GEN_9413; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10055 = unuse_way == 2'h1 ? _GEN_4406 : _GEN_9414; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10056 = unuse_way == 2'h1 ? _GEN_4407 : _GEN_9415; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10057 = unuse_way == 2'h1 ? _GEN_4408 : _GEN_9416; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10058 = unuse_way == 2'h1 ? _GEN_4409 : _GEN_9417; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10059 = unuse_way == 2'h1 ? _GEN_4410 : _GEN_9418; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10060 = unuse_way == 2'h1 ? _GEN_4411 : _GEN_9419; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10061 = unuse_way == 2'h1 ? _GEN_4412 : _GEN_9420; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10062 = unuse_way == 2'h1 ? _GEN_4413 : _GEN_9421; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10063 = unuse_way == 2'h1 ? _GEN_4414 : _GEN_9422; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10064 = unuse_way == 2'h1 ? _GEN_4415 : _GEN_9423; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10065 = unuse_way == 2'h1 ? _GEN_4416 : _GEN_9424; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10066 = unuse_way == 2'h1 ? _GEN_4417 : _GEN_9425; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10067 = unuse_way == 2'h1 ? _GEN_4418 : _GEN_9426; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10068 = unuse_way == 2'h1 ? _GEN_4419 : _GEN_9427; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10069 = unuse_way == 2'h1 ? _GEN_4420 : _GEN_9428; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10070 = unuse_way == 2'h1 ? _GEN_4421 : _GEN_9429; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10071 = unuse_way == 2'h1 ? _GEN_4422 : _GEN_9430; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10072 = unuse_way == 2'h1 ? _GEN_4423 : _GEN_9431; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10073 = unuse_way == 2'h1 ? _GEN_4424 : _GEN_9432; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10074 = unuse_way == 2'h1 ? _GEN_4425 : _GEN_9433; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10075 = unuse_way == 2'h1 ? _GEN_4426 : _GEN_9434; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10076 = unuse_way == 2'h1 ? _GEN_4427 : _GEN_9435; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10077 = unuse_way == 2'h1 ? _GEN_4428 : _GEN_9436; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10078 = unuse_way == 2'h1 ? _GEN_4429 : _GEN_9437; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10079 = unuse_way == 2'h1 ? _GEN_4430 : _GEN_9438; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10080 = unuse_way == 2'h1 ? _GEN_4431 : _GEN_9439; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10081 = unuse_way == 2'h1 ? _GEN_4432 : _GEN_9440; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10082 = unuse_way == 2'h1 ? _GEN_4433 : _GEN_9441; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10083 = unuse_way == 2'h1 ? _GEN_4434 : _GEN_9442; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10084 = unuse_way == 2'h1 ? _GEN_4435 : _GEN_9443; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10085 = unuse_way == 2'h1 ? _GEN_4436 : _GEN_9444; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10086 = unuse_way == 2'h1 ? _GEN_4437 : _GEN_9445; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10087 = unuse_way == 2'h1 ? _GEN_4438 : _GEN_9446; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10088 = unuse_way == 2'h1 ? _GEN_4439 : _GEN_9447; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10089 = unuse_way == 2'h1 ? _GEN_4440 : _GEN_9448; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10090 = unuse_way == 2'h1 ? _GEN_4441 : _GEN_9449; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10091 = unuse_way == 2'h1 ? _GEN_4442 : _GEN_9450; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10092 = unuse_way == 2'h1 ? _GEN_4443 : _GEN_9451; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10093 = unuse_way == 2'h1 ? _GEN_4444 : _GEN_9452; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10094 = unuse_way == 2'h1 ? _GEN_4445 : _GEN_9453; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10095 = unuse_way == 2'h1 ? _GEN_4446 : _GEN_9454; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10096 = unuse_way == 2'h1 ? _GEN_4447 : _GEN_9455; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10097 = unuse_way == 2'h1 ? _GEN_4448 : _GEN_9456; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10098 = unuse_way == 2'h1 ? _GEN_4449 : _GEN_9457; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10099 = unuse_way == 2'h1 ? _GEN_4450 : _GEN_9458; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10100 = unuse_way == 2'h1 ? _GEN_4451 : _GEN_9459; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10101 = unuse_way == 2'h1 ? _GEN_4452 : _GEN_9460; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10102 = unuse_way == 2'h1 ? _GEN_4453 : _GEN_9461; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10103 = unuse_way == 2'h1 ? _GEN_4454 : _GEN_9462; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10104 = unuse_way == 2'h1 ? _GEN_4455 : _GEN_9463; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10105 = unuse_way == 2'h1 ? _GEN_4456 : _GEN_9464; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10106 = unuse_way == 2'h1 ? _GEN_4457 : _GEN_9465; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10107 = unuse_way == 2'h1 ? _GEN_4458 : _GEN_9466; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10108 = unuse_way == 2'h1 ? _GEN_4459 : _GEN_9467; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10109 = unuse_way == 2'h1 ? _GEN_4460 : _GEN_9468; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10110 = unuse_way == 2'h1 ? _GEN_4461 : _GEN_9469; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10111 = unuse_way == 2'h1 ? _GEN_4462 : _GEN_9470; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10112 = unuse_way == 2'h1 ? _GEN_4463 : _GEN_9471; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10113 = unuse_way == 2'h1 ? _GEN_4464 : _GEN_9472; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10114 = unuse_way == 2'h1 ? _GEN_4465 : _GEN_9473; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10115 = unuse_way == 2'h1 ? _GEN_4466 : _GEN_9474; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10116 = unuse_way == 2'h1 ? _GEN_4467 : _GEN_9475; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10117 = unuse_way == 2'h1 ? _GEN_4468 : _GEN_9476; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10118 = unuse_way == 2'h1 ? _GEN_4469 : _GEN_9477; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10119 = unuse_way == 2'h1 ? _GEN_4470 : _GEN_9478; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10120 = unuse_way == 2'h1 ? _GEN_4471 : _GEN_9479; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10121 = unuse_way == 2'h1 ? _GEN_4472 : _GEN_9480; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10122 = unuse_way == 2'h1 ? _GEN_4473 : _GEN_9481; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10123 = unuse_way == 2'h1 ? _GEN_4474 : _GEN_9482; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10124 = unuse_way == 2'h1 ? _GEN_4475 : _GEN_9483; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10125 = unuse_way == 2'h1 ? _GEN_4476 : _GEN_9484; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10126 = unuse_way == 2'h1 ? _GEN_4477 : _GEN_9485; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10127 = unuse_way == 2'h1 ? _GEN_4478 : _GEN_9486; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10128 = unuse_way == 2'h1 ? _GEN_4479 : _GEN_9487; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10129 = unuse_way == 2'h1 ? _GEN_4480 : _GEN_9488; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10130 = unuse_way == 2'h1 ? _GEN_4481 : _GEN_9489; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10131 = unuse_way == 2'h1 ? _GEN_4482 : _GEN_9490; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10132 = unuse_way == 2'h1 ? _GEN_4483 : _GEN_9491; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10133 = unuse_way == 2'h1 ? _GEN_4484 : _GEN_9492; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10134 = unuse_way == 2'h1 ? _GEN_4485 : _GEN_9493; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10135 = unuse_way == 2'h1 ? _GEN_4486 : _GEN_9494; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10136 = unuse_way == 2'h1 ? _GEN_4487 : _GEN_9495; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10137 = unuse_way == 2'h1 ? _GEN_4488 : _GEN_9496; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10138 = unuse_way == 2'h1 ? _GEN_4489 : _GEN_9497; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10139 = unuse_way == 2'h1 ? _GEN_4490 : _GEN_9498; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10140 = unuse_way == 2'h1 ? _GEN_4491 : _GEN_9499; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10141 = unuse_way == 2'h1 ? _GEN_4492 : _GEN_9500; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_10142 = unuse_way == 2'h1 ? _GEN_4493 : _GEN_9501; // @[d_cache.scala 150:34]
  wire  _GEN_10143 = unuse_way == 2'h1 ? _GEN_4494 : _GEN_9630; // @[d_cache.scala 150:34]
  wire  _GEN_10144 = unuse_way == 2'h1 ? _GEN_4495 : _GEN_9631; // @[d_cache.scala 150:34]
  wire  _GEN_10145 = unuse_way == 2'h1 ? _GEN_4496 : _GEN_9632; // @[d_cache.scala 150:34]
  wire  _GEN_10146 = unuse_way == 2'h1 ? _GEN_4497 : _GEN_9633; // @[d_cache.scala 150:34]
  wire  _GEN_10147 = unuse_way == 2'h1 ? _GEN_4498 : _GEN_9634; // @[d_cache.scala 150:34]
  wire  _GEN_10148 = unuse_way == 2'h1 ? _GEN_4499 : _GEN_9635; // @[d_cache.scala 150:34]
  wire  _GEN_10149 = unuse_way == 2'h1 ? _GEN_4500 : _GEN_9636; // @[d_cache.scala 150:34]
  wire  _GEN_10150 = unuse_way == 2'h1 ? _GEN_4501 : _GEN_9637; // @[d_cache.scala 150:34]
  wire  _GEN_10151 = unuse_way == 2'h1 ? _GEN_4502 : _GEN_9638; // @[d_cache.scala 150:34]
  wire  _GEN_10152 = unuse_way == 2'h1 ? _GEN_4503 : _GEN_9639; // @[d_cache.scala 150:34]
  wire  _GEN_10153 = unuse_way == 2'h1 ? _GEN_4504 : _GEN_9640; // @[d_cache.scala 150:34]
  wire  _GEN_10154 = unuse_way == 2'h1 ? _GEN_4505 : _GEN_9641; // @[d_cache.scala 150:34]
  wire  _GEN_10155 = unuse_way == 2'h1 ? _GEN_4506 : _GEN_9642; // @[d_cache.scala 150:34]
  wire  _GEN_10156 = unuse_way == 2'h1 ? _GEN_4507 : _GEN_9643; // @[d_cache.scala 150:34]
  wire  _GEN_10157 = unuse_way == 2'h1 ? _GEN_4508 : _GEN_9644; // @[d_cache.scala 150:34]
  wire  _GEN_10158 = unuse_way == 2'h1 ? _GEN_4509 : _GEN_9645; // @[d_cache.scala 150:34]
  wire  _GEN_10159 = unuse_way == 2'h1 ? _GEN_4510 : _GEN_9646; // @[d_cache.scala 150:34]
  wire  _GEN_10160 = unuse_way == 2'h1 ? _GEN_4511 : _GEN_9647; // @[d_cache.scala 150:34]
  wire  _GEN_10161 = unuse_way == 2'h1 ? _GEN_4512 : _GEN_9648; // @[d_cache.scala 150:34]
  wire  _GEN_10162 = unuse_way == 2'h1 ? _GEN_4513 : _GEN_9649; // @[d_cache.scala 150:34]
  wire  _GEN_10163 = unuse_way == 2'h1 ? _GEN_4514 : _GEN_9650; // @[d_cache.scala 150:34]
  wire  _GEN_10164 = unuse_way == 2'h1 ? _GEN_4515 : _GEN_9651; // @[d_cache.scala 150:34]
  wire  _GEN_10165 = unuse_way == 2'h1 ? _GEN_4516 : _GEN_9652; // @[d_cache.scala 150:34]
  wire  _GEN_10166 = unuse_way == 2'h1 ? _GEN_4517 : _GEN_9653; // @[d_cache.scala 150:34]
  wire  _GEN_10167 = unuse_way == 2'h1 ? _GEN_4518 : _GEN_9654; // @[d_cache.scala 150:34]
  wire  _GEN_10168 = unuse_way == 2'h1 ? _GEN_4519 : _GEN_9655; // @[d_cache.scala 150:34]
  wire  _GEN_10169 = unuse_way == 2'h1 ? _GEN_4520 : _GEN_9656; // @[d_cache.scala 150:34]
  wire  _GEN_10170 = unuse_way == 2'h1 ? _GEN_4521 : _GEN_9657; // @[d_cache.scala 150:34]
  wire  _GEN_10171 = unuse_way == 2'h1 ? _GEN_4522 : _GEN_9658; // @[d_cache.scala 150:34]
  wire  _GEN_10172 = unuse_way == 2'h1 ? _GEN_4523 : _GEN_9659; // @[d_cache.scala 150:34]
  wire  _GEN_10173 = unuse_way == 2'h1 ? _GEN_4524 : _GEN_9660; // @[d_cache.scala 150:34]
  wire  _GEN_10174 = unuse_way == 2'h1 ? _GEN_4525 : _GEN_9661; // @[d_cache.scala 150:34]
  wire  _GEN_10175 = unuse_way == 2'h1 ? _GEN_4526 : _GEN_9662; // @[d_cache.scala 150:34]
  wire  _GEN_10176 = unuse_way == 2'h1 ? _GEN_4527 : _GEN_9663; // @[d_cache.scala 150:34]
  wire  _GEN_10177 = unuse_way == 2'h1 ? _GEN_4528 : _GEN_9664; // @[d_cache.scala 150:34]
  wire  _GEN_10178 = unuse_way == 2'h1 ? _GEN_4529 : _GEN_9665; // @[d_cache.scala 150:34]
  wire  _GEN_10179 = unuse_way == 2'h1 ? _GEN_4530 : _GEN_9666; // @[d_cache.scala 150:34]
  wire  _GEN_10180 = unuse_way == 2'h1 ? _GEN_4531 : _GEN_9667; // @[d_cache.scala 150:34]
  wire  _GEN_10181 = unuse_way == 2'h1 ? _GEN_4532 : _GEN_9668; // @[d_cache.scala 150:34]
  wire  _GEN_10182 = unuse_way == 2'h1 ? _GEN_4533 : _GEN_9669; // @[d_cache.scala 150:34]
  wire  _GEN_10183 = unuse_way == 2'h1 ? _GEN_4534 : _GEN_9670; // @[d_cache.scala 150:34]
  wire  _GEN_10184 = unuse_way == 2'h1 ? _GEN_4535 : _GEN_9671; // @[d_cache.scala 150:34]
  wire  _GEN_10185 = unuse_way == 2'h1 ? _GEN_4536 : _GEN_9672; // @[d_cache.scala 150:34]
  wire  _GEN_10186 = unuse_way == 2'h1 ? _GEN_4537 : _GEN_9673; // @[d_cache.scala 150:34]
  wire  _GEN_10187 = unuse_way == 2'h1 ? _GEN_4538 : _GEN_9674; // @[d_cache.scala 150:34]
  wire  _GEN_10188 = unuse_way == 2'h1 ? _GEN_4539 : _GEN_9675; // @[d_cache.scala 150:34]
  wire  _GEN_10189 = unuse_way == 2'h1 ? _GEN_4540 : _GEN_9676; // @[d_cache.scala 150:34]
  wire  _GEN_10190 = unuse_way == 2'h1 ? _GEN_4541 : _GEN_9677; // @[d_cache.scala 150:34]
  wire  _GEN_10191 = unuse_way == 2'h1 ? _GEN_4542 : _GEN_9678; // @[d_cache.scala 150:34]
  wire  _GEN_10192 = unuse_way == 2'h1 ? _GEN_4543 : _GEN_9679; // @[d_cache.scala 150:34]
  wire  _GEN_10193 = unuse_way == 2'h1 ? _GEN_4544 : _GEN_9680; // @[d_cache.scala 150:34]
  wire  _GEN_10194 = unuse_way == 2'h1 ? _GEN_4545 : _GEN_9681; // @[d_cache.scala 150:34]
  wire  _GEN_10195 = unuse_way == 2'h1 ? _GEN_4546 : _GEN_9682; // @[d_cache.scala 150:34]
  wire  _GEN_10196 = unuse_way == 2'h1 ? _GEN_4547 : _GEN_9683; // @[d_cache.scala 150:34]
  wire  _GEN_10197 = unuse_way == 2'h1 ? _GEN_4548 : _GEN_9684; // @[d_cache.scala 150:34]
  wire  _GEN_10198 = unuse_way == 2'h1 ? _GEN_4549 : _GEN_9685; // @[d_cache.scala 150:34]
  wire  _GEN_10199 = unuse_way == 2'h1 ? _GEN_4550 : _GEN_9686; // @[d_cache.scala 150:34]
  wire  _GEN_10200 = unuse_way == 2'h1 ? _GEN_4551 : _GEN_9687; // @[d_cache.scala 150:34]
  wire  _GEN_10201 = unuse_way == 2'h1 ? _GEN_4552 : _GEN_9688; // @[d_cache.scala 150:34]
  wire  _GEN_10202 = unuse_way == 2'h1 ? _GEN_4553 : _GEN_9689; // @[d_cache.scala 150:34]
  wire  _GEN_10203 = unuse_way == 2'h1 ? _GEN_4554 : _GEN_9690; // @[d_cache.scala 150:34]
  wire  _GEN_10204 = unuse_way == 2'h1 ? _GEN_4555 : _GEN_9691; // @[d_cache.scala 150:34]
  wire  _GEN_10205 = unuse_way == 2'h1 ? _GEN_4556 : _GEN_9692; // @[d_cache.scala 150:34]
  wire  _GEN_10206 = unuse_way == 2'h1 ? _GEN_4557 : _GEN_9693; // @[d_cache.scala 150:34]
  wire  _GEN_10207 = unuse_way == 2'h1 ? _GEN_4558 : _GEN_9694; // @[d_cache.scala 150:34]
  wire  _GEN_10208 = unuse_way == 2'h1 ? _GEN_4559 : _GEN_9695; // @[d_cache.scala 150:34]
  wire  _GEN_10209 = unuse_way == 2'h1 ? _GEN_4560 : _GEN_9696; // @[d_cache.scala 150:34]
  wire  _GEN_10210 = unuse_way == 2'h1 ? _GEN_4561 : _GEN_9697; // @[d_cache.scala 150:34]
  wire  _GEN_10211 = unuse_way == 2'h1 ? _GEN_4562 : _GEN_9698; // @[d_cache.scala 150:34]
  wire  _GEN_10212 = unuse_way == 2'h1 ? _GEN_4563 : _GEN_9699; // @[d_cache.scala 150:34]
  wire  _GEN_10213 = unuse_way == 2'h1 ? _GEN_4564 : _GEN_9700; // @[d_cache.scala 150:34]
  wire  _GEN_10214 = unuse_way == 2'h1 ? _GEN_4565 : _GEN_9701; // @[d_cache.scala 150:34]
  wire  _GEN_10215 = unuse_way == 2'h1 ? _GEN_4566 : _GEN_9702; // @[d_cache.scala 150:34]
  wire  _GEN_10216 = unuse_way == 2'h1 ? _GEN_4567 : _GEN_9703; // @[d_cache.scala 150:34]
  wire  _GEN_10217 = unuse_way == 2'h1 ? _GEN_4568 : _GEN_9704; // @[d_cache.scala 150:34]
  wire  _GEN_10218 = unuse_way == 2'h1 ? _GEN_4569 : _GEN_9705; // @[d_cache.scala 150:34]
  wire  _GEN_10219 = unuse_way == 2'h1 ? _GEN_4570 : _GEN_9706; // @[d_cache.scala 150:34]
  wire  _GEN_10220 = unuse_way == 2'h1 ? _GEN_4571 : _GEN_9707; // @[d_cache.scala 150:34]
  wire  _GEN_10221 = unuse_way == 2'h1 ? _GEN_4572 : _GEN_9708; // @[d_cache.scala 150:34]
  wire  _GEN_10222 = unuse_way == 2'h1 ? _GEN_4573 : _GEN_9709; // @[d_cache.scala 150:34]
  wire  _GEN_10223 = unuse_way == 2'h1 ? _GEN_4574 : _GEN_9710; // @[d_cache.scala 150:34]
  wire  _GEN_10224 = unuse_way == 2'h1 ? _GEN_4575 : _GEN_9711; // @[d_cache.scala 150:34]
  wire  _GEN_10225 = unuse_way == 2'h1 ? _GEN_4576 : _GEN_9712; // @[d_cache.scala 150:34]
  wire  _GEN_10226 = unuse_way == 2'h1 ? _GEN_4577 : _GEN_9713; // @[d_cache.scala 150:34]
  wire  _GEN_10227 = unuse_way == 2'h1 ? _GEN_4578 : _GEN_9714; // @[d_cache.scala 150:34]
  wire  _GEN_10228 = unuse_way == 2'h1 ? _GEN_4579 : _GEN_9715; // @[d_cache.scala 150:34]
  wire  _GEN_10229 = unuse_way == 2'h1 ? _GEN_4580 : _GEN_9716; // @[d_cache.scala 150:34]
  wire  _GEN_10230 = unuse_way == 2'h1 ? _GEN_4581 : _GEN_9717; // @[d_cache.scala 150:34]
  wire  _GEN_10231 = unuse_way == 2'h1 ? _GEN_4582 : _GEN_9718; // @[d_cache.scala 150:34]
  wire  _GEN_10232 = unuse_way == 2'h1 ? _GEN_4583 : _GEN_9719; // @[d_cache.scala 150:34]
  wire  _GEN_10233 = unuse_way == 2'h1 ? _GEN_4584 : _GEN_9720; // @[d_cache.scala 150:34]
  wire  _GEN_10234 = unuse_way == 2'h1 ? _GEN_4585 : _GEN_9721; // @[d_cache.scala 150:34]
  wire  _GEN_10235 = unuse_way == 2'h1 ? _GEN_4586 : _GEN_9722; // @[d_cache.scala 150:34]
  wire  _GEN_10236 = unuse_way == 2'h1 ? _GEN_4587 : _GEN_9723; // @[d_cache.scala 150:34]
  wire  _GEN_10237 = unuse_way == 2'h1 ? _GEN_4588 : _GEN_9724; // @[d_cache.scala 150:34]
  wire  _GEN_10238 = unuse_way == 2'h1 ? _GEN_4589 : _GEN_9725; // @[d_cache.scala 150:34]
  wire  _GEN_10239 = unuse_way == 2'h1 ? _GEN_4590 : _GEN_9726; // @[d_cache.scala 150:34]
  wire  _GEN_10240 = unuse_way == 2'h1 ? _GEN_4591 : _GEN_9727; // @[d_cache.scala 150:34]
  wire  _GEN_10241 = unuse_way == 2'h1 ? _GEN_4592 : _GEN_9728; // @[d_cache.scala 150:34]
  wire  _GEN_10242 = unuse_way == 2'h1 ? _GEN_4593 : _GEN_9729; // @[d_cache.scala 150:34]
  wire  _GEN_10243 = unuse_way == 2'h1 ? _GEN_4594 : _GEN_9730; // @[d_cache.scala 150:34]
  wire  _GEN_10244 = unuse_way == 2'h1 ? _GEN_4595 : _GEN_9731; // @[d_cache.scala 150:34]
  wire  _GEN_10245 = unuse_way == 2'h1 ? _GEN_4596 : _GEN_9732; // @[d_cache.scala 150:34]
  wire  _GEN_10246 = unuse_way == 2'h1 ? _GEN_4597 : _GEN_9733; // @[d_cache.scala 150:34]
  wire  _GEN_10247 = unuse_way == 2'h1 ? _GEN_4598 : _GEN_9734; // @[d_cache.scala 150:34]
  wire  _GEN_10248 = unuse_way == 2'h1 ? _GEN_4599 : _GEN_9735; // @[d_cache.scala 150:34]
  wire  _GEN_10249 = unuse_way == 2'h1 ? _GEN_4600 : _GEN_9736; // @[d_cache.scala 150:34]
  wire  _GEN_10250 = unuse_way == 2'h1 ? _GEN_4601 : _GEN_9737; // @[d_cache.scala 150:34]
  wire  _GEN_10251 = unuse_way == 2'h1 ? _GEN_4602 : _GEN_9738; // @[d_cache.scala 150:34]
  wire  _GEN_10252 = unuse_way == 2'h1 ? _GEN_4603 : _GEN_9739; // @[d_cache.scala 150:34]
  wire  _GEN_10253 = unuse_way == 2'h1 ? _GEN_4604 : _GEN_9740; // @[d_cache.scala 150:34]
  wire  _GEN_10254 = unuse_way == 2'h1 ? _GEN_4605 : _GEN_9741; // @[d_cache.scala 150:34]
  wire  _GEN_10255 = unuse_way == 2'h1 ? _GEN_4606 : _GEN_9742; // @[d_cache.scala 150:34]
  wire  _GEN_10256 = unuse_way == 2'h1 ? _GEN_4607 : _GEN_9743; // @[d_cache.scala 150:34]
  wire  _GEN_10257 = unuse_way == 2'h1 ? _GEN_4608 : _GEN_9744; // @[d_cache.scala 150:34]
  wire  _GEN_10258 = unuse_way == 2'h1 ? _GEN_4609 : _GEN_9745; // @[d_cache.scala 150:34]
  wire  _GEN_10259 = unuse_way == 2'h1 ? _GEN_4610 : _GEN_9746; // @[d_cache.scala 150:34]
  wire  _GEN_10260 = unuse_way == 2'h1 ? _GEN_4611 : _GEN_9747; // @[d_cache.scala 150:34]
  wire  _GEN_10261 = unuse_way == 2'h1 ? _GEN_4612 : _GEN_9748; // @[d_cache.scala 150:34]
  wire  _GEN_10262 = unuse_way == 2'h1 ? _GEN_4613 : _GEN_9749; // @[d_cache.scala 150:34]
  wire  _GEN_10263 = unuse_way == 2'h1 ? _GEN_4614 : _GEN_9750; // @[d_cache.scala 150:34]
  wire  _GEN_10264 = unuse_way == 2'h1 ? _GEN_4615 : _GEN_9751; // @[d_cache.scala 150:34]
  wire  _GEN_10265 = unuse_way == 2'h1 ? _GEN_4616 : _GEN_9752; // @[d_cache.scala 150:34]
  wire  _GEN_10266 = unuse_way == 2'h1 ? _GEN_4617 : _GEN_9753; // @[d_cache.scala 150:34]
  wire  _GEN_10267 = unuse_way == 2'h1 ? _GEN_4618 : _GEN_9754; // @[d_cache.scala 150:34]
  wire  _GEN_10268 = unuse_way == 2'h1 ? _GEN_4619 : _GEN_9755; // @[d_cache.scala 150:34]
  wire  _GEN_10269 = unuse_way == 2'h1 ? _GEN_4620 : _GEN_9756; // @[d_cache.scala 150:34]
  wire  _GEN_10270 = unuse_way == 2'h1 ? _GEN_4621 : _GEN_9757; // @[d_cache.scala 150:34]
  wire  _GEN_10271 = unuse_way == 2'h1 | _GEN_9243; // @[d_cache.scala 150:34 155:23]
  wire [63:0] _GEN_10272 = unuse_way == 2'h1 ? ram_1_0 : _GEN_8859; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10273 = unuse_way == 2'h1 ? ram_1_1 : _GEN_8860; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10274 = unuse_way == 2'h1 ? ram_1_2 : _GEN_8861; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10275 = unuse_way == 2'h1 ? ram_1_3 : _GEN_8862; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10276 = unuse_way == 2'h1 ? ram_1_4 : _GEN_8863; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10277 = unuse_way == 2'h1 ? ram_1_5 : _GEN_8864; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10278 = unuse_way == 2'h1 ? ram_1_6 : _GEN_8865; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10279 = unuse_way == 2'h1 ? ram_1_7 : _GEN_8866; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10280 = unuse_way == 2'h1 ? ram_1_8 : _GEN_8867; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10281 = unuse_way == 2'h1 ? ram_1_9 : _GEN_8868; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10282 = unuse_way == 2'h1 ? ram_1_10 : _GEN_8869; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10283 = unuse_way == 2'h1 ? ram_1_11 : _GEN_8870; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10284 = unuse_way == 2'h1 ? ram_1_12 : _GEN_8871; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10285 = unuse_way == 2'h1 ? ram_1_13 : _GEN_8872; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10286 = unuse_way == 2'h1 ? ram_1_14 : _GEN_8873; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10287 = unuse_way == 2'h1 ? ram_1_15 : _GEN_8874; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10288 = unuse_way == 2'h1 ? ram_1_16 : _GEN_8875; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10289 = unuse_way == 2'h1 ? ram_1_17 : _GEN_8876; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10290 = unuse_way == 2'h1 ? ram_1_18 : _GEN_8877; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10291 = unuse_way == 2'h1 ? ram_1_19 : _GEN_8878; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10292 = unuse_way == 2'h1 ? ram_1_20 : _GEN_8879; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10293 = unuse_way == 2'h1 ? ram_1_21 : _GEN_8880; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10294 = unuse_way == 2'h1 ? ram_1_22 : _GEN_8881; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10295 = unuse_way == 2'h1 ? ram_1_23 : _GEN_8882; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10296 = unuse_way == 2'h1 ? ram_1_24 : _GEN_8883; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10297 = unuse_way == 2'h1 ? ram_1_25 : _GEN_8884; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10298 = unuse_way == 2'h1 ? ram_1_26 : _GEN_8885; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10299 = unuse_way == 2'h1 ? ram_1_27 : _GEN_8886; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10300 = unuse_way == 2'h1 ? ram_1_28 : _GEN_8887; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10301 = unuse_way == 2'h1 ? ram_1_29 : _GEN_8888; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10302 = unuse_way == 2'h1 ? ram_1_30 : _GEN_8889; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10303 = unuse_way == 2'h1 ? ram_1_31 : _GEN_8890; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10304 = unuse_way == 2'h1 ? ram_1_32 : _GEN_8891; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10305 = unuse_way == 2'h1 ? ram_1_33 : _GEN_8892; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10306 = unuse_way == 2'h1 ? ram_1_34 : _GEN_8893; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10307 = unuse_way == 2'h1 ? ram_1_35 : _GEN_8894; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10308 = unuse_way == 2'h1 ? ram_1_36 : _GEN_8895; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10309 = unuse_way == 2'h1 ? ram_1_37 : _GEN_8896; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10310 = unuse_way == 2'h1 ? ram_1_38 : _GEN_8897; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10311 = unuse_way == 2'h1 ? ram_1_39 : _GEN_8898; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10312 = unuse_way == 2'h1 ? ram_1_40 : _GEN_8899; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10313 = unuse_way == 2'h1 ? ram_1_41 : _GEN_8900; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10314 = unuse_way == 2'h1 ? ram_1_42 : _GEN_8901; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10315 = unuse_way == 2'h1 ? ram_1_43 : _GEN_8902; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10316 = unuse_way == 2'h1 ? ram_1_44 : _GEN_8903; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10317 = unuse_way == 2'h1 ? ram_1_45 : _GEN_8904; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10318 = unuse_way == 2'h1 ? ram_1_46 : _GEN_8905; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10319 = unuse_way == 2'h1 ? ram_1_47 : _GEN_8906; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10320 = unuse_way == 2'h1 ? ram_1_48 : _GEN_8907; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10321 = unuse_way == 2'h1 ? ram_1_49 : _GEN_8908; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10322 = unuse_way == 2'h1 ? ram_1_50 : _GEN_8909; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10323 = unuse_way == 2'h1 ? ram_1_51 : _GEN_8910; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10324 = unuse_way == 2'h1 ? ram_1_52 : _GEN_8911; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10325 = unuse_way == 2'h1 ? ram_1_53 : _GEN_8912; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10326 = unuse_way == 2'h1 ? ram_1_54 : _GEN_8913; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10327 = unuse_way == 2'h1 ? ram_1_55 : _GEN_8914; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10328 = unuse_way == 2'h1 ? ram_1_56 : _GEN_8915; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10329 = unuse_way == 2'h1 ? ram_1_57 : _GEN_8916; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10330 = unuse_way == 2'h1 ? ram_1_58 : _GEN_8917; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10331 = unuse_way == 2'h1 ? ram_1_59 : _GEN_8918; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10332 = unuse_way == 2'h1 ? ram_1_60 : _GEN_8919; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10333 = unuse_way == 2'h1 ? ram_1_61 : _GEN_8920; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10334 = unuse_way == 2'h1 ? ram_1_62 : _GEN_8921; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10335 = unuse_way == 2'h1 ? ram_1_63 : _GEN_8922; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10336 = unuse_way == 2'h1 ? ram_1_64 : _GEN_8923; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10337 = unuse_way == 2'h1 ? ram_1_65 : _GEN_8924; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10338 = unuse_way == 2'h1 ? ram_1_66 : _GEN_8925; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10339 = unuse_way == 2'h1 ? ram_1_67 : _GEN_8926; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10340 = unuse_way == 2'h1 ? ram_1_68 : _GEN_8927; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10341 = unuse_way == 2'h1 ? ram_1_69 : _GEN_8928; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10342 = unuse_way == 2'h1 ? ram_1_70 : _GEN_8929; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10343 = unuse_way == 2'h1 ? ram_1_71 : _GEN_8930; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10344 = unuse_way == 2'h1 ? ram_1_72 : _GEN_8931; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10345 = unuse_way == 2'h1 ? ram_1_73 : _GEN_8932; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10346 = unuse_way == 2'h1 ? ram_1_74 : _GEN_8933; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10347 = unuse_way == 2'h1 ? ram_1_75 : _GEN_8934; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10348 = unuse_way == 2'h1 ? ram_1_76 : _GEN_8935; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10349 = unuse_way == 2'h1 ? ram_1_77 : _GEN_8936; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10350 = unuse_way == 2'h1 ? ram_1_78 : _GEN_8937; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10351 = unuse_way == 2'h1 ? ram_1_79 : _GEN_8938; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10352 = unuse_way == 2'h1 ? ram_1_80 : _GEN_8939; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10353 = unuse_way == 2'h1 ? ram_1_81 : _GEN_8940; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10354 = unuse_way == 2'h1 ? ram_1_82 : _GEN_8941; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10355 = unuse_way == 2'h1 ? ram_1_83 : _GEN_8942; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10356 = unuse_way == 2'h1 ? ram_1_84 : _GEN_8943; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10357 = unuse_way == 2'h1 ? ram_1_85 : _GEN_8944; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10358 = unuse_way == 2'h1 ? ram_1_86 : _GEN_8945; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10359 = unuse_way == 2'h1 ? ram_1_87 : _GEN_8946; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10360 = unuse_way == 2'h1 ? ram_1_88 : _GEN_8947; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10361 = unuse_way == 2'h1 ? ram_1_89 : _GEN_8948; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10362 = unuse_way == 2'h1 ? ram_1_90 : _GEN_8949; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10363 = unuse_way == 2'h1 ? ram_1_91 : _GEN_8950; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10364 = unuse_way == 2'h1 ? ram_1_92 : _GEN_8951; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10365 = unuse_way == 2'h1 ? ram_1_93 : _GEN_8952; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10366 = unuse_way == 2'h1 ? ram_1_94 : _GEN_8953; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10367 = unuse_way == 2'h1 ? ram_1_95 : _GEN_8954; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10368 = unuse_way == 2'h1 ? ram_1_96 : _GEN_8955; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10369 = unuse_way == 2'h1 ? ram_1_97 : _GEN_8956; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10370 = unuse_way == 2'h1 ? ram_1_98 : _GEN_8957; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10371 = unuse_way == 2'h1 ? ram_1_99 : _GEN_8958; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10372 = unuse_way == 2'h1 ? ram_1_100 : _GEN_8959; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10373 = unuse_way == 2'h1 ? ram_1_101 : _GEN_8960; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10374 = unuse_way == 2'h1 ? ram_1_102 : _GEN_8961; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10375 = unuse_way == 2'h1 ? ram_1_103 : _GEN_8962; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10376 = unuse_way == 2'h1 ? ram_1_104 : _GEN_8963; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10377 = unuse_way == 2'h1 ? ram_1_105 : _GEN_8964; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10378 = unuse_way == 2'h1 ? ram_1_106 : _GEN_8965; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10379 = unuse_way == 2'h1 ? ram_1_107 : _GEN_8966; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10380 = unuse_way == 2'h1 ? ram_1_108 : _GEN_8967; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10381 = unuse_way == 2'h1 ? ram_1_109 : _GEN_8968; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10382 = unuse_way == 2'h1 ? ram_1_110 : _GEN_8969; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10383 = unuse_way == 2'h1 ? ram_1_111 : _GEN_8970; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10384 = unuse_way == 2'h1 ? ram_1_112 : _GEN_8971; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10385 = unuse_way == 2'h1 ? ram_1_113 : _GEN_8972; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10386 = unuse_way == 2'h1 ? ram_1_114 : _GEN_8973; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10387 = unuse_way == 2'h1 ? ram_1_115 : _GEN_8974; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10388 = unuse_way == 2'h1 ? ram_1_116 : _GEN_8975; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10389 = unuse_way == 2'h1 ? ram_1_117 : _GEN_8976; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10390 = unuse_way == 2'h1 ? ram_1_118 : _GEN_8977; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10391 = unuse_way == 2'h1 ? ram_1_119 : _GEN_8978; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10392 = unuse_way == 2'h1 ? ram_1_120 : _GEN_8979; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10393 = unuse_way == 2'h1 ? ram_1_121 : _GEN_8980; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10394 = unuse_way == 2'h1 ? ram_1_122 : _GEN_8981; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10395 = unuse_way == 2'h1 ? ram_1_123 : _GEN_8982; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10396 = unuse_way == 2'h1 ? ram_1_124 : _GEN_8983; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10397 = unuse_way == 2'h1 ? ram_1_125 : _GEN_8984; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10398 = unuse_way == 2'h1 ? ram_1_126 : _GEN_8985; // @[d_cache.scala 150:34 20:24]
  wire [63:0] _GEN_10399 = unuse_way == 2'h1 ? ram_1_127 : _GEN_8986; // @[d_cache.scala 150:34 20:24]
  wire [31:0] _GEN_10400 = unuse_way == 2'h1 ? tag_1_0 : _GEN_8987; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10401 = unuse_way == 2'h1 ? tag_1_1 : _GEN_8988; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10402 = unuse_way == 2'h1 ? tag_1_2 : _GEN_8989; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10403 = unuse_way == 2'h1 ? tag_1_3 : _GEN_8990; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10404 = unuse_way == 2'h1 ? tag_1_4 : _GEN_8991; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10405 = unuse_way == 2'h1 ? tag_1_5 : _GEN_8992; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10406 = unuse_way == 2'h1 ? tag_1_6 : _GEN_8993; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10407 = unuse_way == 2'h1 ? tag_1_7 : _GEN_8994; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10408 = unuse_way == 2'h1 ? tag_1_8 : _GEN_8995; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10409 = unuse_way == 2'h1 ? tag_1_9 : _GEN_8996; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10410 = unuse_way == 2'h1 ? tag_1_10 : _GEN_8997; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10411 = unuse_way == 2'h1 ? tag_1_11 : _GEN_8998; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10412 = unuse_way == 2'h1 ? tag_1_12 : _GEN_8999; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10413 = unuse_way == 2'h1 ? tag_1_13 : _GEN_9000; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10414 = unuse_way == 2'h1 ? tag_1_14 : _GEN_9001; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10415 = unuse_way == 2'h1 ? tag_1_15 : _GEN_9002; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10416 = unuse_way == 2'h1 ? tag_1_16 : _GEN_9003; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10417 = unuse_way == 2'h1 ? tag_1_17 : _GEN_9004; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10418 = unuse_way == 2'h1 ? tag_1_18 : _GEN_9005; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10419 = unuse_way == 2'h1 ? tag_1_19 : _GEN_9006; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10420 = unuse_way == 2'h1 ? tag_1_20 : _GEN_9007; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10421 = unuse_way == 2'h1 ? tag_1_21 : _GEN_9008; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10422 = unuse_way == 2'h1 ? tag_1_22 : _GEN_9009; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10423 = unuse_way == 2'h1 ? tag_1_23 : _GEN_9010; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10424 = unuse_way == 2'h1 ? tag_1_24 : _GEN_9011; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10425 = unuse_way == 2'h1 ? tag_1_25 : _GEN_9012; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10426 = unuse_way == 2'h1 ? tag_1_26 : _GEN_9013; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10427 = unuse_way == 2'h1 ? tag_1_27 : _GEN_9014; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10428 = unuse_way == 2'h1 ? tag_1_28 : _GEN_9015; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10429 = unuse_way == 2'h1 ? tag_1_29 : _GEN_9016; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10430 = unuse_way == 2'h1 ? tag_1_30 : _GEN_9017; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10431 = unuse_way == 2'h1 ? tag_1_31 : _GEN_9018; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10432 = unuse_way == 2'h1 ? tag_1_32 : _GEN_9019; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10433 = unuse_way == 2'h1 ? tag_1_33 : _GEN_9020; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10434 = unuse_way == 2'h1 ? tag_1_34 : _GEN_9021; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10435 = unuse_way == 2'h1 ? tag_1_35 : _GEN_9022; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10436 = unuse_way == 2'h1 ? tag_1_36 : _GEN_9023; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10437 = unuse_way == 2'h1 ? tag_1_37 : _GEN_9024; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10438 = unuse_way == 2'h1 ? tag_1_38 : _GEN_9025; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10439 = unuse_way == 2'h1 ? tag_1_39 : _GEN_9026; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10440 = unuse_way == 2'h1 ? tag_1_40 : _GEN_9027; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10441 = unuse_way == 2'h1 ? tag_1_41 : _GEN_9028; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10442 = unuse_way == 2'h1 ? tag_1_42 : _GEN_9029; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10443 = unuse_way == 2'h1 ? tag_1_43 : _GEN_9030; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10444 = unuse_way == 2'h1 ? tag_1_44 : _GEN_9031; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10445 = unuse_way == 2'h1 ? tag_1_45 : _GEN_9032; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10446 = unuse_way == 2'h1 ? tag_1_46 : _GEN_9033; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10447 = unuse_way == 2'h1 ? tag_1_47 : _GEN_9034; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10448 = unuse_way == 2'h1 ? tag_1_48 : _GEN_9035; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10449 = unuse_way == 2'h1 ? tag_1_49 : _GEN_9036; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10450 = unuse_way == 2'h1 ? tag_1_50 : _GEN_9037; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10451 = unuse_way == 2'h1 ? tag_1_51 : _GEN_9038; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10452 = unuse_way == 2'h1 ? tag_1_52 : _GEN_9039; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10453 = unuse_way == 2'h1 ? tag_1_53 : _GEN_9040; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10454 = unuse_way == 2'h1 ? tag_1_54 : _GEN_9041; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10455 = unuse_way == 2'h1 ? tag_1_55 : _GEN_9042; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10456 = unuse_way == 2'h1 ? tag_1_56 : _GEN_9043; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10457 = unuse_way == 2'h1 ? tag_1_57 : _GEN_9044; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10458 = unuse_way == 2'h1 ? tag_1_58 : _GEN_9045; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10459 = unuse_way == 2'h1 ? tag_1_59 : _GEN_9046; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10460 = unuse_way == 2'h1 ? tag_1_60 : _GEN_9047; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10461 = unuse_way == 2'h1 ? tag_1_61 : _GEN_9048; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10462 = unuse_way == 2'h1 ? tag_1_62 : _GEN_9049; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10463 = unuse_way == 2'h1 ? tag_1_63 : _GEN_9050; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10464 = unuse_way == 2'h1 ? tag_1_64 : _GEN_9051; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10465 = unuse_way == 2'h1 ? tag_1_65 : _GEN_9052; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10466 = unuse_way == 2'h1 ? tag_1_66 : _GEN_9053; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10467 = unuse_way == 2'h1 ? tag_1_67 : _GEN_9054; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10468 = unuse_way == 2'h1 ? tag_1_68 : _GEN_9055; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10469 = unuse_way == 2'h1 ? tag_1_69 : _GEN_9056; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10470 = unuse_way == 2'h1 ? tag_1_70 : _GEN_9057; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10471 = unuse_way == 2'h1 ? tag_1_71 : _GEN_9058; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10472 = unuse_way == 2'h1 ? tag_1_72 : _GEN_9059; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10473 = unuse_way == 2'h1 ? tag_1_73 : _GEN_9060; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10474 = unuse_way == 2'h1 ? tag_1_74 : _GEN_9061; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10475 = unuse_way == 2'h1 ? tag_1_75 : _GEN_9062; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10476 = unuse_way == 2'h1 ? tag_1_76 : _GEN_9063; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10477 = unuse_way == 2'h1 ? tag_1_77 : _GEN_9064; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10478 = unuse_way == 2'h1 ? tag_1_78 : _GEN_9065; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10479 = unuse_way == 2'h1 ? tag_1_79 : _GEN_9066; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10480 = unuse_way == 2'h1 ? tag_1_80 : _GEN_9067; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10481 = unuse_way == 2'h1 ? tag_1_81 : _GEN_9068; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10482 = unuse_way == 2'h1 ? tag_1_82 : _GEN_9069; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10483 = unuse_way == 2'h1 ? tag_1_83 : _GEN_9070; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10484 = unuse_way == 2'h1 ? tag_1_84 : _GEN_9071; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10485 = unuse_way == 2'h1 ? tag_1_85 : _GEN_9072; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10486 = unuse_way == 2'h1 ? tag_1_86 : _GEN_9073; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10487 = unuse_way == 2'h1 ? tag_1_87 : _GEN_9074; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10488 = unuse_way == 2'h1 ? tag_1_88 : _GEN_9075; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10489 = unuse_way == 2'h1 ? tag_1_89 : _GEN_9076; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10490 = unuse_way == 2'h1 ? tag_1_90 : _GEN_9077; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10491 = unuse_way == 2'h1 ? tag_1_91 : _GEN_9078; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10492 = unuse_way == 2'h1 ? tag_1_92 : _GEN_9079; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10493 = unuse_way == 2'h1 ? tag_1_93 : _GEN_9080; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10494 = unuse_way == 2'h1 ? tag_1_94 : _GEN_9081; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10495 = unuse_way == 2'h1 ? tag_1_95 : _GEN_9082; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10496 = unuse_way == 2'h1 ? tag_1_96 : _GEN_9083; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10497 = unuse_way == 2'h1 ? tag_1_97 : _GEN_9084; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10498 = unuse_way == 2'h1 ? tag_1_98 : _GEN_9085; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10499 = unuse_way == 2'h1 ? tag_1_99 : _GEN_9086; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10500 = unuse_way == 2'h1 ? tag_1_100 : _GEN_9087; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10501 = unuse_way == 2'h1 ? tag_1_101 : _GEN_9088; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10502 = unuse_way == 2'h1 ? tag_1_102 : _GEN_9089; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10503 = unuse_way == 2'h1 ? tag_1_103 : _GEN_9090; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10504 = unuse_way == 2'h1 ? tag_1_104 : _GEN_9091; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10505 = unuse_way == 2'h1 ? tag_1_105 : _GEN_9092; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10506 = unuse_way == 2'h1 ? tag_1_106 : _GEN_9093; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10507 = unuse_way == 2'h1 ? tag_1_107 : _GEN_9094; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10508 = unuse_way == 2'h1 ? tag_1_108 : _GEN_9095; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10509 = unuse_way == 2'h1 ? tag_1_109 : _GEN_9096; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10510 = unuse_way == 2'h1 ? tag_1_110 : _GEN_9097; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10511 = unuse_way == 2'h1 ? tag_1_111 : _GEN_9098; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10512 = unuse_way == 2'h1 ? tag_1_112 : _GEN_9099; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10513 = unuse_way == 2'h1 ? tag_1_113 : _GEN_9100; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10514 = unuse_way == 2'h1 ? tag_1_114 : _GEN_9101; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10515 = unuse_way == 2'h1 ? tag_1_115 : _GEN_9102; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10516 = unuse_way == 2'h1 ? tag_1_116 : _GEN_9103; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10517 = unuse_way == 2'h1 ? tag_1_117 : _GEN_9104; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10518 = unuse_way == 2'h1 ? tag_1_118 : _GEN_9105; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10519 = unuse_way == 2'h1 ? tag_1_119 : _GEN_9106; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10520 = unuse_way == 2'h1 ? tag_1_120 : _GEN_9107; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10521 = unuse_way == 2'h1 ? tag_1_121 : _GEN_9108; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10522 = unuse_way == 2'h1 ? tag_1_122 : _GEN_9109; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10523 = unuse_way == 2'h1 ? tag_1_123 : _GEN_9110; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10524 = unuse_way == 2'h1 ? tag_1_124 : _GEN_9111; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10525 = unuse_way == 2'h1 ? tag_1_125 : _GEN_9112; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10526 = unuse_way == 2'h1 ? tag_1_126 : _GEN_9113; // @[d_cache.scala 150:34 29:24]
  wire [31:0] _GEN_10527 = unuse_way == 2'h1 ? tag_1_127 : _GEN_9114; // @[d_cache.scala 150:34 29:24]
  wire  _GEN_10528 = unuse_way == 2'h1 ? valid_1_0 : _GEN_9115; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10529 = unuse_way == 2'h1 ? valid_1_1 : _GEN_9116; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10530 = unuse_way == 2'h1 ? valid_1_2 : _GEN_9117; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10531 = unuse_way == 2'h1 ? valid_1_3 : _GEN_9118; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10532 = unuse_way == 2'h1 ? valid_1_4 : _GEN_9119; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10533 = unuse_way == 2'h1 ? valid_1_5 : _GEN_9120; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10534 = unuse_way == 2'h1 ? valid_1_6 : _GEN_9121; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10535 = unuse_way == 2'h1 ? valid_1_7 : _GEN_9122; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10536 = unuse_way == 2'h1 ? valid_1_8 : _GEN_9123; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10537 = unuse_way == 2'h1 ? valid_1_9 : _GEN_9124; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10538 = unuse_way == 2'h1 ? valid_1_10 : _GEN_9125; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10539 = unuse_way == 2'h1 ? valid_1_11 : _GEN_9126; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10540 = unuse_way == 2'h1 ? valid_1_12 : _GEN_9127; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10541 = unuse_way == 2'h1 ? valid_1_13 : _GEN_9128; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10542 = unuse_way == 2'h1 ? valid_1_14 : _GEN_9129; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10543 = unuse_way == 2'h1 ? valid_1_15 : _GEN_9130; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10544 = unuse_way == 2'h1 ? valid_1_16 : _GEN_9131; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10545 = unuse_way == 2'h1 ? valid_1_17 : _GEN_9132; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10546 = unuse_way == 2'h1 ? valid_1_18 : _GEN_9133; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10547 = unuse_way == 2'h1 ? valid_1_19 : _GEN_9134; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10548 = unuse_way == 2'h1 ? valid_1_20 : _GEN_9135; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10549 = unuse_way == 2'h1 ? valid_1_21 : _GEN_9136; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10550 = unuse_way == 2'h1 ? valid_1_22 : _GEN_9137; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10551 = unuse_way == 2'h1 ? valid_1_23 : _GEN_9138; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10552 = unuse_way == 2'h1 ? valid_1_24 : _GEN_9139; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10553 = unuse_way == 2'h1 ? valid_1_25 : _GEN_9140; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10554 = unuse_way == 2'h1 ? valid_1_26 : _GEN_9141; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10555 = unuse_way == 2'h1 ? valid_1_27 : _GEN_9142; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10556 = unuse_way == 2'h1 ? valid_1_28 : _GEN_9143; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10557 = unuse_way == 2'h1 ? valid_1_29 : _GEN_9144; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10558 = unuse_way == 2'h1 ? valid_1_30 : _GEN_9145; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10559 = unuse_way == 2'h1 ? valid_1_31 : _GEN_9146; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10560 = unuse_way == 2'h1 ? valid_1_32 : _GEN_9147; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10561 = unuse_way == 2'h1 ? valid_1_33 : _GEN_9148; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10562 = unuse_way == 2'h1 ? valid_1_34 : _GEN_9149; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10563 = unuse_way == 2'h1 ? valid_1_35 : _GEN_9150; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10564 = unuse_way == 2'h1 ? valid_1_36 : _GEN_9151; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10565 = unuse_way == 2'h1 ? valid_1_37 : _GEN_9152; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10566 = unuse_way == 2'h1 ? valid_1_38 : _GEN_9153; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10567 = unuse_way == 2'h1 ? valid_1_39 : _GEN_9154; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10568 = unuse_way == 2'h1 ? valid_1_40 : _GEN_9155; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10569 = unuse_way == 2'h1 ? valid_1_41 : _GEN_9156; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10570 = unuse_way == 2'h1 ? valid_1_42 : _GEN_9157; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10571 = unuse_way == 2'h1 ? valid_1_43 : _GEN_9158; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10572 = unuse_way == 2'h1 ? valid_1_44 : _GEN_9159; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10573 = unuse_way == 2'h1 ? valid_1_45 : _GEN_9160; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10574 = unuse_way == 2'h1 ? valid_1_46 : _GEN_9161; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10575 = unuse_way == 2'h1 ? valid_1_47 : _GEN_9162; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10576 = unuse_way == 2'h1 ? valid_1_48 : _GEN_9163; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10577 = unuse_way == 2'h1 ? valid_1_49 : _GEN_9164; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10578 = unuse_way == 2'h1 ? valid_1_50 : _GEN_9165; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10579 = unuse_way == 2'h1 ? valid_1_51 : _GEN_9166; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10580 = unuse_way == 2'h1 ? valid_1_52 : _GEN_9167; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10581 = unuse_way == 2'h1 ? valid_1_53 : _GEN_9168; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10582 = unuse_way == 2'h1 ? valid_1_54 : _GEN_9169; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10583 = unuse_way == 2'h1 ? valid_1_55 : _GEN_9170; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10584 = unuse_way == 2'h1 ? valid_1_56 : _GEN_9171; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10585 = unuse_way == 2'h1 ? valid_1_57 : _GEN_9172; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10586 = unuse_way == 2'h1 ? valid_1_58 : _GEN_9173; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10587 = unuse_way == 2'h1 ? valid_1_59 : _GEN_9174; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10588 = unuse_way == 2'h1 ? valid_1_60 : _GEN_9175; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10589 = unuse_way == 2'h1 ? valid_1_61 : _GEN_9176; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10590 = unuse_way == 2'h1 ? valid_1_62 : _GEN_9177; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10591 = unuse_way == 2'h1 ? valid_1_63 : _GEN_9178; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10592 = unuse_way == 2'h1 ? valid_1_64 : _GEN_9179; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10593 = unuse_way == 2'h1 ? valid_1_65 : _GEN_9180; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10594 = unuse_way == 2'h1 ? valid_1_66 : _GEN_9181; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10595 = unuse_way == 2'h1 ? valid_1_67 : _GEN_9182; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10596 = unuse_way == 2'h1 ? valid_1_68 : _GEN_9183; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10597 = unuse_way == 2'h1 ? valid_1_69 : _GEN_9184; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10598 = unuse_way == 2'h1 ? valid_1_70 : _GEN_9185; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10599 = unuse_way == 2'h1 ? valid_1_71 : _GEN_9186; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10600 = unuse_way == 2'h1 ? valid_1_72 : _GEN_9187; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10601 = unuse_way == 2'h1 ? valid_1_73 : _GEN_9188; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10602 = unuse_way == 2'h1 ? valid_1_74 : _GEN_9189; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10603 = unuse_way == 2'h1 ? valid_1_75 : _GEN_9190; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10604 = unuse_way == 2'h1 ? valid_1_76 : _GEN_9191; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10605 = unuse_way == 2'h1 ? valid_1_77 : _GEN_9192; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10606 = unuse_way == 2'h1 ? valid_1_78 : _GEN_9193; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10607 = unuse_way == 2'h1 ? valid_1_79 : _GEN_9194; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10608 = unuse_way == 2'h1 ? valid_1_80 : _GEN_9195; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10609 = unuse_way == 2'h1 ? valid_1_81 : _GEN_9196; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10610 = unuse_way == 2'h1 ? valid_1_82 : _GEN_9197; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10611 = unuse_way == 2'h1 ? valid_1_83 : _GEN_9198; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10612 = unuse_way == 2'h1 ? valid_1_84 : _GEN_9199; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10613 = unuse_way == 2'h1 ? valid_1_85 : _GEN_9200; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10614 = unuse_way == 2'h1 ? valid_1_86 : _GEN_9201; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10615 = unuse_way == 2'h1 ? valid_1_87 : _GEN_9202; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10616 = unuse_way == 2'h1 ? valid_1_88 : _GEN_9203; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10617 = unuse_way == 2'h1 ? valid_1_89 : _GEN_9204; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10618 = unuse_way == 2'h1 ? valid_1_90 : _GEN_9205; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10619 = unuse_way == 2'h1 ? valid_1_91 : _GEN_9206; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10620 = unuse_way == 2'h1 ? valid_1_92 : _GEN_9207; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10621 = unuse_way == 2'h1 ? valid_1_93 : _GEN_9208; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10622 = unuse_way == 2'h1 ? valid_1_94 : _GEN_9209; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10623 = unuse_way == 2'h1 ? valid_1_95 : _GEN_9210; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10624 = unuse_way == 2'h1 ? valid_1_96 : _GEN_9211; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10625 = unuse_way == 2'h1 ? valid_1_97 : _GEN_9212; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10626 = unuse_way == 2'h1 ? valid_1_98 : _GEN_9213; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10627 = unuse_way == 2'h1 ? valid_1_99 : _GEN_9214; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10628 = unuse_way == 2'h1 ? valid_1_100 : _GEN_9215; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10629 = unuse_way == 2'h1 ? valid_1_101 : _GEN_9216; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10630 = unuse_way == 2'h1 ? valid_1_102 : _GEN_9217; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10631 = unuse_way == 2'h1 ? valid_1_103 : _GEN_9218; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10632 = unuse_way == 2'h1 ? valid_1_104 : _GEN_9219; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10633 = unuse_way == 2'h1 ? valid_1_105 : _GEN_9220; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10634 = unuse_way == 2'h1 ? valid_1_106 : _GEN_9221; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10635 = unuse_way == 2'h1 ? valid_1_107 : _GEN_9222; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10636 = unuse_way == 2'h1 ? valid_1_108 : _GEN_9223; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10637 = unuse_way == 2'h1 ? valid_1_109 : _GEN_9224; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10638 = unuse_way == 2'h1 ? valid_1_110 : _GEN_9225; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10639 = unuse_way == 2'h1 ? valid_1_111 : _GEN_9226; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10640 = unuse_way == 2'h1 ? valid_1_112 : _GEN_9227; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10641 = unuse_way == 2'h1 ? valid_1_113 : _GEN_9228; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10642 = unuse_way == 2'h1 ? valid_1_114 : _GEN_9229; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10643 = unuse_way == 2'h1 ? valid_1_115 : _GEN_9230; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10644 = unuse_way == 2'h1 ? valid_1_116 : _GEN_9231; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10645 = unuse_way == 2'h1 ? valid_1_117 : _GEN_9232; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10646 = unuse_way == 2'h1 ? valid_1_118 : _GEN_9233; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10647 = unuse_way == 2'h1 ? valid_1_119 : _GEN_9234; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10648 = unuse_way == 2'h1 ? valid_1_120 : _GEN_9235; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10649 = unuse_way == 2'h1 ? valid_1_121 : _GEN_9236; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10650 = unuse_way == 2'h1 ? valid_1_122 : _GEN_9237; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10651 = unuse_way == 2'h1 ? valid_1_123 : _GEN_9238; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10652 = unuse_way == 2'h1 ? valid_1_124 : _GEN_9239; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10653 = unuse_way == 2'h1 ? valid_1_125 : _GEN_9240; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10654 = unuse_way == 2'h1 ? valid_1_126 : _GEN_9241; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_10655 = unuse_way == 2'h1 ? valid_1_127 : _GEN_9242; // @[d_cache.scala 150:34 31:26]
  wire [63:0] _GEN_10656 = unuse_way == 2'h1 ? write_back_data : _GEN_9244; // @[d_cache.scala 150:34 37:34]
  wire [41:0] _GEN_10657 = unuse_way == 2'h1 ? {{10'd0}, write_back_addr} : _GEN_9245; // @[d_cache.scala 150:34 38:34]
  wire  _GEN_10658 = unuse_way == 2'h1 ? dirty_0_0 : _GEN_9502; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10659 = unuse_way == 2'h1 ? dirty_0_1 : _GEN_9503; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10660 = unuse_way == 2'h1 ? dirty_0_2 : _GEN_9504; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10661 = unuse_way == 2'h1 ? dirty_0_3 : _GEN_9505; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10662 = unuse_way == 2'h1 ? dirty_0_4 : _GEN_9506; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10663 = unuse_way == 2'h1 ? dirty_0_5 : _GEN_9507; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10664 = unuse_way == 2'h1 ? dirty_0_6 : _GEN_9508; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10665 = unuse_way == 2'h1 ? dirty_0_7 : _GEN_9509; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10666 = unuse_way == 2'h1 ? dirty_0_8 : _GEN_9510; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10667 = unuse_way == 2'h1 ? dirty_0_9 : _GEN_9511; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10668 = unuse_way == 2'h1 ? dirty_0_10 : _GEN_9512; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10669 = unuse_way == 2'h1 ? dirty_0_11 : _GEN_9513; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10670 = unuse_way == 2'h1 ? dirty_0_12 : _GEN_9514; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10671 = unuse_way == 2'h1 ? dirty_0_13 : _GEN_9515; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10672 = unuse_way == 2'h1 ? dirty_0_14 : _GEN_9516; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10673 = unuse_way == 2'h1 ? dirty_0_15 : _GEN_9517; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10674 = unuse_way == 2'h1 ? dirty_0_16 : _GEN_9518; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10675 = unuse_way == 2'h1 ? dirty_0_17 : _GEN_9519; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10676 = unuse_way == 2'h1 ? dirty_0_18 : _GEN_9520; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10677 = unuse_way == 2'h1 ? dirty_0_19 : _GEN_9521; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10678 = unuse_way == 2'h1 ? dirty_0_20 : _GEN_9522; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10679 = unuse_way == 2'h1 ? dirty_0_21 : _GEN_9523; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10680 = unuse_way == 2'h1 ? dirty_0_22 : _GEN_9524; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10681 = unuse_way == 2'h1 ? dirty_0_23 : _GEN_9525; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10682 = unuse_way == 2'h1 ? dirty_0_24 : _GEN_9526; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10683 = unuse_way == 2'h1 ? dirty_0_25 : _GEN_9527; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10684 = unuse_way == 2'h1 ? dirty_0_26 : _GEN_9528; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10685 = unuse_way == 2'h1 ? dirty_0_27 : _GEN_9529; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10686 = unuse_way == 2'h1 ? dirty_0_28 : _GEN_9530; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10687 = unuse_way == 2'h1 ? dirty_0_29 : _GEN_9531; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10688 = unuse_way == 2'h1 ? dirty_0_30 : _GEN_9532; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10689 = unuse_way == 2'h1 ? dirty_0_31 : _GEN_9533; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10690 = unuse_way == 2'h1 ? dirty_0_32 : _GEN_9534; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10691 = unuse_way == 2'h1 ? dirty_0_33 : _GEN_9535; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10692 = unuse_way == 2'h1 ? dirty_0_34 : _GEN_9536; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10693 = unuse_way == 2'h1 ? dirty_0_35 : _GEN_9537; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10694 = unuse_way == 2'h1 ? dirty_0_36 : _GEN_9538; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10695 = unuse_way == 2'h1 ? dirty_0_37 : _GEN_9539; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10696 = unuse_way == 2'h1 ? dirty_0_38 : _GEN_9540; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10697 = unuse_way == 2'h1 ? dirty_0_39 : _GEN_9541; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10698 = unuse_way == 2'h1 ? dirty_0_40 : _GEN_9542; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10699 = unuse_way == 2'h1 ? dirty_0_41 : _GEN_9543; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10700 = unuse_way == 2'h1 ? dirty_0_42 : _GEN_9544; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10701 = unuse_way == 2'h1 ? dirty_0_43 : _GEN_9545; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10702 = unuse_way == 2'h1 ? dirty_0_44 : _GEN_9546; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10703 = unuse_way == 2'h1 ? dirty_0_45 : _GEN_9547; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10704 = unuse_way == 2'h1 ? dirty_0_46 : _GEN_9548; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10705 = unuse_way == 2'h1 ? dirty_0_47 : _GEN_9549; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10706 = unuse_way == 2'h1 ? dirty_0_48 : _GEN_9550; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10707 = unuse_way == 2'h1 ? dirty_0_49 : _GEN_9551; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10708 = unuse_way == 2'h1 ? dirty_0_50 : _GEN_9552; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10709 = unuse_way == 2'h1 ? dirty_0_51 : _GEN_9553; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10710 = unuse_way == 2'h1 ? dirty_0_52 : _GEN_9554; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10711 = unuse_way == 2'h1 ? dirty_0_53 : _GEN_9555; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10712 = unuse_way == 2'h1 ? dirty_0_54 : _GEN_9556; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10713 = unuse_way == 2'h1 ? dirty_0_55 : _GEN_9557; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10714 = unuse_way == 2'h1 ? dirty_0_56 : _GEN_9558; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10715 = unuse_way == 2'h1 ? dirty_0_57 : _GEN_9559; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10716 = unuse_way == 2'h1 ? dirty_0_58 : _GEN_9560; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10717 = unuse_way == 2'h1 ? dirty_0_59 : _GEN_9561; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10718 = unuse_way == 2'h1 ? dirty_0_60 : _GEN_9562; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10719 = unuse_way == 2'h1 ? dirty_0_61 : _GEN_9563; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10720 = unuse_way == 2'h1 ? dirty_0_62 : _GEN_9564; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10721 = unuse_way == 2'h1 ? dirty_0_63 : _GEN_9565; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10722 = unuse_way == 2'h1 ? dirty_0_64 : _GEN_9566; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10723 = unuse_way == 2'h1 ? dirty_0_65 : _GEN_9567; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10724 = unuse_way == 2'h1 ? dirty_0_66 : _GEN_9568; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10725 = unuse_way == 2'h1 ? dirty_0_67 : _GEN_9569; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10726 = unuse_way == 2'h1 ? dirty_0_68 : _GEN_9570; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10727 = unuse_way == 2'h1 ? dirty_0_69 : _GEN_9571; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10728 = unuse_way == 2'h1 ? dirty_0_70 : _GEN_9572; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10729 = unuse_way == 2'h1 ? dirty_0_71 : _GEN_9573; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10730 = unuse_way == 2'h1 ? dirty_0_72 : _GEN_9574; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10731 = unuse_way == 2'h1 ? dirty_0_73 : _GEN_9575; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10732 = unuse_way == 2'h1 ? dirty_0_74 : _GEN_9576; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10733 = unuse_way == 2'h1 ? dirty_0_75 : _GEN_9577; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10734 = unuse_way == 2'h1 ? dirty_0_76 : _GEN_9578; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10735 = unuse_way == 2'h1 ? dirty_0_77 : _GEN_9579; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10736 = unuse_way == 2'h1 ? dirty_0_78 : _GEN_9580; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10737 = unuse_way == 2'h1 ? dirty_0_79 : _GEN_9581; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10738 = unuse_way == 2'h1 ? dirty_0_80 : _GEN_9582; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10739 = unuse_way == 2'h1 ? dirty_0_81 : _GEN_9583; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10740 = unuse_way == 2'h1 ? dirty_0_82 : _GEN_9584; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10741 = unuse_way == 2'h1 ? dirty_0_83 : _GEN_9585; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10742 = unuse_way == 2'h1 ? dirty_0_84 : _GEN_9586; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10743 = unuse_way == 2'h1 ? dirty_0_85 : _GEN_9587; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10744 = unuse_way == 2'h1 ? dirty_0_86 : _GEN_9588; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10745 = unuse_way == 2'h1 ? dirty_0_87 : _GEN_9589; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10746 = unuse_way == 2'h1 ? dirty_0_88 : _GEN_9590; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10747 = unuse_way == 2'h1 ? dirty_0_89 : _GEN_9591; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10748 = unuse_way == 2'h1 ? dirty_0_90 : _GEN_9592; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10749 = unuse_way == 2'h1 ? dirty_0_91 : _GEN_9593; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10750 = unuse_way == 2'h1 ? dirty_0_92 : _GEN_9594; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10751 = unuse_way == 2'h1 ? dirty_0_93 : _GEN_9595; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10752 = unuse_way == 2'h1 ? dirty_0_94 : _GEN_9596; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10753 = unuse_way == 2'h1 ? dirty_0_95 : _GEN_9597; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10754 = unuse_way == 2'h1 ? dirty_0_96 : _GEN_9598; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10755 = unuse_way == 2'h1 ? dirty_0_97 : _GEN_9599; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10756 = unuse_way == 2'h1 ? dirty_0_98 : _GEN_9600; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10757 = unuse_way == 2'h1 ? dirty_0_99 : _GEN_9601; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10758 = unuse_way == 2'h1 ? dirty_0_100 : _GEN_9602; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10759 = unuse_way == 2'h1 ? dirty_0_101 : _GEN_9603; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10760 = unuse_way == 2'h1 ? dirty_0_102 : _GEN_9604; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10761 = unuse_way == 2'h1 ? dirty_0_103 : _GEN_9605; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10762 = unuse_way == 2'h1 ? dirty_0_104 : _GEN_9606; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10763 = unuse_way == 2'h1 ? dirty_0_105 : _GEN_9607; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10764 = unuse_way == 2'h1 ? dirty_0_106 : _GEN_9608; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10765 = unuse_way == 2'h1 ? dirty_0_107 : _GEN_9609; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10766 = unuse_way == 2'h1 ? dirty_0_108 : _GEN_9610; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10767 = unuse_way == 2'h1 ? dirty_0_109 : _GEN_9611; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10768 = unuse_way == 2'h1 ? dirty_0_110 : _GEN_9612; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10769 = unuse_way == 2'h1 ? dirty_0_111 : _GEN_9613; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10770 = unuse_way == 2'h1 ? dirty_0_112 : _GEN_9614; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10771 = unuse_way == 2'h1 ? dirty_0_113 : _GEN_9615; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10772 = unuse_way == 2'h1 ? dirty_0_114 : _GEN_9616; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10773 = unuse_way == 2'h1 ? dirty_0_115 : _GEN_9617; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10774 = unuse_way == 2'h1 ? dirty_0_116 : _GEN_9618; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10775 = unuse_way == 2'h1 ? dirty_0_117 : _GEN_9619; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10776 = unuse_way == 2'h1 ? dirty_0_118 : _GEN_9620; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10777 = unuse_way == 2'h1 ? dirty_0_119 : _GEN_9621; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10778 = unuse_way == 2'h1 ? dirty_0_120 : _GEN_9622; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10779 = unuse_way == 2'h1 ? dirty_0_121 : _GEN_9623; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10780 = unuse_way == 2'h1 ? dirty_0_122 : _GEN_9624; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10781 = unuse_way == 2'h1 ? dirty_0_123 : _GEN_9625; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10782 = unuse_way == 2'h1 ? dirty_0_124 : _GEN_9626; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10783 = unuse_way == 2'h1 ? dirty_0_125 : _GEN_9627; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10784 = unuse_way == 2'h1 ? dirty_0_126 : _GEN_9628; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10785 = unuse_way == 2'h1 ? dirty_0_127 : _GEN_9629; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_10786 = unuse_way == 2'h1 ? dirty_1_0 : _GEN_9758; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10787 = unuse_way == 2'h1 ? dirty_1_1 : _GEN_9759; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10788 = unuse_way == 2'h1 ? dirty_1_2 : _GEN_9760; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10789 = unuse_way == 2'h1 ? dirty_1_3 : _GEN_9761; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10790 = unuse_way == 2'h1 ? dirty_1_4 : _GEN_9762; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10791 = unuse_way == 2'h1 ? dirty_1_5 : _GEN_9763; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10792 = unuse_way == 2'h1 ? dirty_1_6 : _GEN_9764; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10793 = unuse_way == 2'h1 ? dirty_1_7 : _GEN_9765; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10794 = unuse_way == 2'h1 ? dirty_1_8 : _GEN_9766; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10795 = unuse_way == 2'h1 ? dirty_1_9 : _GEN_9767; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10796 = unuse_way == 2'h1 ? dirty_1_10 : _GEN_9768; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10797 = unuse_way == 2'h1 ? dirty_1_11 : _GEN_9769; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10798 = unuse_way == 2'h1 ? dirty_1_12 : _GEN_9770; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10799 = unuse_way == 2'h1 ? dirty_1_13 : _GEN_9771; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10800 = unuse_way == 2'h1 ? dirty_1_14 : _GEN_9772; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10801 = unuse_way == 2'h1 ? dirty_1_15 : _GEN_9773; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10802 = unuse_way == 2'h1 ? dirty_1_16 : _GEN_9774; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10803 = unuse_way == 2'h1 ? dirty_1_17 : _GEN_9775; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10804 = unuse_way == 2'h1 ? dirty_1_18 : _GEN_9776; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10805 = unuse_way == 2'h1 ? dirty_1_19 : _GEN_9777; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10806 = unuse_way == 2'h1 ? dirty_1_20 : _GEN_9778; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10807 = unuse_way == 2'h1 ? dirty_1_21 : _GEN_9779; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10808 = unuse_way == 2'h1 ? dirty_1_22 : _GEN_9780; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10809 = unuse_way == 2'h1 ? dirty_1_23 : _GEN_9781; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10810 = unuse_way == 2'h1 ? dirty_1_24 : _GEN_9782; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10811 = unuse_way == 2'h1 ? dirty_1_25 : _GEN_9783; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10812 = unuse_way == 2'h1 ? dirty_1_26 : _GEN_9784; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10813 = unuse_way == 2'h1 ? dirty_1_27 : _GEN_9785; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10814 = unuse_way == 2'h1 ? dirty_1_28 : _GEN_9786; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10815 = unuse_way == 2'h1 ? dirty_1_29 : _GEN_9787; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10816 = unuse_way == 2'h1 ? dirty_1_30 : _GEN_9788; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10817 = unuse_way == 2'h1 ? dirty_1_31 : _GEN_9789; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10818 = unuse_way == 2'h1 ? dirty_1_32 : _GEN_9790; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10819 = unuse_way == 2'h1 ? dirty_1_33 : _GEN_9791; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10820 = unuse_way == 2'h1 ? dirty_1_34 : _GEN_9792; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10821 = unuse_way == 2'h1 ? dirty_1_35 : _GEN_9793; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10822 = unuse_way == 2'h1 ? dirty_1_36 : _GEN_9794; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10823 = unuse_way == 2'h1 ? dirty_1_37 : _GEN_9795; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10824 = unuse_way == 2'h1 ? dirty_1_38 : _GEN_9796; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10825 = unuse_way == 2'h1 ? dirty_1_39 : _GEN_9797; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10826 = unuse_way == 2'h1 ? dirty_1_40 : _GEN_9798; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10827 = unuse_way == 2'h1 ? dirty_1_41 : _GEN_9799; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10828 = unuse_way == 2'h1 ? dirty_1_42 : _GEN_9800; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10829 = unuse_way == 2'h1 ? dirty_1_43 : _GEN_9801; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10830 = unuse_way == 2'h1 ? dirty_1_44 : _GEN_9802; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10831 = unuse_way == 2'h1 ? dirty_1_45 : _GEN_9803; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10832 = unuse_way == 2'h1 ? dirty_1_46 : _GEN_9804; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10833 = unuse_way == 2'h1 ? dirty_1_47 : _GEN_9805; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10834 = unuse_way == 2'h1 ? dirty_1_48 : _GEN_9806; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10835 = unuse_way == 2'h1 ? dirty_1_49 : _GEN_9807; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10836 = unuse_way == 2'h1 ? dirty_1_50 : _GEN_9808; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10837 = unuse_way == 2'h1 ? dirty_1_51 : _GEN_9809; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10838 = unuse_way == 2'h1 ? dirty_1_52 : _GEN_9810; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10839 = unuse_way == 2'h1 ? dirty_1_53 : _GEN_9811; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10840 = unuse_way == 2'h1 ? dirty_1_54 : _GEN_9812; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10841 = unuse_way == 2'h1 ? dirty_1_55 : _GEN_9813; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10842 = unuse_way == 2'h1 ? dirty_1_56 : _GEN_9814; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10843 = unuse_way == 2'h1 ? dirty_1_57 : _GEN_9815; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10844 = unuse_way == 2'h1 ? dirty_1_58 : _GEN_9816; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10845 = unuse_way == 2'h1 ? dirty_1_59 : _GEN_9817; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10846 = unuse_way == 2'h1 ? dirty_1_60 : _GEN_9818; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10847 = unuse_way == 2'h1 ? dirty_1_61 : _GEN_9819; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10848 = unuse_way == 2'h1 ? dirty_1_62 : _GEN_9820; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10849 = unuse_way == 2'h1 ? dirty_1_63 : _GEN_9821; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10850 = unuse_way == 2'h1 ? dirty_1_64 : _GEN_9822; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10851 = unuse_way == 2'h1 ? dirty_1_65 : _GEN_9823; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10852 = unuse_way == 2'h1 ? dirty_1_66 : _GEN_9824; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10853 = unuse_way == 2'h1 ? dirty_1_67 : _GEN_9825; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10854 = unuse_way == 2'h1 ? dirty_1_68 : _GEN_9826; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10855 = unuse_way == 2'h1 ? dirty_1_69 : _GEN_9827; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10856 = unuse_way == 2'h1 ? dirty_1_70 : _GEN_9828; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10857 = unuse_way == 2'h1 ? dirty_1_71 : _GEN_9829; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10858 = unuse_way == 2'h1 ? dirty_1_72 : _GEN_9830; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10859 = unuse_way == 2'h1 ? dirty_1_73 : _GEN_9831; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10860 = unuse_way == 2'h1 ? dirty_1_74 : _GEN_9832; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10861 = unuse_way == 2'h1 ? dirty_1_75 : _GEN_9833; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10862 = unuse_way == 2'h1 ? dirty_1_76 : _GEN_9834; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10863 = unuse_way == 2'h1 ? dirty_1_77 : _GEN_9835; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10864 = unuse_way == 2'h1 ? dirty_1_78 : _GEN_9836; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10865 = unuse_way == 2'h1 ? dirty_1_79 : _GEN_9837; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10866 = unuse_way == 2'h1 ? dirty_1_80 : _GEN_9838; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10867 = unuse_way == 2'h1 ? dirty_1_81 : _GEN_9839; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10868 = unuse_way == 2'h1 ? dirty_1_82 : _GEN_9840; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10869 = unuse_way == 2'h1 ? dirty_1_83 : _GEN_9841; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10870 = unuse_way == 2'h1 ? dirty_1_84 : _GEN_9842; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10871 = unuse_way == 2'h1 ? dirty_1_85 : _GEN_9843; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10872 = unuse_way == 2'h1 ? dirty_1_86 : _GEN_9844; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10873 = unuse_way == 2'h1 ? dirty_1_87 : _GEN_9845; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10874 = unuse_way == 2'h1 ? dirty_1_88 : _GEN_9846; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10875 = unuse_way == 2'h1 ? dirty_1_89 : _GEN_9847; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10876 = unuse_way == 2'h1 ? dirty_1_90 : _GEN_9848; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10877 = unuse_way == 2'h1 ? dirty_1_91 : _GEN_9849; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10878 = unuse_way == 2'h1 ? dirty_1_92 : _GEN_9850; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10879 = unuse_way == 2'h1 ? dirty_1_93 : _GEN_9851; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10880 = unuse_way == 2'h1 ? dirty_1_94 : _GEN_9852; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10881 = unuse_way == 2'h1 ? dirty_1_95 : _GEN_9853; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10882 = unuse_way == 2'h1 ? dirty_1_96 : _GEN_9854; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10883 = unuse_way == 2'h1 ? dirty_1_97 : _GEN_9855; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10884 = unuse_way == 2'h1 ? dirty_1_98 : _GEN_9856; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10885 = unuse_way == 2'h1 ? dirty_1_99 : _GEN_9857; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10886 = unuse_way == 2'h1 ? dirty_1_100 : _GEN_9858; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10887 = unuse_way == 2'h1 ? dirty_1_101 : _GEN_9859; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10888 = unuse_way == 2'h1 ? dirty_1_102 : _GEN_9860; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10889 = unuse_way == 2'h1 ? dirty_1_103 : _GEN_9861; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10890 = unuse_way == 2'h1 ? dirty_1_104 : _GEN_9862; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10891 = unuse_way == 2'h1 ? dirty_1_105 : _GEN_9863; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10892 = unuse_way == 2'h1 ? dirty_1_106 : _GEN_9864; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10893 = unuse_way == 2'h1 ? dirty_1_107 : _GEN_9865; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10894 = unuse_way == 2'h1 ? dirty_1_108 : _GEN_9866; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10895 = unuse_way == 2'h1 ? dirty_1_109 : _GEN_9867; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10896 = unuse_way == 2'h1 ? dirty_1_110 : _GEN_9868; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10897 = unuse_way == 2'h1 ? dirty_1_111 : _GEN_9869; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10898 = unuse_way == 2'h1 ? dirty_1_112 : _GEN_9870; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10899 = unuse_way == 2'h1 ? dirty_1_113 : _GEN_9871; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10900 = unuse_way == 2'h1 ? dirty_1_114 : _GEN_9872; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10901 = unuse_way == 2'h1 ? dirty_1_115 : _GEN_9873; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10902 = unuse_way == 2'h1 ? dirty_1_116 : _GEN_9874; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10903 = unuse_way == 2'h1 ? dirty_1_117 : _GEN_9875; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10904 = unuse_way == 2'h1 ? dirty_1_118 : _GEN_9876; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10905 = unuse_way == 2'h1 ? dirty_1_119 : _GEN_9877; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10906 = unuse_way == 2'h1 ? dirty_1_120 : _GEN_9878; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10907 = unuse_way == 2'h1 ? dirty_1_121 : _GEN_9879; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10908 = unuse_way == 2'h1 ? dirty_1_122 : _GEN_9880; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10909 = unuse_way == 2'h1 ? dirty_1_123 : _GEN_9881; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10910 = unuse_way == 2'h1 ? dirty_1_124 : _GEN_9882; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10911 = unuse_way == 2'h1 ? dirty_1_125 : _GEN_9883; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10912 = unuse_way == 2'h1 ? dirty_1_126 : _GEN_9884; // @[d_cache.scala 150:34 33:26]
  wire  _GEN_10913 = unuse_way == 2'h1 ? dirty_1_127 : _GEN_9885; // @[d_cache.scala 150:34 33:26]
  wire [2:0] _GEN_10914 = io_from_axi_bvalid ? 3'h7 : state; // @[d_cache.scala 202:37 203:23 82:24]
  wire [2:0] _GEN_10915 = 3'h7 == state ? 3'h1 : state; // @[d_cache.scala 87:18 207:19 82:24]
  wire [2:0] _GEN_10916 = 3'h6 == state ? _GEN_10914 : _GEN_10915; // @[d_cache.scala 87:18]
  wire [2:0] _GEN_10917 = 3'h5 == state ? _GEN_9886 : _GEN_10916; // @[d_cache.scala 87:18]
  wire [63:0] _GEN_10918 = 3'h5 == state ? _GEN_9887 : ram_0_0; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10919 = 3'h5 == state ? _GEN_9888 : ram_0_1; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10920 = 3'h5 == state ? _GEN_9889 : ram_0_2; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10921 = 3'h5 == state ? _GEN_9890 : ram_0_3; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10922 = 3'h5 == state ? _GEN_9891 : ram_0_4; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10923 = 3'h5 == state ? _GEN_9892 : ram_0_5; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10924 = 3'h5 == state ? _GEN_9893 : ram_0_6; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10925 = 3'h5 == state ? _GEN_9894 : ram_0_7; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10926 = 3'h5 == state ? _GEN_9895 : ram_0_8; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10927 = 3'h5 == state ? _GEN_9896 : ram_0_9; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10928 = 3'h5 == state ? _GEN_9897 : ram_0_10; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10929 = 3'h5 == state ? _GEN_9898 : ram_0_11; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10930 = 3'h5 == state ? _GEN_9899 : ram_0_12; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10931 = 3'h5 == state ? _GEN_9900 : ram_0_13; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10932 = 3'h5 == state ? _GEN_9901 : ram_0_14; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10933 = 3'h5 == state ? _GEN_9902 : ram_0_15; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10934 = 3'h5 == state ? _GEN_9903 : ram_0_16; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10935 = 3'h5 == state ? _GEN_9904 : ram_0_17; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10936 = 3'h5 == state ? _GEN_9905 : ram_0_18; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10937 = 3'h5 == state ? _GEN_9906 : ram_0_19; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10938 = 3'h5 == state ? _GEN_9907 : ram_0_20; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10939 = 3'h5 == state ? _GEN_9908 : ram_0_21; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10940 = 3'h5 == state ? _GEN_9909 : ram_0_22; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10941 = 3'h5 == state ? _GEN_9910 : ram_0_23; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10942 = 3'h5 == state ? _GEN_9911 : ram_0_24; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10943 = 3'h5 == state ? _GEN_9912 : ram_0_25; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10944 = 3'h5 == state ? _GEN_9913 : ram_0_26; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10945 = 3'h5 == state ? _GEN_9914 : ram_0_27; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10946 = 3'h5 == state ? _GEN_9915 : ram_0_28; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10947 = 3'h5 == state ? _GEN_9916 : ram_0_29; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10948 = 3'h5 == state ? _GEN_9917 : ram_0_30; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10949 = 3'h5 == state ? _GEN_9918 : ram_0_31; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10950 = 3'h5 == state ? _GEN_9919 : ram_0_32; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10951 = 3'h5 == state ? _GEN_9920 : ram_0_33; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10952 = 3'h5 == state ? _GEN_9921 : ram_0_34; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10953 = 3'h5 == state ? _GEN_9922 : ram_0_35; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10954 = 3'h5 == state ? _GEN_9923 : ram_0_36; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10955 = 3'h5 == state ? _GEN_9924 : ram_0_37; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10956 = 3'h5 == state ? _GEN_9925 : ram_0_38; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10957 = 3'h5 == state ? _GEN_9926 : ram_0_39; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10958 = 3'h5 == state ? _GEN_9927 : ram_0_40; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10959 = 3'h5 == state ? _GEN_9928 : ram_0_41; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10960 = 3'h5 == state ? _GEN_9929 : ram_0_42; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10961 = 3'h5 == state ? _GEN_9930 : ram_0_43; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10962 = 3'h5 == state ? _GEN_9931 : ram_0_44; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10963 = 3'h5 == state ? _GEN_9932 : ram_0_45; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10964 = 3'h5 == state ? _GEN_9933 : ram_0_46; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10965 = 3'h5 == state ? _GEN_9934 : ram_0_47; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10966 = 3'h5 == state ? _GEN_9935 : ram_0_48; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10967 = 3'h5 == state ? _GEN_9936 : ram_0_49; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10968 = 3'h5 == state ? _GEN_9937 : ram_0_50; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10969 = 3'h5 == state ? _GEN_9938 : ram_0_51; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10970 = 3'h5 == state ? _GEN_9939 : ram_0_52; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10971 = 3'h5 == state ? _GEN_9940 : ram_0_53; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10972 = 3'h5 == state ? _GEN_9941 : ram_0_54; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10973 = 3'h5 == state ? _GEN_9942 : ram_0_55; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10974 = 3'h5 == state ? _GEN_9943 : ram_0_56; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10975 = 3'h5 == state ? _GEN_9944 : ram_0_57; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10976 = 3'h5 == state ? _GEN_9945 : ram_0_58; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10977 = 3'h5 == state ? _GEN_9946 : ram_0_59; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10978 = 3'h5 == state ? _GEN_9947 : ram_0_60; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10979 = 3'h5 == state ? _GEN_9948 : ram_0_61; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10980 = 3'h5 == state ? _GEN_9949 : ram_0_62; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10981 = 3'h5 == state ? _GEN_9950 : ram_0_63; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10982 = 3'h5 == state ? _GEN_9951 : ram_0_64; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10983 = 3'h5 == state ? _GEN_9952 : ram_0_65; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10984 = 3'h5 == state ? _GEN_9953 : ram_0_66; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10985 = 3'h5 == state ? _GEN_9954 : ram_0_67; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10986 = 3'h5 == state ? _GEN_9955 : ram_0_68; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10987 = 3'h5 == state ? _GEN_9956 : ram_0_69; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10988 = 3'h5 == state ? _GEN_9957 : ram_0_70; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10989 = 3'h5 == state ? _GEN_9958 : ram_0_71; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10990 = 3'h5 == state ? _GEN_9959 : ram_0_72; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10991 = 3'h5 == state ? _GEN_9960 : ram_0_73; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10992 = 3'h5 == state ? _GEN_9961 : ram_0_74; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10993 = 3'h5 == state ? _GEN_9962 : ram_0_75; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10994 = 3'h5 == state ? _GEN_9963 : ram_0_76; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10995 = 3'h5 == state ? _GEN_9964 : ram_0_77; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10996 = 3'h5 == state ? _GEN_9965 : ram_0_78; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10997 = 3'h5 == state ? _GEN_9966 : ram_0_79; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10998 = 3'h5 == state ? _GEN_9967 : ram_0_80; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_10999 = 3'h5 == state ? _GEN_9968 : ram_0_81; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11000 = 3'h5 == state ? _GEN_9969 : ram_0_82; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11001 = 3'h5 == state ? _GEN_9970 : ram_0_83; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11002 = 3'h5 == state ? _GEN_9971 : ram_0_84; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11003 = 3'h5 == state ? _GEN_9972 : ram_0_85; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11004 = 3'h5 == state ? _GEN_9973 : ram_0_86; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11005 = 3'h5 == state ? _GEN_9974 : ram_0_87; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11006 = 3'h5 == state ? _GEN_9975 : ram_0_88; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11007 = 3'h5 == state ? _GEN_9976 : ram_0_89; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11008 = 3'h5 == state ? _GEN_9977 : ram_0_90; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11009 = 3'h5 == state ? _GEN_9978 : ram_0_91; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11010 = 3'h5 == state ? _GEN_9979 : ram_0_92; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11011 = 3'h5 == state ? _GEN_9980 : ram_0_93; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11012 = 3'h5 == state ? _GEN_9981 : ram_0_94; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11013 = 3'h5 == state ? _GEN_9982 : ram_0_95; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11014 = 3'h5 == state ? _GEN_9983 : ram_0_96; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11015 = 3'h5 == state ? _GEN_9984 : ram_0_97; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11016 = 3'h5 == state ? _GEN_9985 : ram_0_98; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11017 = 3'h5 == state ? _GEN_9986 : ram_0_99; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11018 = 3'h5 == state ? _GEN_9987 : ram_0_100; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11019 = 3'h5 == state ? _GEN_9988 : ram_0_101; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11020 = 3'h5 == state ? _GEN_9989 : ram_0_102; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11021 = 3'h5 == state ? _GEN_9990 : ram_0_103; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11022 = 3'h5 == state ? _GEN_9991 : ram_0_104; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11023 = 3'h5 == state ? _GEN_9992 : ram_0_105; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11024 = 3'h5 == state ? _GEN_9993 : ram_0_106; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11025 = 3'h5 == state ? _GEN_9994 : ram_0_107; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11026 = 3'h5 == state ? _GEN_9995 : ram_0_108; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11027 = 3'h5 == state ? _GEN_9996 : ram_0_109; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11028 = 3'h5 == state ? _GEN_9997 : ram_0_110; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11029 = 3'h5 == state ? _GEN_9998 : ram_0_111; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11030 = 3'h5 == state ? _GEN_9999 : ram_0_112; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11031 = 3'h5 == state ? _GEN_10000 : ram_0_113; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11032 = 3'h5 == state ? _GEN_10001 : ram_0_114; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11033 = 3'h5 == state ? _GEN_10002 : ram_0_115; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11034 = 3'h5 == state ? _GEN_10003 : ram_0_116; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11035 = 3'h5 == state ? _GEN_10004 : ram_0_117; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11036 = 3'h5 == state ? _GEN_10005 : ram_0_118; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11037 = 3'h5 == state ? _GEN_10006 : ram_0_119; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11038 = 3'h5 == state ? _GEN_10007 : ram_0_120; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11039 = 3'h5 == state ? _GEN_10008 : ram_0_121; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11040 = 3'h5 == state ? _GEN_10009 : ram_0_122; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11041 = 3'h5 == state ? _GEN_10010 : ram_0_123; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11042 = 3'h5 == state ? _GEN_10011 : ram_0_124; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11043 = 3'h5 == state ? _GEN_10012 : ram_0_125; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11044 = 3'h5 == state ? _GEN_10013 : ram_0_126; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11045 = 3'h5 == state ? _GEN_10014 : ram_0_127; // @[d_cache.scala 87:18 19:24]
  wire [31:0] _GEN_11046 = 3'h5 == state ? _GEN_10015 : tag_0_0; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11047 = 3'h5 == state ? _GEN_10016 : tag_0_1; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11048 = 3'h5 == state ? _GEN_10017 : tag_0_2; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11049 = 3'h5 == state ? _GEN_10018 : tag_0_3; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11050 = 3'h5 == state ? _GEN_10019 : tag_0_4; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11051 = 3'h5 == state ? _GEN_10020 : tag_0_5; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11052 = 3'h5 == state ? _GEN_10021 : tag_0_6; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11053 = 3'h5 == state ? _GEN_10022 : tag_0_7; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11054 = 3'h5 == state ? _GEN_10023 : tag_0_8; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11055 = 3'h5 == state ? _GEN_10024 : tag_0_9; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11056 = 3'h5 == state ? _GEN_10025 : tag_0_10; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11057 = 3'h5 == state ? _GEN_10026 : tag_0_11; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11058 = 3'h5 == state ? _GEN_10027 : tag_0_12; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11059 = 3'h5 == state ? _GEN_10028 : tag_0_13; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11060 = 3'h5 == state ? _GEN_10029 : tag_0_14; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11061 = 3'h5 == state ? _GEN_10030 : tag_0_15; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11062 = 3'h5 == state ? _GEN_10031 : tag_0_16; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11063 = 3'h5 == state ? _GEN_10032 : tag_0_17; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11064 = 3'h5 == state ? _GEN_10033 : tag_0_18; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11065 = 3'h5 == state ? _GEN_10034 : tag_0_19; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11066 = 3'h5 == state ? _GEN_10035 : tag_0_20; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11067 = 3'h5 == state ? _GEN_10036 : tag_0_21; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11068 = 3'h5 == state ? _GEN_10037 : tag_0_22; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11069 = 3'h5 == state ? _GEN_10038 : tag_0_23; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11070 = 3'h5 == state ? _GEN_10039 : tag_0_24; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11071 = 3'h5 == state ? _GEN_10040 : tag_0_25; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11072 = 3'h5 == state ? _GEN_10041 : tag_0_26; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11073 = 3'h5 == state ? _GEN_10042 : tag_0_27; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11074 = 3'h5 == state ? _GEN_10043 : tag_0_28; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11075 = 3'h5 == state ? _GEN_10044 : tag_0_29; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11076 = 3'h5 == state ? _GEN_10045 : tag_0_30; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11077 = 3'h5 == state ? _GEN_10046 : tag_0_31; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11078 = 3'h5 == state ? _GEN_10047 : tag_0_32; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11079 = 3'h5 == state ? _GEN_10048 : tag_0_33; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11080 = 3'h5 == state ? _GEN_10049 : tag_0_34; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11081 = 3'h5 == state ? _GEN_10050 : tag_0_35; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11082 = 3'h5 == state ? _GEN_10051 : tag_0_36; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11083 = 3'h5 == state ? _GEN_10052 : tag_0_37; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11084 = 3'h5 == state ? _GEN_10053 : tag_0_38; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11085 = 3'h5 == state ? _GEN_10054 : tag_0_39; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11086 = 3'h5 == state ? _GEN_10055 : tag_0_40; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11087 = 3'h5 == state ? _GEN_10056 : tag_0_41; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11088 = 3'h5 == state ? _GEN_10057 : tag_0_42; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11089 = 3'h5 == state ? _GEN_10058 : tag_0_43; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11090 = 3'h5 == state ? _GEN_10059 : tag_0_44; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11091 = 3'h5 == state ? _GEN_10060 : tag_0_45; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11092 = 3'h5 == state ? _GEN_10061 : tag_0_46; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11093 = 3'h5 == state ? _GEN_10062 : tag_0_47; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11094 = 3'h5 == state ? _GEN_10063 : tag_0_48; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11095 = 3'h5 == state ? _GEN_10064 : tag_0_49; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11096 = 3'h5 == state ? _GEN_10065 : tag_0_50; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11097 = 3'h5 == state ? _GEN_10066 : tag_0_51; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11098 = 3'h5 == state ? _GEN_10067 : tag_0_52; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11099 = 3'h5 == state ? _GEN_10068 : tag_0_53; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11100 = 3'h5 == state ? _GEN_10069 : tag_0_54; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11101 = 3'h5 == state ? _GEN_10070 : tag_0_55; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11102 = 3'h5 == state ? _GEN_10071 : tag_0_56; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11103 = 3'h5 == state ? _GEN_10072 : tag_0_57; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11104 = 3'h5 == state ? _GEN_10073 : tag_0_58; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11105 = 3'h5 == state ? _GEN_10074 : tag_0_59; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11106 = 3'h5 == state ? _GEN_10075 : tag_0_60; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11107 = 3'h5 == state ? _GEN_10076 : tag_0_61; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11108 = 3'h5 == state ? _GEN_10077 : tag_0_62; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11109 = 3'h5 == state ? _GEN_10078 : tag_0_63; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11110 = 3'h5 == state ? _GEN_10079 : tag_0_64; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11111 = 3'h5 == state ? _GEN_10080 : tag_0_65; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11112 = 3'h5 == state ? _GEN_10081 : tag_0_66; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11113 = 3'h5 == state ? _GEN_10082 : tag_0_67; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11114 = 3'h5 == state ? _GEN_10083 : tag_0_68; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11115 = 3'h5 == state ? _GEN_10084 : tag_0_69; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11116 = 3'h5 == state ? _GEN_10085 : tag_0_70; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11117 = 3'h5 == state ? _GEN_10086 : tag_0_71; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11118 = 3'h5 == state ? _GEN_10087 : tag_0_72; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11119 = 3'h5 == state ? _GEN_10088 : tag_0_73; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11120 = 3'h5 == state ? _GEN_10089 : tag_0_74; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11121 = 3'h5 == state ? _GEN_10090 : tag_0_75; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11122 = 3'h5 == state ? _GEN_10091 : tag_0_76; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11123 = 3'h5 == state ? _GEN_10092 : tag_0_77; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11124 = 3'h5 == state ? _GEN_10093 : tag_0_78; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11125 = 3'h5 == state ? _GEN_10094 : tag_0_79; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11126 = 3'h5 == state ? _GEN_10095 : tag_0_80; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11127 = 3'h5 == state ? _GEN_10096 : tag_0_81; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11128 = 3'h5 == state ? _GEN_10097 : tag_0_82; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11129 = 3'h5 == state ? _GEN_10098 : tag_0_83; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11130 = 3'h5 == state ? _GEN_10099 : tag_0_84; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11131 = 3'h5 == state ? _GEN_10100 : tag_0_85; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11132 = 3'h5 == state ? _GEN_10101 : tag_0_86; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11133 = 3'h5 == state ? _GEN_10102 : tag_0_87; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11134 = 3'h5 == state ? _GEN_10103 : tag_0_88; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11135 = 3'h5 == state ? _GEN_10104 : tag_0_89; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11136 = 3'h5 == state ? _GEN_10105 : tag_0_90; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11137 = 3'h5 == state ? _GEN_10106 : tag_0_91; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11138 = 3'h5 == state ? _GEN_10107 : tag_0_92; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11139 = 3'h5 == state ? _GEN_10108 : tag_0_93; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11140 = 3'h5 == state ? _GEN_10109 : tag_0_94; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11141 = 3'h5 == state ? _GEN_10110 : tag_0_95; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11142 = 3'h5 == state ? _GEN_10111 : tag_0_96; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11143 = 3'h5 == state ? _GEN_10112 : tag_0_97; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11144 = 3'h5 == state ? _GEN_10113 : tag_0_98; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11145 = 3'h5 == state ? _GEN_10114 : tag_0_99; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11146 = 3'h5 == state ? _GEN_10115 : tag_0_100; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11147 = 3'h5 == state ? _GEN_10116 : tag_0_101; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11148 = 3'h5 == state ? _GEN_10117 : tag_0_102; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11149 = 3'h5 == state ? _GEN_10118 : tag_0_103; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11150 = 3'h5 == state ? _GEN_10119 : tag_0_104; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11151 = 3'h5 == state ? _GEN_10120 : tag_0_105; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11152 = 3'h5 == state ? _GEN_10121 : tag_0_106; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11153 = 3'h5 == state ? _GEN_10122 : tag_0_107; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11154 = 3'h5 == state ? _GEN_10123 : tag_0_108; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11155 = 3'h5 == state ? _GEN_10124 : tag_0_109; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11156 = 3'h5 == state ? _GEN_10125 : tag_0_110; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11157 = 3'h5 == state ? _GEN_10126 : tag_0_111; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11158 = 3'h5 == state ? _GEN_10127 : tag_0_112; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11159 = 3'h5 == state ? _GEN_10128 : tag_0_113; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11160 = 3'h5 == state ? _GEN_10129 : tag_0_114; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11161 = 3'h5 == state ? _GEN_10130 : tag_0_115; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11162 = 3'h5 == state ? _GEN_10131 : tag_0_116; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11163 = 3'h5 == state ? _GEN_10132 : tag_0_117; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11164 = 3'h5 == state ? _GEN_10133 : tag_0_118; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11165 = 3'h5 == state ? _GEN_10134 : tag_0_119; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11166 = 3'h5 == state ? _GEN_10135 : tag_0_120; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11167 = 3'h5 == state ? _GEN_10136 : tag_0_121; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11168 = 3'h5 == state ? _GEN_10137 : tag_0_122; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11169 = 3'h5 == state ? _GEN_10138 : tag_0_123; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11170 = 3'h5 == state ? _GEN_10139 : tag_0_124; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11171 = 3'h5 == state ? _GEN_10140 : tag_0_125; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11172 = 3'h5 == state ? _GEN_10141 : tag_0_126; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_11173 = 3'h5 == state ? _GEN_10142 : tag_0_127; // @[d_cache.scala 87:18 28:24]
  wire  _GEN_11174 = 3'h5 == state ? _GEN_10143 : valid_0_0; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11175 = 3'h5 == state ? _GEN_10144 : valid_0_1; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11176 = 3'h5 == state ? _GEN_10145 : valid_0_2; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11177 = 3'h5 == state ? _GEN_10146 : valid_0_3; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11178 = 3'h5 == state ? _GEN_10147 : valid_0_4; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11179 = 3'h5 == state ? _GEN_10148 : valid_0_5; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11180 = 3'h5 == state ? _GEN_10149 : valid_0_6; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11181 = 3'h5 == state ? _GEN_10150 : valid_0_7; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11182 = 3'h5 == state ? _GEN_10151 : valid_0_8; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11183 = 3'h5 == state ? _GEN_10152 : valid_0_9; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11184 = 3'h5 == state ? _GEN_10153 : valid_0_10; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11185 = 3'h5 == state ? _GEN_10154 : valid_0_11; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11186 = 3'h5 == state ? _GEN_10155 : valid_0_12; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11187 = 3'h5 == state ? _GEN_10156 : valid_0_13; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11188 = 3'h5 == state ? _GEN_10157 : valid_0_14; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11189 = 3'h5 == state ? _GEN_10158 : valid_0_15; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11190 = 3'h5 == state ? _GEN_10159 : valid_0_16; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11191 = 3'h5 == state ? _GEN_10160 : valid_0_17; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11192 = 3'h5 == state ? _GEN_10161 : valid_0_18; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11193 = 3'h5 == state ? _GEN_10162 : valid_0_19; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11194 = 3'h5 == state ? _GEN_10163 : valid_0_20; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11195 = 3'h5 == state ? _GEN_10164 : valid_0_21; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11196 = 3'h5 == state ? _GEN_10165 : valid_0_22; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11197 = 3'h5 == state ? _GEN_10166 : valid_0_23; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11198 = 3'h5 == state ? _GEN_10167 : valid_0_24; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11199 = 3'h5 == state ? _GEN_10168 : valid_0_25; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11200 = 3'h5 == state ? _GEN_10169 : valid_0_26; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11201 = 3'h5 == state ? _GEN_10170 : valid_0_27; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11202 = 3'h5 == state ? _GEN_10171 : valid_0_28; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11203 = 3'h5 == state ? _GEN_10172 : valid_0_29; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11204 = 3'h5 == state ? _GEN_10173 : valid_0_30; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11205 = 3'h5 == state ? _GEN_10174 : valid_0_31; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11206 = 3'h5 == state ? _GEN_10175 : valid_0_32; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11207 = 3'h5 == state ? _GEN_10176 : valid_0_33; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11208 = 3'h5 == state ? _GEN_10177 : valid_0_34; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11209 = 3'h5 == state ? _GEN_10178 : valid_0_35; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11210 = 3'h5 == state ? _GEN_10179 : valid_0_36; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11211 = 3'h5 == state ? _GEN_10180 : valid_0_37; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11212 = 3'h5 == state ? _GEN_10181 : valid_0_38; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11213 = 3'h5 == state ? _GEN_10182 : valid_0_39; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11214 = 3'h5 == state ? _GEN_10183 : valid_0_40; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11215 = 3'h5 == state ? _GEN_10184 : valid_0_41; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11216 = 3'h5 == state ? _GEN_10185 : valid_0_42; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11217 = 3'h5 == state ? _GEN_10186 : valid_0_43; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11218 = 3'h5 == state ? _GEN_10187 : valid_0_44; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11219 = 3'h5 == state ? _GEN_10188 : valid_0_45; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11220 = 3'h5 == state ? _GEN_10189 : valid_0_46; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11221 = 3'h5 == state ? _GEN_10190 : valid_0_47; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11222 = 3'h5 == state ? _GEN_10191 : valid_0_48; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11223 = 3'h5 == state ? _GEN_10192 : valid_0_49; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11224 = 3'h5 == state ? _GEN_10193 : valid_0_50; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11225 = 3'h5 == state ? _GEN_10194 : valid_0_51; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11226 = 3'h5 == state ? _GEN_10195 : valid_0_52; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11227 = 3'h5 == state ? _GEN_10196 : valid_0_53; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11228 = 3'h5 == state ? _GEN_10197 : valid_0_54; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11229 = 3'h5 == state ? _GEN_10198 : valid_0_55; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11230 = 3'h5 == state ? _GEN_10199 : valid_0_56; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11231 = 3'h5 == state ? _GEN_10200 : valid_0_57; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11232 = 3'h5 == state ? _GEN_10201 : valid_0_58; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11233 = 3'h5 == state ? _GEN_10202 : valid_0_59; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11234 = 3'h5 == state ? _GEN_10203 : valid_0_60; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11235 = 3'h5 == state ? _GEN_10204 : valid_0_61; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11236 = 3'h5 == state ? _GEN_10205 : valid_0_62; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11237 = 3'h5 == state ? _GEN_10206 : valid_0_63; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11238 = 3'h5 == state ? _GEN_10207 : valid_0_64; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11239 = 3'h5 == state ? _GEN_10208 : valid_0_65; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11240 = 3'h5 == state ? _GEN_10209 : valid_0_66; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11241 = 3'h5 == state ? _GEN_10210 : valid_0_67; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11242 = 3'h5 == state ? _GEN_10211 : valid_0_68; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11243 = 3'h5 == state ? _GEN_10212 : valid_0_69; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11244 = 3'h5 == state ? _GEN_10213 : valid_0_70; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11245 = 3'h5 == state ? _GEN_10214 : valid_0_71; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11246 = 3'h5 == state ? _GEN_10215 : valid_0_72; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11247 = 3'h5 == state ? _GEN_10216 : valid_0_73; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11248 = 3'h5 == state ? _GEN_10217 : valid_0_74; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11249 = 3'h5 == state ? _GEN_10218 : valid_0_75; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11250 = 3'h5 == state ? _GEN_10219 : valid_0_76; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11251 = 3'h5 == state ? _GEN_10220 : valid_0_77; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11252 = 3'h5 == state ? _GEN_10221 : valid_0_78; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11253 = 3'h5 == state ? _GEN_10222 : valid_0_79; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11254 = 3'h5 == state ? _GEN_10223 : valid_0_80; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11255 = 3'h5 == state ? _GEN_10224 : valid_0_81; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11256 = 3'h5 == state ? _GEN_10225 : valid_0_82; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11257 = 3'h5 == state ? _GEN_10226 : valid_0_83; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11258 = 3'h5 == state ? _GEN_10227 : valid_0_84; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11259 = 3'h5 == state ? _GEN_10228 : valid_0_85; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11260 = 3'h5 == state ? _GEN_10229 : valid_0_86; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11261 = 3'h5 == state ? _GEN_10230 : valid_0_87; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11262 = 3'h5 == state ? _GEN_10231 : valid_0_88; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11263 = 3'h5 == state ? _GEN_10232 : valid_0_89; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11264 = 3'h5 == state ? _GEN_10233 : valid_0_90; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11265 = 3'h5 == state ? _GEN_10234 : valid_0_91; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11266 = 3'h5 == state ? _GEN_10235 : valid_0_92; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11267 = 3'h5 == state ? _GEN_10236 : valid_0_93; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11268 = 3'h5 == state ? _GEN_10237 : valid_0_94; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11269 = 3'h5 == state ? _GEN_10238 : valid_0_95; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11270 = 3'h5 == state ? _GEN_10239 : valid_0_96; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11271 = 3'h5 == state ? _GEN_10240 : valid_0_97; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11272 = 3'h5 == state ? _GEN_10241 : valid_0_98; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11273 = 3'h5 == state ? _GEN_10242 : valid_0_99; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11274 = 3'h5 == state ? _GEN_10243 : valid_0_100; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11275 = 3'h5 == state ? _GEN_10244 : valid_0_101; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11276 = 3'h5 == state ? _GEN_10245 : valid_0_102; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11277 = 3'h5 == state ? _GEN_10246 : valid_0_103; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11278 = 3'h5 == state ? _GEN_10247 : valid_0_104; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11279 = 3'h5 == state ? _GEN_10248 : valid_0_105; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11280 = 3'h5 == state ? _GEN_10249 : valid_0_106; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11281 = 3'h5 == state ? _GEN_10250 : valid_0_107; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11282 = 3'h5 == state ? _GEN_10251 : valid_0_108; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11283 = 3'h5 == state ? _GEN_10252 : valid_0_109; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11284 = 3'h5 == state ? _GEN_10253 : valid_0_110; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11285 = 3'h5 == state ? _GEN_10254 : valid_0_111; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11286 = 3'h5 == state ? _GEN_10255 : valid_0_112; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11287 = 3'h5 == state ? _GEN_10256 : valid_0_113; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11288 = 3'h5 == state ? _GEN_10257 : valid_0_114; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11289 = 3'h5 == state ? _GEN_10258 : valid_0_115; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11290 = 3'h5 == state ? _GEN_10259 : valid_0_116; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11291 = 3'h5 == state ? _GEN_10260 : valid_0_117; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11292 = 3'h5 == state ? _GEN_10261 : valid_0_118; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11293 = 3'h5 == state ? _GEN_10262 : valid_0_119; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11294 = 3'h5 == state ? _GEN_10263 : valid_0_120; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11295 = 3'h5 == state ? _GEN_10264 : valid_0_121; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11296 = 3'h5 == state ? _GEN_10265 : valid_0_122; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11297 = 3'h5 == state ? _GEN_10266 : valid_0_123; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11298 = 3'h5 == state ? _GEN_10267 : valid_0_124; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11299 = 3'h5 == state ? _GEN_10268 : valid_0_125; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11300 = 3'h5 == state ? _GEN_10269 : valid_0_126; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11301 = 3'h5 == state ? _GEN_10270 : valid_0_127; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_11302 = 3'h5 == state ? _GEN_10271 : quene; // @[d_cache.scala 87:18 43:24]
  wire [63:0] _GEN_11303 = 3'h5 == state ? _GEN_10272 : ram_1_0; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11304 = 3'h5 == state ? _GEN_10273 : ram_1_1; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11305 = 3'h5 == state ? _GEN_10274 : ram_1_2; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11306 = 3'h5 == state ? _GEN_10275 : ram_1_3; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11307 = 3'h5 == state ? _GEN_10276 : ram_1_4; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11308 = 3'h5 == state ? _GEN_10277 : ram_1_5; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11309 = 3'h5 == state ? _GEN_10278 : ram_1_6; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11310 = 3'h5 == state ? _GEN_10279 : ram_1_7; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11311 = 3'h5 == state ? _GEN_10280 : ram_1_8; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11312 = 3'h5 == state ? _GEN_10281 : ram_1_9; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11313 = 3'h5 == state ? _GEN_10282 : ram_1_10; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11314 = 3'h5 == state ? _GEN_10283 : ram_1_11; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11315 = 3'h5 == state ? _GEN_10284 : ram_1_12; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11316 = 3'h5 == state ? _GEN_10285 : ram_1_13; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11317 = 3'h5 == state ? _GEN_10286 : ram_1_14; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11318 = 3'h5 == state ? _GEN_10287 : ram_1_15; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11319 = 3'h5 == state ? _GEN_10288 : ram_1_16; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11320 = 3'h5 == state ? _GEN_10289 : ram_1_17; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11321 = 3'h5 == state ? _GEN_10290 : ram_1_18; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11322 = 3'h5 == state ? _GEN_10291 : ram_1_19; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11323 = 3'h5 == state ? _GEN_10292 : ram_1_20; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11324 = 3'h5 == state ? _GEN_10293 : ram_1_21; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11325 = 3'h5 == state ? _GEN_10294 : ram_1_22; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11326 = 3'h5 == state ? _GEN_10295 : ram_1_23; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11327 = 3'h5 == state ? _GEN_10296 : ram_1_24; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11328 = 3'h5 == state ? _GEN_10297 : ram_1_25; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11329 = 3'h5 == state ? _GEN_10298 : ram_1_26; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11330 = 3'h5 == state ? _GEN_10299 : ram_1_27; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11331 = 3'h5 == state ? _GEN_10300 : ram_1_28; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11332 = 3'h5 == state ? _GEN_10301 : ram_1_29; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11333 = 3'h5 == state ? _GEN_10302 : ram_1_30; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11334 = 3'h5 == state ? _GEN_10303 : ram_1_31; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11335 = 3'h5 == state ? _GEN_10304 : ram_1_32; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11336 = 3'h5 == state ? _GEN_10305 : ram_1_33; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11337 = 3'h5 == state ? _GEN_10306 : ram_1_34; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11338 = 3'h5 == state ? _GEN_10307 : ram_1_35; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11339 = 3'h5 == state ? _GEN_10308 : ram_1_36; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11340 = 3'h5 == state ? _GEN_10309 : ram_1_37; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11341 = 3'h5 == state ? _GEN_10310 : ram_1_38; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11342 = 3'h5 == state ? _GEN_10311 : ram_1_39; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11343 = 3'h5 == state ? _GEN_10312 : ram_1_40; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11344 = 3'h5 == state ? _GEN_10313 : ram_1_41; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11345 = 3'h5 == state ? _GEN_10314 : ram_1_42; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11346 = 3'h5 == state ? _GEN_10315 : ram_1_43; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11347 = 3'h5 == state ? _GEN_10316 : ram_1_44; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11348 = 3'h5 == state ? _GEN_10317 : ram_1_45; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11349 = 3'h5 == state ? _GEN_10318 : ram_1_46; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11350 = 3'h5 == state ? _GEN_10319 : ram_1_47; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11351 = 3'h5 == state ? _GEN_10320 : ram_1_48; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11352 = 3'h5 == state ? _GEN_10321 : ram_1_49; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11353 = 3'h5 == state ? _GEN_10322 : ram_1_50; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11354 = 3'h5 == state ? _GEN_10323 : ram_1_51; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11355 = 3'h5 == state ? _GEN_10324 : ram_1_52; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11356 = 3'h5 == state ? _GEN_10325 : ram_1_53; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11357 = 3'h5 == state ? _GEN_10326 : ram_1_54; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11358 = 3'h5 == state ? _GEN_10327 : ram_1_55; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11359 = 3'h5 == state ? _GEN_10328 : ram_1_56; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11360 = 3'h5 == state ? _GEN_10329 : ram_1_57; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11361 = 3'h5 == state ? _GEN_10330 : ram_1_58; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11362 = 3'h5 == state ? _GEN_10331 : ram_1_59; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11363 = 3'h5 == state ? _GEN_10332 : ram_1_60; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11364 = 3'h5 == state ? _GEN_10333 : ram_1_61; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11365 = 3'h5 == state ? _GEN_10334 : ram_1_62; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11366 = 3'h5 == state ? _GEN_10335 : ram_1_63; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11367 = 3'h5 == state ? _GEN_10336 : ram_1_64; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11368 = 3'h5 == state ? _GEN_10337 : ram_1_65; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11369 = 3'h5 == state ? _GEN_10338 : ram_1_66; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11370 = 3'h5 == state ? _GEN_10339 : ram_1_67; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11371 = 3'h5 == state ? _GEN_10340 : ram_1_68; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11372 = 3'h5 == state ? _GEN_10341 : ram_1_69; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11373 = 3'h5 == state ? _GEN_10342 : ram_1_70; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11374 = 3'h5 == state ? _GEN_10343 : ram_1_71; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11375 = 3'h5 == state ? _GEN_10344 : ram_1_72; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11376 = 3'h5 == state ? _GEN_10345 : ram_1_73; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11377 = 3'h5 == state ? _GEN_10346 : ram_1_74; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11378 = 3'h5 == state ? _GEN_10347 : ram_1_75; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11379 = 3'h5 == state ? _GEN_10348 : ram_1_76; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11380 = 3'h5 == state ? _GEN_10349 : ram_1_77; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11381 = 3'h5 == state ? _GEN_10350 : ram_1_78; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11382 = 3'h5 == state ? _GEN_10351 : ram_1_79; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11383 = 3'h5 == state ? _GEN_10352 : ram_1_80; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11384 = 3'h5 == state ? _GEN_10353 : ram_1_81; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11385 = 3'h5 == state ? _GEN_10354 : ram_1_82; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11386 = 3'h5 == state ? _GEN_10355 : ram_1_83; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11387 = 3'h5 == state ? _GEN_10356 : ram_1_84; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11388 = 3'h5 == state ? _GEN_10357 : ram_1_85; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11389 = 3'h5 == state ? _GEN_10358 : ram_1_86; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11390 = 3'h5 == state ? _GEN_10359 : ram_1_87; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11391 = 3'h5 == state ? _GEN_10360 : ram_1_88; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11392 = 3'h5 == state ? _GEN_10361 : ram_1_89; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11393 = 3'h5 == state ? _GEN_10362 : ram_1_90; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11394 = 3'h5 == state ? _GEN_10363 : ram_1_91; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11395 = 3'h5 == state ? _GEN_10364 : ram_1_92; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11396 = 3'h5 == state ? _GEN_10365 : ram_1_93; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11397 = 3'h5 == state ? _GEN_10366 : ram_1_94; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11398 = 3'h5 == state ? _GEN_10367 : ram_1_95; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11399 = 3'h5 == state ? _GEN_10368 : ram_1_96; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11400 = 3'h5 == state ? _GEN_10369 : ram_1_97; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11401 = 3'h5 == state ? _GEN_10370 : ram_1_98; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11402 = 3'h5 == state ? _GEN_10371 : ram_1_99; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11403 = 3'h5 == state ? _GEN_10372 : ram_1_100; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11404 = 3'h5 == state ? _GEN_10373 : ram_1_101; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11405 = 3'h5 == state ? _GEN_10374 : ram_1_102; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11406 = 3'h5 == state ? _GEN_10375 : ram_1_103; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11407 = 3'h5 == state ? _GEN_10376 : ram_1_104; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11408 = 3'h5 == state ? _GEN_10377 : ram_1_105; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11409 = 3'h5 == state ? _GEN_10378 : ram_1_106; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11410 = 3'h5 == state ? _GEN_10379 : ram_1_107; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11411 = 3'h5 == state ? _GEN_10380 : ram_1_108; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11412 = 3'h5 == state ? _GEN_10381 : ram_1_109; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11413 = 3'h5 == state ? _GEN_10382 : ram_1_110; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11414 = 3'h5 == state ? _GEN_10383 : ram_1_111; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11415 = 3'h5 == state ? _GEN_10384 : ram_1_112; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11416 = 3'h5 == state ? _GEN_10385 : ram_1_113; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11417 = 3'h5 == state ? _GEN_10386 : ram_1_114; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11418 = 3'h5 == state ? _GEN_10387 : ram_1_115; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11419 = 3'h5 == state ? _GEN_10388 : ram_1_116; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11420 = 3'h5 == state ? _GEN_10389 : ram_1_117; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11421 = 3'h5 == state ? _GEN_10390 : ram_1_118; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11422 = 3'h5 == state ? _GEN_10391 : ram_1_119; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11423 = 3'h5 == state ? _GEN_10392 : ram_1_120; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11424 = 3'h5 == state ? _GEN_10393 : ram_1_121; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11425 = 3'h5 == state ? _GEN_10394 : ram_1_122; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11426 = 3'h5 == state ? _GEN_10395 : ram_1_123; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11427 = 3'h5 == state ? _GEN_10396 : ram_1_124; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11428 = 3'h5 == state ? _GEN_10397 : ram_1_125; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11429 = 3'h5 == state ? _GEN_10398 : ram_1_126; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_11430 = 3'h5 == state ? _GEN_10399 : ram_1_127; // @[d_cache.scala 87:18 20:24]
  wire [31:0] _GEN_11431 = 3'h5 == state ? _GEN_10400 : tag_1_0; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11432 = 3'h5 == state ? _GEN_10401 : tag_1_1; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11433 = 3'h5 == state ? _GEN_10402 : tag_1_2; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11434 = 3'h5 == state ? _GEN_10403 : tag_1_3; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11435 = 3'h5 == state ? _GEN_10404 : tag_1_4; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11436 = 3'h5 == state ? _GEN_10405 : tag_1_5; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11437 = 3'h5 == state ? _GEN_10406 : tag_1_6; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11438 = 3'h5 == state ? _GEN_10407 : tag_1_7; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11439 = 3'h5 == state ? _GEN_10408 : tag_1_8; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11440 = 3'h5 == state ? _GEN_10409 : tag_1_9; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11441 = 3'h5 == state ? _GEN_10410 : tag_1_10; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11442 = 3'h5 == state ? _GEN_10411 : tag_1_11; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11443 = 3'h5 == state ? _GEN_10412 : tag_1_12; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11444 = 3'h5 == state ? _GEN_10413 : tag_1_13; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11445 = 3'h5 == state ? _GEN_10414 : tag_1_14; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11446 = 3'h5 == state ? _GEN_10415 : tag_1_15; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11447 = 3'h5 == state ? _GEN_10416 : tag_1_16; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11448 = 3'h5 == state ? _GEN_10417 : tag_1_17; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11449 = 3'h5 == state ? _GEN_10418 : tag_1_18; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11450 = 3'h5 == state ? _GEN_10419 : tag_1_19; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11451 = 3'h5 == state ? _GEN_10420 : tag_1_20; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11452 = 3'h5 == state ? _GEN_10421 : tag_1_21; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11453 = 3'h5 == state ? _GEN_10422 : tag_1_22; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11454 = 3'h5 == state ? _GEN_10423 : tag_1_23; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11455 = 3'h5 == state ? _GEN_10424 : tag_1_24; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11456 = 3'h5 == state ? _GEN_10425 : tag_1_25; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11457 = 3'h5 == state ? _GEN_10426 : tag_1_26; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11458 = 3'h5 == state ? _GEN_10427 : tag_1_27; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11459 = 3'h5 == state ? _GEN_10428 : tag_1_28; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11460 = 3'h5 == state ? _GEN_10429 : tag_1_29; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11461 = 3'h5 == state ? _GEN_10430 : tag_1_30; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11462 = 3'h5 == state ? _GEN_10431 : tag_1_31; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11463 = 3'h5 == state ? _GEN_10432 : tag_1_32; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11464 = 3'h5 == state ? _GEN_10433 : tag_1_33; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11465 = 3'h5 == state ? _GEN_10434 : tag_1_34; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11466 = 3'h5 == state ? _GEN_10435 : tag_1_35; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11467 = 3'h5 == state ? _GEN_10436 : tag_1_36; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11468 = 3'h5 == state ? _GEN_10437 : tag_1_37; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11469 = 3'h5 == state ? _GEN_10438 : tag_1_38; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11470 = 3'h5 == state ? _GEN_10439 : tag_1_39; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11471 = 3'h5 == state ? _GEN_10440 : tag_1_40; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11472 = 3'h5 == state ? _GEN_10441 : tag_1_41; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11473 = 3'h5 == state ? _GEN_10442 : tag_1_42; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11474 = 3'h5 == state ? _GEN_10443 : tag_1_43; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11475 = 3'h5 == state ? _GEN_10444 : tag_1_44; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11476 = 3'h5 == state ? _GEN_10445 : tag_1_45; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11477 = 3'h5 == state ? _GEN_10446 : tag_1_46; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11478 = 3'h5 == state ? _GEN_10447 : tag_1_47; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11479 = 3'h5 == state ? _GEN_10448 : tag_1_48; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11480 = 3'h5 == state ? _GEN_10449 : tag_1_49; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11481 = 3'h5 == state ? _GEN_10450 : tag_1_50; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11482 = 3'h5 == state ? _GEN_10451 : tag_1_51; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11483 = 3'h5 == state ? _GEN_10452 : tag_1_52; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11484 = 3'h5 == state ? _GEN_10453 : tag_1_53; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11485 = 3'h5 == state ? _GEN_10454 : tag_1_54; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11486 = 3'h5 == state ? _GEN_10455 : tag_1_55; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11487 = 3'h5 == state ? _GEN_10456 : tag_1_56; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11488 = 3'h5 == state ? _GEN_10457 : tag_1_57; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11489 = 3'h5 == state ? _GEN_10458 : tag_1_58; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11490 = 3'h5 == state ? _GEN_10459 : tag_1_59; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11491 = 3'h5 == state ? _GEN_10460 : tag_1_60; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11492 = 3'h5 == state ? _GEN_10461 : tag_1_61; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11493 = 3'h5 == state ? _GEN_10462 : tag_1_62; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11494 = 3'h5 == state ? _GEN_10463 : tag_1_63; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11495 = 3'h5 == state ? _GEN_10464 : tag_1_64; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11496 = 3'h5 == state ? _GEN_10465 : tag_1_65; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11497 = 3'h5 == state ? _GEN_10466 : tag_1_66; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11498 = 3'h5 == state ? _GEN_10467 : tag_1_67; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11499 = 3'h5 == state ? _GEN_10468 : tag_1_68; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11500 = 3'h5 == state ? _GEN_10469 : tag_1_69; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11501 = 3'h5 == state ? _GEN_10470 : tag_1_70; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11502 = 3'h5 == state ? _GEN_10471 : tag_1_71; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11503 = 3'h5 == state ? _GEN_10472 : tag_1_72; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11504 = 3'h5 == state ? _GEN_10473 : tag_1_73; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11505 = 3'h5 == state ? _GEN_10474 : tag_1_74; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11506 = 3'h5 == state ? _GEN_10475 : tag_1_75; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11507 = 3'h5 == state ? _GEN_10476 : tag_1_76; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11508 = 3'h5 == state ? _GEN_10477 : tag_1_77; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11509 = 3'h5 == state ? _GEN_10478 : tag_1_78; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11510 = 3'h5 == state ? _GEN_10479 : tag_1_79; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11511 = 3'h5 == state ? _GEN_10480 : tag_1_80; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11512 = 3'h5 == state ? _GEN_10481 : tag_1_81; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11513 = 3'h5 == state ? _GEN_10482 : tag_1_82; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11514 = 3'h5 == state ? _GEN_10483 : tag_1_83; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11515 = 3'h5 == state ? _GEN_10484 : tag_1_84; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11516 = 3'h5 == state ? _GEN_10485 : tag_1_85; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11517 = 3'h5 == state ? _GEN_10486 : tag_1_86; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11518 = 3'h5 == state ? _GEN_10487 : tag_1_87; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11519 = 3'h5 == state ? _GEN_10488 : tag_1_88; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11520 = 3'h5 == state ? _GEN_10489 : tag_1_89; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11521 = 3'h5 == state ? _GEN_10490 : tag_1_90; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11522 = 3'h5 == state ? _GEN_10491 : tag_1_91; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11523 = 3'h5 == state ? _GEN_10492 : tag_1_92; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11524 = 3'h5 == state ? _GEN_10493 : tag_1_93; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11525 = 3'h5 == state ? _GEN_10494 : tag_1_94; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11526 = 3'h5 == state ? _GEN_10495 : tag_1_95; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11527 = 3'h5 == state ? _GEN_10496 : tag_1_96; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11528 = 3'h5 == state ? _GEN_10497 : tag_1_97; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11529 = 3'h5 == state ? _GEN_10498 : tag_1_98; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11530 = 3'h5 == state ? _GEN_10499 : tag_1_99; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11531 = 3'h5 == state ? _GEN_10500 : tag_1_100; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11532 = 3'h5 == state ? _GEN_10501 : tag_1_101; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11533 = 3'h5 == state ? _GEN_10502 : tag_1_102; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11534 = 3'h5 == state ? _GEN_10503 : tag_1_103; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11535 = 3'h5 == state ? _GEN_10504 : tag_1_104; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11536 = 3'h5 == state ? _GEN_10505 : tag_1_105; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11537 = 3'h5 == state ? _GEN_10506 : tag_1_106; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11538 = 3'h5 == state ? _GEN_10507 : tag_1_107; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11539 = 3'h5 == state ? _GEN_10508 : tag_1_108; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11540 = 3'h5 == state ? _GEN_10509 : tag_1_109; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11541 = 3'h5 == state ? _GEN_10510 : tag_1_110; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11542 = 3'h5 == state ? _GEN_10511 : tag_1_111; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11543 = 3'h5 == state ? _GEN_10512 : tag_1_112; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11544 = 3'h5 == state ? _GEN_10513 : tag_1_113; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11545 = 3'h5 == state ? _GEN_10514 : tag_1_114; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11546 = 3'h5 == state ? _GEN_10515 : tag_1_115; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11547 = 3'h5 == state ? _GEN_10516 : tag_1_116; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11548 = 3'h5 == state ? _GEN_10517 : tag_1_117; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11549 = 3'h5 == state ? _GEN_10518 : tag_1_118; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11550 = 3'h5 == state ? _GEN_10519 : tag_1_119; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11551 = 3'h5 == state ? _GEN_10520 : tag_1_120; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11552 = 3'h5 == state ? _GEN_10521 : tag_1_121; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11553 = 3'h5 == state ? _GEN_10522 : tag_1_122; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11554 = 3'h5 == state ? _GEN_10523 : tag_1_123; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11555 = 3'h5 == state ? _GEN_10524 : tag_1_124; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11556 = 3'h5 == state ? _GEN_10525 : tag_1_125; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11557 = 3'h5 == state ? _GEN_10526 : tag_1_126; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_11558 = 3'h5 == state ? _GEN_10527 : tag_1_127; // @[d_cache.scala 87:18 29:24]
  wire  _GEN_11559 = 3'h5 == state ? _GEN_10528 : valid_1_0; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11560 = 3'h5 == state ? _GEN_10529 : valid_1_1; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11561 = 3'h5 == state ? _GEN_10530 : valid_1_2; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11562 = 3'h5 == state ? _GEN_10531 : valid_1_3; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11563 = 3'h5 == state ? _GEN_10532 : valid_1_4; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11564 = 3'h5 == state ? _GEN_10533 : valid_1_5; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11565 = 3'h5 == state ? _GEN_10534 : valid_1_6; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11566 = 3'h5 == state ? _GEN_10535 : valid_1_7; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11567 = 3'h5 == state ? _GEN_10536 : valid_1_8; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11568 = 3'h5 == state ? _GEN_10537 : valid_1_9; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11569 = 3'h5 == state ? _GEN_10538 : valid_1_10; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11570 = 3'h5 == state ? _GEN_10539 : valid_1_11; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11571 = 3'h5 == state ? _GEN_10540 : valid_1_12; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11572 = 3'h5 == state ? _GEN_10541 : valid_1_13; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11573 = 3'h5 == state ? _GEN_10542 : valid_1_14; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11574 = 3'h5 == state ? _GEN_10543 : valid_1_15; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11575 = 3'h5 == state ? _GEN_10544 : valid_1_16; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11576 = 3'h5 == state ? _GEN_10545 : valid_1_17; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11577 = 3'h5 == state ? _GEN_10546 : valid_1_18; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11578 = 3'h5 == state ? _GEN_10547 : valid_1_19; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11579 = 3'h5 == state ? _GEN_10548 : valid_1_20; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11580 = 3'h5 == state ? _GEN_10549 : valid_1_21; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11581 = 3'h5 == state ? _GEN_10550 : valid_1_22; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11582 = 3'h5 == state ? _GEN_10551 : valid_1_23; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11583 = 3'h5 == state ? _GEN_10552 : valid_1_24; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11584 = 3'h5 == state ? _GEN_10553 : valid_1_25; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11585 = 3'h5 == state ? _GEN_10554 : valid_1_26; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11586 = 3'h5 == state ? _GEN_10555 : valid_1_27; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11587 = 3'h5 == state ? _GEN_10556 : valid_1_28; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11588 = 3'h5 == state ? _GEN_10557 : valid_1_29; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11589 = 3'h5 == state ? _GEN_10558 : valid_1_30; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11590 = 3'h5 == state ? _GEN_10559 : valid_1_31; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11591 = 3'h5 == state ? _GEN_10560 : valid_1_32; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11592 = 3'h5 == state ? _GEN_10561 : valid_1_33; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11593 = 3'h5 == state ? _GEN_10562 : valid_1_34; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11594 = 3'h5 == state ? _GEN_10563 : valid_1_35; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11595 = 3'h5 == state ? _GEN_10564 : valid_1_36; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11596 = 3'h5 == state ? _GEN_10565 : valid_1_37; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11597 = 3'h5 == state ? _GEN_10566 : valid_1_38; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11598 = 3'h5 == state ? _GEN_10567 : valid_1_39; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11599 = 3'h5 == state ? _GEN_10568 : valid_1_40; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11600 = 3'h5 == state ? _GEN_10569 : valid_1_41; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11601 = 3'h5 == state ? _GEN_10570 : valid_1_42; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11602 = 3'h5 == state ? _GEN_10571 : valid_1_43; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11603 = 3'h5 == state ? _GEN_10572 : valid_1_44; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11604 = 3'h5 == state ? _GEN_10573 : valid_1_45; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11605 = 3'h5 == state ? _GEN_10574 : valid_1_46; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11606 = 3'h5 == state ? _GEN_10575 : valid_1_47; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11607 = 3'h5 == state ? _GEN_10576 : valid_1_48; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11608 = 3'h5 == state ? _GEN_10577 : valid_1_49; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11609 = 3'h5 == state ? _GEN_10578 : valid_1_50; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11610 = 3'h5 == state ? _GEN_10579 : valid_1_51; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11611 = 3'h5 == state ? _GEN_10580 : valid_1_52; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11612 = 3'h5 == state ? _GEN_10581 : valid_1_53; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11613 = 3'h5 == state ? _GEN_10582 : valid_1_54; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11614 = 3'h5 == state ? _GEN_10583 : valid_1_55; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11615 = 3'h5 == state ? _GEN_10584 : valid_1_56; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11616 = 3'h5 == state ? _GEN_10585 : valid_1_57; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11617 = 3'h5 == state ? _GEN_10586 : valid_1_58; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11618 = 3'h5 == state ? _GEN_10587 : valid_1_59; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11619 = 3'h5 == state ? _GEN_10588 : valid_1_60; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11620 = 3'h5 == state ? _GEN_10589 : valid_1_61; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11621 = 3'h5 == state ? _GEN_10590 : valid_1_62; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11622 = 3'h5 == state ? _GEN_10591 : valid_1_63; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11623 = 3'h5 == state ? _GEN_10592 : valid_1_64; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11624 = 3'h5 == state ? _GEN_10593 : valid_1_65; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11625 = 3'h5 == state ? _GEN_10594 : valid_1_66; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11626 = 3'h5 == state ? _GEN_10595 : valid_1_67; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11627 = 3'h5 == state ? _GEN_10596 : valid_1_68; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11628 = 3'h5 == state ? _GEN_10597 : valid_1_69; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11629 = 3'h5 == state ? _GEN_10598 : valid_1_70; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11630 = 3'h5 == state ? _GEN_10599 : valid_1_71; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11631 = 3'h5 == state ? _GEN_10600 : valid_1_72; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11632 = 3'h5 == state ? _GEN_10601 : valid_1_73; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11633 = 3'h5 == state ? _GEN_10602 : valid_1_74; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11634 = 3'h5 == state ? _GEN_10603 : valid_1_75; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11635 = 3'h5 == state ? _GEN_10604 : valid_1_76; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11636 = 3'h5 == state ? _GEN_10605 : valid_1_77; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11637 = 3'h5 == state ? _GEN_10606 : valid_1_78; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11638 = 3'h5 == state ? _GEN_10607 : valid_1_79; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11639 = 3'h5 == state ? _GEN_10608 : valid_1_80; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11640 = 3'h5 == state ? _GEN_10609 : valid_1_81; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11641 = 3'h5 == state ? _GEN_10610 : valid_1_82; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11642 = 3'h5 == state ? _GEN_10611 : valid_1_83; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11643 = 3'h5 == state ? _GEN_10612 : valid_1_84; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11644 = 3'h5 == state ? _GEN_10613 : valid_1_85; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11645 = 3'h5 == state ? _GEN_10614 : valid_1_86; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11646 = 3'h5 == state ? _GEN_10615 : valid_1_87; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11647 = 3'h5 == state ? _GEN_10616 : valid_1_88; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11648 = 3'h5 == state ? _GEN_10617 : valid_1_89; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11649 = 3'h5 == state ? _GEN_10618 : valid_1_90; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11650 = 3'h5 == state ? _GEN_10619 : valid_1_91; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11651 = 3'h5 == state ? _GEN_10620 : valid_1_92; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11652 = 3'h5 == state ? _GEN_10621 : valid_1_93; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11653 = 3'h5 == state ? _GEN_10622 : valid_1_94; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11654 = 3'h5 == state ? _GEN_10623 : valid_1_95; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11655 = 3'h5 == state ? _GEN_10624 : valid_1_96; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11656 = 3'h5 == state ? _GEN_10625 : valid_1_97; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11657 = 3'h5 == state ? _GEN_10626 : valid_1_98; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11658 = 3'h5 == state ? _GEN_10627 : valid_1_99; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11659 = 3'h5 == state ? _GEN_10628 : valid_1_100; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11660 = 3'h5 == state ? _GEN_10629 : valid_1_101; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11661 = 3'h5 == state ? _GEN_10630 : valid_1_102; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11662 = 3'h5 == state ? _GEN_10631 : valid_1_103; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11663 = 3'h5 == state ? _GEN_10632 : valid_1_104; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11664 = 3'h5 == state ? _GEN_10633 : valid_1_105; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11665 = 3'h5 == state ? _GEN_10634 : valid_1_106; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11666 = 3'h5 == state ? _GEN_10635 : valid_1_107; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11667 = 3'h5 == state ? _GEN_10636 : valid_1_108; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11668 = 3'h5 == state ? _GEN_10637 : valid_1_109; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11669 = 3'h5 == state ? _GEN_10638 : valid_1_110; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11670 = 3'h5 == state ? _GEN_10639 : valid_1_111; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11671 = 3'h5 == state ? _GEN_10640 : valid_1_112; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11672 = 3'h5 == state ? _GEN_10641 : valid_1_113; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11673 = 3'h5 == state ? _GEN_10642 : valid_1_114; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11674 = 3'h5 == state ? _GEN_10643 : valid_1_115; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11675 = 3'h5 == state ? _GEN_10644 : valid_1_116; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11676 = 3'h5 == state ? _GEN_10645 : valid_1_117; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11677 = 3'h5 == state ? _GEN_10646 : valid_1_118; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11678 = 3'h5 == state ? _GEN_10647 : valid_1_119; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11679 = 3'h5 == state ? _GEN_10648 : valid_1_120; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11680 = 3'h5 == state ? _GEN_10649 : valid_1_121; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11681 = 3'h5 == state ? _GEN_10650 : valid_1_122; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11682 = 3'h5 == state ? _GEN_10651 : valid_1_123; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11683 = 3'h5 == state ? _GEN_10652 : valid_1_124; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11684 = 3'h5 == state ? _GEN_10653 : valid_1_125; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11685 = 3'h5 == state ? _GEN_10654 : valid_1_126; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_11686 = 3'h5 == state ? _GEN_10655 : valid_1_127; // @[d_cache.scala 87:18 31:26]
  wire [63:0] _GEN_11687 = 3'h5 == state ? _GEN_10656 : write_back_data; // @[d_cache.scala 87:18 37:34]
  wire [41:0] _GEN_11688 = 3'h5 == state ? _GEN_10657 : {{10'd0}, write_back_addr}; // @[d_cache.scala 87:18 38:34]
  wire  _GEN_11689 = 3'h5 == state ? _GEN_10658 : dirty_0_0; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11690 = 3'h5 == state ? _GEN_10659 : dirty_0_1; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11691 = 3'h5 == state ? _GEN_10660 : dirty_0_2; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11692 = 3'h5 == state ? _GEN_10661 : dirty_0_3; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11693 = 3'h5 == state ? _GEN_10662 : dirty_0_4; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11694 = 3'h5 == state ? _GEN_10663 : dirty_0_5; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11695 = 3'h5 == state ? _GEN_10664 : dirty_0_6; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11696 = 3'h5 == state ? _GEN_10665 : dirty_0_7; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11697 = 3'h5 == state ? _GEN_10666 : dirty_0_8; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11698 = 3'h5 == state ? _GEN_10667 : dirty_0_9; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11699 = 3'h5 == state ? _GEN_10668 : dirty_0_10; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11700 = 3'h5 == state ? _GEN_10669 : dirty_0_11; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11701 = 3'h5 == state ? _GEN_10670 : dirty_0_12; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11702 = 3'h5 == state ? _GEN_10671 : dirty_0_13; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11703 = 3'h5 == state ? _GEN_10672 : dirty_0_14; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11704 = 3'h5 == state ? _GEN_10673 : dirty_0_15; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11705 = 3'h5 == state ? _GEN_10674 : dirty_0_16; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11706 = 3'h5 == state ? _GEN_10675 : dirty_0_17; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11707 = 3'h5 == state ? _GEN_10676 : dirty_0_18; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11708 = 3'h5 == state ? _GEN_10677 : dirty_0_19; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11709 = 3'h5 == state ? _GEN_10678 : dirty_0_20; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11710 = 3'h5 == state ? _GEN_10679 : dirty_0_21; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11711 = 3'h5 == state ? _GEN_10680 : dirty_0_22; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11712 = 3'h5 == state ? _GEN_10681 : dirty_0_23; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11713 = 3'h5 == state ? _GEN_10682 : dirty_0_24; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11714 = 3'h5 == state ? _GEN_10683 : dirty_0_25; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11715 = 3'h5 == state ? _GEN_10684 : dirty_0_26; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11716 = 3'h5 == state ? _GEN_10685 : dirty_0_27; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11717 = 3'h5 == state ? _GEN_10686 : dirty_0_28; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11718 = 3'h5 == state ? _GEN_10687 : dirty_0_29; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11719 = 3'h5 == state ? _GEN_10688 : dirty_0_30; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11720 = 3'h5 == state ? _GEN_10689 : dirty_0_31; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11721 = 3'h5 == state ? _GEN_10690 : dirty_0_32; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11722 = 3'h5 == state ? _GEN_10691 : dirty_0_33; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11723 = 3'h5 == state ? _GEN_10692 : dirty_0_34; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11724 = 3'h5 == state ? _GEN_10693 : dirty_0_35; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11725 = 3'h5 == state ? _GEN_10694 : dirty_0_36; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11726 = 3'h5 == state ? _GEN_10695 : dirty_0_37; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11727 = 3'h5 == state ? _GEN_10696 : dirty_0_38; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11728 = 3'h5 == state ? _GEN_10697 : dirty_0_39; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11729 = 3'h5 == state ? _GEN_10698 : dirty_0_40; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11730 = 3'h5 == state ? _GEN_10699 : dirty_0_41; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11731 = 3'h5 == state ? _GEN_10700 : dirty_0_42; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11732 = 3'h5 == state ? _GEN_10701 : dirty_0_43; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11733 = 3'h5 == state ? _GEN_10702 : dirty_0_44; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11734 = 3'h5 == state ? _GEN_10703 : dirty_0_45; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11735 = 3'h5 == state ? _GEN_10704 : dirty_0_46; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11736 = 3'h5 == state ? _GEN_10705 : dirty_0_47; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11737 = 3'h5 == state ? _GEN_10706 : dirty_0_48; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11738 = 3'h5 == state ? _GEN_10707 : dirty_0_49; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11739 = 3'h5 == state ? _GEN_10708 : dirty_0_50; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11740 = 3'h5 == state ? _GEN_10709 : dirty_0_51; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11741 = 3'h5 == state ? _GEN_10710 : dirty_0_52; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11742 = 3'h5 == state ? _GEN_10711 : dirty_0_53; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11743 = 3'h5 == state ? _GEN_10712 : dirty_0_54; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11744 = 3'h5 == state ? _GEN_10713 : dirty_0_55; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11745 = 3'h5 == state ? _GEN_10714 : dirty_0_56; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11746 = 3'h5 == state ? _GEN_10715 : dirty_0_57; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11747 = 3'h5 == state ? _GEN_10716 : dirty_0_58; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11748 = 3'h5 == state ? _GEN_10717 : dirty_0_59; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11749 = 3'h5 == state ? _GEN_10718 : dirty_0_60; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11750 = 3'h5 == state ? _GEN_10719 : dirty_0_61; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11751 = 3'h5 == state ? _GEN_10720 : dirty_0_62; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11752 = 3'h5 == state ? _GEN_10721 : dirty_0_63; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11753 = 3'h5 == state ? _GEN_10722 : dirty_0_64; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11754 = 3'h5 == state ? _GEN_10723 : dirty_0_65; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11755 = 3'h5 == state ? _GEN_10724 : dirty_0_66; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11756 = 3'h5 == state ? _GEN_10725 : dirty_0_67; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11757 = 3'h5 == state ? _GEN_10726 : dirty_0_68; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11758 = 3'h5 == state ? _GEN_10727 : dirty_0_69; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11759 = 3'h5 == state ? _GEN_10728 : dirty_0_70; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11760 = 3'h5 == state ? _GEN_10729 : dirty_0_71; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11761 = 3'h5 == state ? _GEN_10730 : dirty_0_72; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11762 = 3'h5 == state ? _GEN_10731 : dirty_0_73; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11763 = 3'h5 == state ? _GEN_10732 : dirty_0_74; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11764 = 3'h5 == state ? _GEN_10733 : dirty_0_75; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11765 = 3'h5 == state ? _GEN_10734 : dirty_0_76; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11766 = 3'h5 == state ? _GEN_10735 : dirty_0_77; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11767 = 3'h5 == state ? _GEN_10736 : dirty_0_78; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11768 = 3'h5 == state ? _GEN_10737 : dirty_0_79; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11769 = 3'h5 == state ? _GEN_10738 : dirty_0_80; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11770 = 3'h5 == state ? _GEN_10739 : dirty_0_81; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11771 = 3'h5 == state ? _GEN_10740 : dirty_0_82; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11772 = 3'h5 == state ? _GEN_10741 : dirty_0_83; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11773 = 3'h5 == state ? _GEN_10742 : dirty_0_84; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11774 = 3'h5 == state ? _GEN_10743 : dirty_0_85; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11775 = 3'h5 == state ? _GEN_10744 : dirty_0_86; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11776 = 3'h5 == state ? _GEN_10745 : dirty_0_87; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11777 = 3'h5 == state ? _GEN_10746 : dirty_0_88; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11778 = 3'h5 == state ? _GEN_10747 : dirty_0_89; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11779 = 3'h5 == state ? _GEN_10748 : dirty_0_90; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11780 = 3'h5 == state ? _GEN_10749 : dirty_0_91; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11781 = 3'h5 == state ? _GEN_10750 : dirty_0_92; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11782 = 3'h5 == state ? _GEN_10751 : dirty_0_93; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11783 = 3'h5 == state ? _GEN_10752 : dirty_0_94; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11784 = 3'h5 == state ? _GEN_10753 : dirty_0_95; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11785 = 3'h5 == state ? _GEN_10754 : dirty_0_96; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11786 = 3'h5 == state ? _GEN_10755 : dirty_0_97; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11787 = 3'h5 == state ? _GEN_10756 : dirty_0_98; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11788 = 3'h5 == state ? _GEN_10757 : dirty_0_99; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11789 = 3'h5 == state ? _GEN_10758 : dirty_0_100; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11790 = 3'h5 == state ? _GEN_10759 : dirty_0_101; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11791 = 3'h5 == state ? _GEN_10760 : dirty_0_102; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11792 = 3'h5 == state ? _GEN_10761 : dirty_0_103; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11793 = 3'h5 == state ? _GEN_10762 : dirty_0_104; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11794 = 3'h5 == state ? _GEN_10763 : dirty_0_105; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11795 = 3'h5 == state ? _GEN_10764 : dirty_0_106; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11796 = 3'h5 == state ? _GEN_10765 : dirty_0_107; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11797 = 3'h5 == state ? _GEN_10766 : dirty_0_108; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11798 = 3'h5 == state ? _GEN_10767 : dirty_0_109; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11799 = 3'h5 == state ? _GEN_10768 : dirty_0_110; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11800 = 3'h5 == state ? _GEN_10769 : dirty_0_111; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11801 = 3'h5 == state ? _GEN_10770 : dirty_0_112; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11802 = 3'h5 == state ? _GEN_10771 : dirty_0_113; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11803 = 3'h5 == state ? _GEN_10772 : dirty_0_114; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11804 = 3'h5 == state ? _GEN_10773 : dirty_0_115; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11805 = 3'h5 == state ? _GEN_10774 : dirty_0_116; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11806 = 3'h5 == state ? _GEN_10775 : dirty_0_117; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11807 = 3'h5 == state ? _GEN_10776 : dirty_0_118; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11808 = 3'h5 == state ? _GEN_10777 : dirty_0_119; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11809 = 3'h5 == state ? _GEN_10778 : dirty_0_120; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11810 = 3'h5 == state ? _GEN_10779 : dirty_0_121; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11811 = 3'h5 == state ? _GEN_10780 : dirty_0_122; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11812 = 3'h5 == state ? _GEN_10781 : dirty_0_123; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11813 = 3'h5 == state ? _GEN_10782 : dirty_0_124; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11814 = 3'h5 == state ? _GEN_10783 : dirty_0_125; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11815 = 3'h5 == state ? _GEN_10784 : dirty_0_126; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11816 = 3'h5 == state ? _GEN_10785 : dirty_0_127; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_11817 = 3'h5 == state ? _GEN_10786 : dirty_1_0; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11818 = 3'h5 == state ? _GEN_10787 : dirty_1_1; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11819 = 3'h5 == state ? _GEN_10788 : dirty_1_2; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11820 = 3'h5 == state ? _GEN_10789 : dirty_1_3; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11821 = 3'h5 == state ? _GEN_10790 : dirty_1_4; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11822 = 3'h5 == state ? _GEN_10791 : dirty_1_5; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11823 = 3'h5 == state ? _GEN_10792 : dirty_1_6; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11824 = 3'h5 == state ? _GEN_10793 : dirty_1_7; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11825 = 3'h5 == state ? _GEN_10794 : dirty_1_8; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11826 = 3'h5 == state ? _GEN_10795 : dirty_1_9; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11827 = 3'h5 == state ? _GEN_10796 : dirty_1_10; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11828 = 3'h5 == state ? _GEN_10797 : dirty_1_11; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11829 = 3'h5 == state ? _GEN_10798 : dirty_1_12; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11830 = 3'h5 == state ? _GEN_10799 : dirty_1_13; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11831 = 3'h5 == state ? _GEN_10800 : dirty_1_14; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11832 = 3'h5 == state ? _GEN_10801 : dirty_1_15; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11833 = 3'h5 == state ? _GEN_10802 : dirty_1_16; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11834 = 3'h5 == state ? _GEN_10803 : dirty_1_17; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11835 = 3'h5 == state ? _GEN_10804 : dirty_1_18; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11836 = 3'h5 == state ? _GEN_10805 : dirty_1_19; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11837 = 3'h5 == state ? _GEN_10806 : dirty_1_20; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11838 = 3'h5 == state ? _GEN_10807 : dirty_1_21; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11839 = 3'h5 == state ? _GEN_10808 : dirty_1_22; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11840 = 3'h5 == state ? _GEN_10809 : dirty_1_23; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11841 = 3'h5 == state ? _GEN_10810 : dirty_1_24; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11842 = 3'h5 == state ? _GEN_10811 : dirty_1_25; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11843 = 3'h5 == state ? _GEN_10812 : dirty_1_26; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11844 = 3'h5 == state ? _GEN_10813 : dirty_1_27; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11845 = 3'h5 == state ? _GEN_10814 : dirty_1_28; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11846 = 3'h5 == state ? _GEN_10815 : dirty_1_29; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11847 = 3'h5 == state ? _GEN_10816 : dirty_1_30; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11848 = 3'h5 == state ? _GEN_10817 : dirty_1_31; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11849 = 3'h5 == state ? _GEN_10818 : dirty_1_32; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11850 = 3'h5 == state ? _GEN_10819 : dirty_1_33; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11851 = 3'h5 == state ? _GEN_10820 : dirty_1_34; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11852 = 3'h5 == state ? _GEN_10821 : dirty_1_35; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11853 = 3'h5 == state ? _GEN_10822 : dirty_1_36; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11854 = 3'h5 == state ? _GEN_10823 : dirty_1_37; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11855 = 3'h5 == state ? _GEN_10824 : dirty_1_38; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11856 = 3'h5 == state ? _GEN_10825 : dirty_1_39; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11857 = 3'h5 == state ? _GEN_10826 : dirty_1_40; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11858 = 3'h5 == state ? _GEN_10827 : dirty_1_41; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11859 = 3'h5 == state ? _GEN_10828 : dirty_1_42; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11860 = 3'h5 == state ? _GEN_10829 : dirty_1_43; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11861 = 3'h5 == state ? _GEN_10830 : dirty_1_44; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11862 = 3'h5 == state ? _GEN_10831 : dirty_1_45; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11863 = 3'h5 == state ? _GEN_10832 : dirty_1_46; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11864 = 3'h5 == state ? _GEN_10833 : dirty_1_47; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11865 = 3'h5 == state ? _GEN_10834 : dirty_1_48; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11866 = 3'h5 == state ? _GEN_10835 : dirty_1_49; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11867 = 3'h5 == state ? _GEN_10836 : dirty_1_50; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11868 = 3'h5 == state ? _GEN_10837 : dirty_1_51; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11869 = 3'h5 == state ? _GEN_10838 : dirty_1_52; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11870 = 3'h5 == state ? _GEN_10839 : dirty_1_53; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11871 = 3'h5 == state ? _GEN_10840 : dirty_1_54; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11872 = 3'h5 == state ? _GEN_10841 : dirty_1_55; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11873 = 3'h5 == state ? _GEN_10842 : dirty_1_56; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11874 = 3'h5 == state ? _GEN_10843 : dirty_1_57; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11875 = 3'h5 == state ? _GEN_10844 : dirty_1_58; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11876 = 3'h5 == state ? _GEN_10845 : dirty_1_59; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11877 = 3'h5 == state ? _GEN_10846 : dirty_1_60; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11878 = 3'h5 == state ? _GEN_10847 : dirty_1_61; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11879 = 3'h5 == state ? _GEN_10848 : dirty_1_62; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11880 = 3'h5 == state ? _GEN_10849 : dirty_1_63; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11881 = 3'h5 == state ? _GEN_10850 : dirty_1_64; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11882 = 3'h5 == state ? _GEN_10851 : dirty_1_65; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11883 = 3'h5 == state ? _GEN_10852 : dirty_1_66; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11884 = 3'h5 == state ? _GEN_10853 : dirty_1_67; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11885 = 3'h5 == state ? _GEN_10854 : dirty_1_68; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11886 = 3'h5 == state ? _GEN_10855 : dirty_1_69; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11887 = 3'h5 == state ? _GEN_10856 : dirty_1_70; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11888 = 3'h5 == state ? _GEN_10857 : dirty_1_71; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11889 = 3'h5 == state ? _GEN_10858 : dirty_1_72; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11890 = 3'h5 == state ? _GEN_10859 : dirty_1_73; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11891 = 3'h5 == state ? _GEN_10860 : dirty_1_74; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11892 = 3'h5 == state ? _GEN_10861 : dirty_1_75; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11893 = 3'h5 == state ? _GEN_10862 : dirty_1_76; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11894 = 3'h5 == state ? _GEN_10863 : dirty_1_77; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11895 = 3'h5 == state ? _GEN_10864 : dirty_1_78; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11896 = 3'h5 == state ? _GEN_10865 : dirty_1_79; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11897 = 3'h5 == state ? _GEN_10866 : dirty_1_80; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11898 = 3'h5 == state ? _GEN_10867 : dirty_1_81; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11899 = 3'h5 == state ? _GEN_10868 : dirty_1_82; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11900 = 3'h5 == state ? _GEN_10869 : dirty_1_83; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11901 = 3'h5 == state ? _GEN_10870 : dirty_1_84; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11902 = 3'h5 == state ? _GEN_10871 : dirty_1_85; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11903 = 3'h5 == state ? _GEN_10872 : dirty_1_86; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11904 = 3'h5 == state ? _GEN_10873 : dirty_1_87; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11905 = 3'h5 == state ? _GEN_10874 : dirty_1_88; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11906 = 3'h5 == state ? _GEN_10875 : dirty_1_89; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11907 = 3'h5 == state ? _GEN_10876 : dirty_1_90; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11908 = 3'h5 == state ? _GEN_10877 : dirty_1_91; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11909 = 3'h5 == state ? _GEN_10878 : dirty_1_92; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11910 = 3'h5 == state ? _GEN_10879 : dirty_1_93; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11911 = 3'h5 == state ? _GEN_10880 : dirty_1_94; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11912 = 3'h5 == state ? _GEN_10881 : dirty_1_95; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11913 = 3'h5 == state ? _GEN_10882 : dirty_1_96; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11914 = 3'h5 == state ? _GEN_10883 : dirty_1_97; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11915 = 3'h5 == state ? _GEN_10884 : dirty_1_98; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11916 = 3'h5 == state ? _GEN_10885 : dirty_1_99; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11917 = 3'h5 == state ? _GEN_10886 : dirty_1_100; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11918 = 3'h5 == state ? _GEN_10887 : dirty_1_101; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11919 = 3'h5 == state ? _GEN_10888 : dirty_1_102; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11920 = 3'h5 == state ? _GEN_10889 : dirty_1_103; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11921 = 3'h5 == state ? _GEN_10890 : dirty_1_104; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11922 = 3'h5 == state ? _GEN_10891 : dirty_1_105; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11923 = 3'h5 == state ? _GEN_10892 : dirty_1_106; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11924 = 3'h5 == state ? _GEN_10893 : dirty_1_107; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11925 = 3'h5 == state ? _GEN_10894 : dirty_1_108; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11926 = 3'h5 == state ? _GEN_10895 : dirty_1_109; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11927 = 3'h5 == state ? _GEN_10896 : dirty_1_110; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11928 = 3'h5 == state ? _GEN_10897 : dirty_1_111; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11929 = 3'h5 == state ? _GEN_10898 : dirty_1_112; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11930 = 3'h5 == state ? _GEN_10899 : dirty_1_113; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11931 = 3'h5 == state ? _GEN_10900 : dirty_1_114; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11932 = 3'h5 == state ? _GEN_10901 : dirty_1_115; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11933 = 3'h5 == state ? _GEN_10902 : dirty_1_116; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11934 = 3'h5 == state ? _GEN_10903 : dirty_1_117; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11935 = 3'h5 == state ? _GEN_10904 : dirty_1_118; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11936 = 3'h5 == state ? _GEN_10905 : dirty_1_119; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11937 = 3'h5 == state ? _GEN_10906 : dirty_1_120; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11938 = 3'h5 == state ? _GEN_10907 : dirty_1_121; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11939 = 3'h5 == state ? _GEN_10908 : dirty_1_122; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11940 = 3'h5 == state ? _GEN_10909 : dirty_1_123; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11941 = 3'h5 == state ? _GEN_10910 : dirty_1_124; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11942 = 3'h5 == state ? _GEN_10911 : dirty_1_125; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11943 = 3'h5 == state ? _GEN_10912 : dirty_1_126; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_11944 = 3'h5 == state ? _GEN_10913 : dirty_1_127; // @[d_cache.scala 87:18 33:26]
  wire [2:0] _GEN_11945 = 3'h4 == state ? _GEN_4237 : _GEN_10917; // @[d_cache.scala 87:18]
  wire [63:0] _GEN_11946 = 3'h4 == state ? ram_0_0 : _GEN_10918; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11947 = 3'h4 == state ? ram_0_1 : _GEN_10919; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11948 = 3'h4 == state ? ram_0_2 : _GEN_10920; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11949 = 3'h4 == state ? ram_0_3 : _GEN_10921; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11950 = 3'h4 == state ? ram_0_4 : _GEN_10922; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11951 = 3'h4 == state ? ram_0_5 : _GEN_10923; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11952 = 3'h4 == state ? ram_0_6 : _GEN_10924; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11953 = 3'h4 == state ? ram_0_7 : _GEN_10925; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11954 = 3'h4 == state ? ram_0_8 : _GEN_10926; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11955 = 3'h4 == state ? ram_0_9 : _GEN_10927; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11956 = 3'h4 == state ? ram_0_10 : _GEN_10928; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11957 = 3'h4 == state ? ram_0_11 : _GEN_10929; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11958 = 3'h4 == state ? ram_0_12 : _GEN_10930; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11959 = 3'h4 == state ? ram_0_13 : _GEN_10931; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11960 = 3'h4 == state ? ram_0_14 : _GEN_10932; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11961 = 3'h4 == state ? ram_0_15 : _GEN_10933; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11962 = 3'h4 == state ? ram_0_16 : _GEN_10934; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11963 = 3'h4 == state ? ram_0_17 : _GEN_10935; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11964 = 3'h4 == state ? ram_0_18 : _GEN_10936; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11965 = 3'h4 == state ? ram_0_19 : _GEN_10937; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11966 = 3'h4 == state ? ram_0_20 : _GEN_10938; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11967 = 3'h4 == state ? ram_0_21 : _GEN_10939; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11968 = 3'h4 == state ? ram_0_22 : _GEN_10940; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11969 = 3'h4 == state ? ram_0_23 : _GEN_10941; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11970 = 3'h4 == state ? ram_0_24 : _GEN_10942; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11971 = 3'h4 == state ? ram_0_25 : _GEN_10943; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11972 = 3'h4 == state ? ram_0_26 : _GEN_10944; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11973 = 3'h4 == state ? ram_0_27 : _GEN_10945; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11974 = 3'h4 == state ? ram_0_28 : _GEN_10946; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11975 = 3'h4 == state ? ram_0_29 : _GEN_10947; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11976 = 3'h4 == state ? ram_0_30 : _GEN_10948; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11977 = 3'h4 == state ? ram_0_31 : _GEN_10949; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11978 = 3'h4 == state ? ram_0_32 : _GEN_10950; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11979 = 3'h4 == state ? ram_0_33 : _GEN_10951; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11980 = 3'h4 == state ? ram_0_34 : _GEN_10952; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11981 = 3'h4 == state ? ram_0_35 : _GEN_10953; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11982 = 3'h4 == state ? ram_0_36 : _GEN_10954; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11983 = 3'h4 == state ? ram_0_37 : _GEN_10955; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11984 = 3'h4 == state ? ram_0_38 : _GEN_10956; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11985 = 3'h4 == state ? ram_0_39 : _GEN_10957; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11986 = 3'h4 == state ? ram_0_40 : _GEN_10958; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11987 = 3'h4 == state ? ram_0_41 : _GEN_10959; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11988 = 3'h4 == state ? ram_0_42 : _GEN_10960; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11989 = 3'h4 == state ? ram_0_43 : _GEN_10961; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11990 = 3'h4 == state ? ram_0_44 : _GEN_10962; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11991 = 3'h4 == state ? ram_0_45 : _GEN_10963; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11992 = 3'h4 == state ? ram_0_46 : _GEN_10964; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11993 = 3'h4 == state ? ram_0_47 : _GEN_10965; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11994 = 3'h4 == state ? ram_0_48 : _GEN_10966; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11995 = 3'h4 == state ? ram_0_49 : _GEN_10967; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11996 = 3'h4 == state ? ram_0_50 : _GEN_10968; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11997 = 3'h4 == state ? ram_0_51 : _GEN_10969; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11998 = 3'h4 == state ? ram_0_52 : _GEN_10970; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_11999 = 3'h4 == state ? ram_0_53 : _GEN_10971; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12000 = 3'h4 == state ? ram_0_54 : _GEN_10972; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12001 = 3'h4 == state ? ram_0_55 : _GEN_10973; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12002 = 3'h4 == state ? ram_0_56 : _GEN_10974; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12003 = 3'h4 == state ? ram_0_57 : _GEN_10975; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12004 = 3'h4 == state ? ram_0_58 : _GEN_10976; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12005 = 3'h4 == state ? ram_0_59 : _GEN_10977; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12006 = 3'h4 == state ? ram_0_60 : _GEN_10978; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12007 = 3'h4 == state ? ram_0_61 : _GEN_10979; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12008 = 3'h4 == state ? ram_0_62 : _GEN_10980; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12009 = 3'h4 == state ? ram_0_63 : _GEN_10981; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12010 = 3'h4 == state ? ram_0_64 : _GEN_10982; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12011 = 3'h4 == state ? ram_0_65 : _GEN_10983; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12012 = 3'h4 == state ? ram_0_66 : _GEN_10984; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12013 = 3'h4 == state ? ram_0_67 : _GEN_10985; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12014 = 3'h4 == state ? ram_0_68 : _GEN_10986; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12015 = 3'h4 == state ? ram_0_69 : _GEN_10987; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12016 = 3'h4 == state ? ram_0_70 : _GEN_10988; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12017 = 3'h4 == state ? ram_0_71 : _GEN_10989; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12018 = 3'h4 == state ? ram_0_72 : _GEN_10990; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12019 = 3'h4 == state ? ram_0_73 : _GEN_10991; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12020 = 3'h4 == state ? ram_0_74 : _GEN_10992; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12021 = 3'h4 == state ? ram_0_75 : _GEN_10993; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12022 = 3'h4 == state ? ram_0_76 : _GEN_10994; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12023 = 3'h4 == state ? ram_0_77 : _GEN_10995; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12024 = 3'h4 == state ? ram_0_78 : _GEN_10996; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12025 = 3'h4 == state ? ram_0_79 : _GEN_10997; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12026 = 3'h4 == state ? ram_0_80 : _GEN_10998; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12027 = 3'h4 == state ? ram_0_81 : _GEN_10999; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12028 = 3'h4 == state ? ram_0_82 : _GEN_11000; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12029 = 3'h4 == state ? ram_0_83 : _GEN_11001; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12030 = 3'h4 == state ? ram_0_84 : _GEN_11002; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12031 = 3'h4 == state ? ram_0_85 : _GEN_11003; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12032 = 3'h4 == state ? ram_0_86 : _GEN_11004; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12033 = 3'h4 == state ? ram_0_87 : _GEN_11005; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12034 = 3'h4 == state ? ram_0_88 : _GEN_11006; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12035 = 3'h4 == state ? ram_0_89 : _GEN_11007; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12036 = 3'h4 == state ? ram_0_90 : _GEN_11008; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12037 = 3'h4 == state ? ram_0_91 : _GEN_11009; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12038 = 3'h4 == state ? ram_0_92 : _GEN_11010; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12039 = 3'h4 == state ? ram_0_93 : _GEN_11011; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12040 = 3'h4 == state ? ram_0_94 : _GEN_11012; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12041 = 3'h4 == state ? ram_0_95 : _GEN_11013; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12042 = 3'h4 == state ? ram_0_96 : _GEN_11014; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12043 = 3'h4 == state ? ram_0_97 : _GEN_11015; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12044 = 3'h4 == state ? ram_0_98 : _GEN_11016; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12045 = 3'h4 == state ? ram_0_99 : _GEN_11017; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12046 = 3'h4 == state ? ram_0_100 : _GEN_11018; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12047 = 3'h4 == state ? ram_0_101 : _GEN_11019; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12048 = 3'h4 == state ? ram_0_102 : _GEN_11020; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12049 = 3'h4 == state ? ram_0_103 : _GEN_11021; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12050 = 3'h4 == state ? ram_0_104 : _GEN_11022; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12051 = 3'h4 == state ? ram_0_105 : _GEN_11023; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12052 = 3'h4 == state ? ram_0_106 : _GEN_11024; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12053 = 3'h4 == state ? ram_0_107 : _GEN_11025; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12054 = 3'h4 == state ? ram_0_108 : _GEN_11026; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12055 = 3'h4 == state ? ram_0_109 : _GEN_11027; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12056 = 3'h4 == state ? ram_0_110 : _GEN_11028; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12057 = 3'h4 == state ? ram_0_111 : _GEN_11029; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12058 = 3'h4 == state ? ram_0_112 : _GEN_11030; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12059 = 3'h4 == state ? ram_0_113 : _GEN_11031; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12060 = 3'h4 == state ? ram_0_114 : _GEN_11032; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12061 = 3'h4 == state ? ram_0_115 : _GEN_11033; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12062 = 3'h4 == state ? ram_0_116 : _GEN_11034; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12063 = 3'h4 == state ? ram_0_117 : _GEN_11035; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12064 = 3'h4 == state ? ram_0_118 : _GEN_11036; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12065 = 3'h4 == state ? ram_0_119 : _GEN_11037; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12066 = 3'h4 == state ? ram_0_120 : _GEN_11038; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12067 = 3'h4 == state ? ram_0_121 : _GEN_11039; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12068 = 3'h4 == state ? ram_0_122 : _GEN_11040; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12069 = 3'h4 == state ? ram_0_123 : _GEN_11041; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12070 = 3'h4 == state ? ram_0_124 : _GEN_11042; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12071 = 3'h4 == state ? ram_0_125 : _GEN_11043; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12072 = 3'h4 == state ? ram_0_126 : _GEN_11044; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12073 = 3'h4 == state ? ram_0_127 : _GEN_11045; // @[d_cache.scala 87:18 19:24]
  wire [31:0] _GEN_12074 = 3'h4 == state ? tag_0_0 : _GEN_11046; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12075 = 3'h4 == state ? tag_0_1 : _GEN_11047; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12076 = 3'h4 == state ? tag_0_2 : _GEN_11048; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12077 = 3'h4 == state ? tag_0_3 : _GEN_11049; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12078 = 3'h4 == state ? tag_0_4 : _GEN_11050; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12079 = 3'h4 == state ? tag_0_5 : _GEN_11051; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12080 = 3'h4 == state ? tag_0_6 : _GEN_11052; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12081 = 3'h4 == state ? tag_0_7 : _GEN_11053; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12082 = 3'h4 == state ? tag_0_8 : _GEN_11054; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12083 = 3'h4 == state ? tag_0_9 : _GEN_11055; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12084 = 3'h4 == state ? tag_0_10 : _GEN_11056; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12085 = 3'h4 == state ? tag_0_11 : _GEN_11057; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12086 = 3'h4 == state ? tag_0_12 : _GEN_11058; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12087 = 3'h4 == state ? tag_0_13 : _GEN_11059; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12088 = 3'h4 == state ? tag_0_14 : _GEN_11060; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12089 = 3'h4 == state ? tag_0_15 : _GEN_11061; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12090 = 3'h4 == state ? tag_0_16 : _GEN_11062; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12091 = 3'h4 == state ? tag_0_17 : _GEN_11063; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12092 = 3'h4 == state ? tag_0_18 : _GEN_11064; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12093 = 3'h4 == state ? tag_0_19 : _GEN_11065; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12094 = 3'h4 == state ? tag_0_20 : _GEN_11066; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12095 = 3'h4 == state ? tag_0_21 : _GEN_11067; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12096 = 3'h4 == state ? tag_0_22 : _GEN_11068; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12097 = 3'h4 == state ? tag_0_23 : _GEN_11069; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12098 = 3'h4 == state ? tag_0_24 : _GEN_11070; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12099 = 3'h4 == state ? tag_0_25 : _GEN_11071; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12100 = 3'h4 == state ? tag_0_26 : _GEN_11072; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12101 = 3'h4 == state ? tag_0_27 : _GEN_11073; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12102 = 3'h4 == state ? tag_0_28 : _GEN_11074; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12103 = 3'h4 == state ? tag_0_29 : _GEN_11075; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12104 = 3'h4 == state ? tag_0_30 : _GEN_11076; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12105 = 3'h4 == state ? tag_0_31 : _GEN_11077; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12106 = 3'h4 == state ? tag_0_32 : _GEN_11078; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12107 = 3'h4 == state ? tag_0_33 : _GEN_11079; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12108 = 3'h4 == state ? tag_0_34 : _GEN_11080; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12109 = 3'h4 == state ? tag_0_35 : _GEN_11081; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12110 = 3'h4 == state ? tag_0_36 : _GEN_11082; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12111 = 3'h4 == state ? tag_0_37 : _GEN_11083; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12112 = 3'h4 == state ? tag_0_38 : _GEN_11084; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12113 = 3'h4 == state ? tag_0_39 : _GEN_11085; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12114 = 3'h4 == state ? tag_0_40 : _GEN_11086; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12115 = 3'h4 == state ? tag_0_41 : _GEN_11087; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12116 = 3'h4 == state ? tag_0_42 : _GEN_11088; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12117 = 3'h4 == state ? tag_0_43 : _GEN_11089; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12118 = 3'h4 == state ? tag_0_44 : _GEN_11090; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12119 = 3'h4 == state ? tag_0_45 : _GEN_11091; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12120 = 3'h4 == state ? tag_0_46 : _GEN_11092; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12121 = 3'h4 == state ? tag_0_47 : _GEN_11093; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12122 = 3'h4 == state ? tag_0_48 : _GEN_11094; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12123 = 3'h4 == state ? tag_0_49 : _GEN_11095; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12124 = 3'h4 == state ? tag_0_50 : _GEN_11096; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12125 = 3'h4 == state ? tag_0_51 : _GEN_11097; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12126 = 3'h4 == state ? tag_0_52 : _GEN_11098; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12127 = 3'h4 == state ? tag_0_53 : _GEN_11099; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12128 = 3'h4 == state ? tag_0_54 : _GEN_11100; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12129 = 3'h4 == state ? tag_0_55 : _GEN_11101; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12130 = 3'h4 == state ? tag_0_56 : _GEN_11102; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12131 = 3'h4 == state ? tag_0_57 : _GEN_11103; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12132 = 3'h4 == state ? tag_0_58 : _GEN_11104; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12133 = 3'h4 == state ? tag_0_59 : _GEN_11105; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12134 = 3'h4 == state ? tag_0_60 : _GEN_11106; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12135 = 3'h4 == state ? tag_0_61 : _GEN_11107; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12136 = 3'h4 == state ? tag_0_62 : _GEN_11108; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12137 = 3'h4 == state ? tag_0_63 : _GEN_11109; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12138 = 3'h4 == state ? tag_0_64 : _GEN_11110; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12139 = 3'h4 == state ? tag_0_65 : _GEN_11111; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12140 = 3'h4 == state ? tag_0_66 : _GEN_11112; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12141 = 3'h4 == state ? tag_0_67 : _GEN_11113; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12142 = 3'h4 == state ? tag_0_68 : _GEN_11114; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12143 = 3'h4 == state ? tag_0_69 : _GEN_11115; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12144 = 3'h4 == state ? tag_0_70 : _GEN_11116; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12145 = 3'h4 == state ? tag_0_71 : _GEN_11117; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12146 = 3'h4 == state ? tag_0_72 : _GEN_11118; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12147 = 3'h4 == state ? tag_0_73 : _GEN_11119; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12148 = 3'h4 == state ? tag_0_74 : _GEN_11120; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12149 = 3'h4 == state ? tag_0_75 : _GEN_11121; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12150 = 3'h4 == state ? tag_0_76 : _GEN_11122; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12151 = 3'h4 == state ? tag_0_77 : _GEN_11123; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12152 = 3'h4 == state ? tag_0_78 : _GEN_11124; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12153 = 3'h4 == state ? tag_0_79 : _GEN_11125; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12154 = 3'h4 == state ? tag_0_80 : _GEN_11126; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12155 = 3'h4 == state ? tag_0_81 : _GEN_11127; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12156 = 3'h4 == state ? tag_0_82 : _GEN_11128; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12157 = 3'h4 == state ? tag_0_83 : _GEN_11129; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12158 = 3'h4 == state ? tag_0_84 : _GEN_11130; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12159 = 3'h4 == state ? tag_0_85 : _GEN_11131; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12160 = 3'h4 == state ? tag_0_86 : _GEN_11132; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12161 = 3'h4 == state ? tag_0_87 : _GEN_11133; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12162 = 3'h4 == state ? tag_0_88 : _GEN_11134; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12163 = 3'h4 == state ? tag_0_89 : _GEN_11135; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12164 = 3'h4 == state ? tag_0_90 : _GEN_11136; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12165 = 3'h4 == state ? tag_0_91 : _GEN_11137; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12166 = 3'h4 == state ? tag_0_92 : _GEN_11138; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12167 = 3'h4 == state ? tag_0_93 : _GEN_11139; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12168 = 3'h4 == state ? tag_0_94 : _GEN_11140; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12169 = 3'h4 == state ? tag_0_95 : _GEN_11141; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12170 = 3'h4 == state ? tag_0_96 : _GEN_11142; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12171 = 3'h4 == state ? tag_0_97 : _GEN_11143; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12172 = 3'h4 == state ? tag_0_98 : _GEN_11144; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12173 = 3'h4 == state ? tag_0_99 : _GEN_11145; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12174 = 3'h4 == state ? tag_0_100 : _GEN_11146; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12175 = 3'h4 == state ? tag_0_101 : _GEN_11147; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12176 = 3'h4 == state ? tag_0_102 : _GEN_11148; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12177 = 3'h4 == state ? tag_0_103 : _GEN_11149; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12178 = 3'h4 == state ? tag_0_104 : _GEN_11150; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12179 = 3'h4 == state ? tag_0_105 : _GEN_11151; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12180 = 3'h4 == state ? tag_0_106 : _GEN_11152; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12181 = 3'h4 == state ? tag_0_107 : _GEN_11153; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12182 = 3'h4 == state ? tag_0_108 : _GEN_11154; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12183 = 3'h4 == state ? tag_0_109 : _GEN_11155; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12184 = 3'h4 == state ? tag_0_110 : _GEN_11156; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12185 = 3'h4 == state ? tag_0_111 : _GEN_11157; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12186 = 3'h4 == state ? tag_0_112 : _GEN_11158; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12187 = 3'h4 == state ? tag_0_113 : _GEN_11159; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12188 = 3'h4 == state ? tag_0_114 : _GEN_11160; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12189 = 3'h4 == state ? tag_0_115 : _GEN_11161; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12190 = 3'h4 == state ? tag_0_116 : _GEN_11162; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12191 = 3'h4 == state ? tag_0_117 : _GEN_11163; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12192 = 3'h4 == state ? tag_0_118 : _GEN_11164; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12193 = 3'h4 == state ? tag_0_119 : _GEN_11165; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12194 = 3'h4 == state ? tag_0_120 : _GEN_11166; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12195 = 3'h4 == state ? tag_0_121 : _GEN_11167; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12196 = 3'h4 == state ? tag_0_122 : _GEN_11168; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12197 = 3'h4 == state ? tag_0_123 : _GEN_11169; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12198 = 3'h4 == state ? tag_0_124 : _GEN_11170; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12199 = 3'h4 == state ? tag_0_125 : _GEN_11171; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12200 = 3'h4 == state ? tag_0_126 : _GEN_11172; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_12201 = 3'h4 == state ? tag_0_127 : _GEN_11173; // @[d_cache.scala 87:18 28:24]
  wire  _GEN_12202 = 3'h4 == state ? valid_0_0 : _GEN_11174; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12203 = 3'h4 == state ? valid_0_1 : _GEN_11175; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12204 = 3'h4 == state ? valid_0_2 : _GEN_11176; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12205 = 3'h4 == state ? valid_0_3 : _GEN_11177; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12206 = 3'h4 == state ? valid_0_4 : _GEN_11178; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12207 = 3'h4 == state ? valid_0_5 : _GEN_11179; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12208 = 3'h4 == state ? valid_0_6 : _GEN_11180; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12209 = 3'h4 == state ? valid_0_7 : _GEN_11181; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12210 = 3'h4 == state ? valid_0_8 : _GEN_11182; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12211 = 3'h4 == state ? valid_0_9 : _GEN_11183; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12212 = 3'h4 == state ? valid_0_10 : _GEN_11184; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12213 = 3'h4 == state ? valid_0_11 : _GEN_11185; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12214 = 3'h4 == state ? valid_0_12 : _GEN_11186; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12215 = 3'h4 == state ? valid_0_13 : _GEN_11187; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12216 = 3'h4 == state ? valid_0_14 : _GEN_11188; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12217 = 3'h4 == state ? valid_0_15 : _GEN_11189; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12218 = 3'h4 == state ? valid_0_16 : _GEN_11190; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12219 = 3'h4 == state ? valid_0_17 : _GEN_11191; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12220 = 3'h4 == state ? valid_0_18 : _GEN_11192; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12221 = 3'h4 == state ? valid_0_19 : _GEN_11193; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12222 = 3'h4 == state ? valid_0_20 : _GEN_11194; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12223 = 3'h4 == state ? valid_0_21 : _GEN_11195; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12224 = 3'h4 == state ? valid_0_22 : _GEN_11196; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12225 = 3'h4 == state ? valid_0_23 : _GEN_11197; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12226 = 3'h4 == state ? valid_0_24 : _GEN_11198; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12227 = 3'h4 == state ? valid_0_25 : _GEN_11199; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12228 = 3'h4 == state ? valid_0_26 : _GEN_11200; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12229 = 3'h4 == state ? valid_0_27 : _GEN_11201; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12230 = 3'h4 == state ? valid_0_28 : _GEN_11202; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12231 = 3'h4 == state ? valid_0_29 : _GEN_11203; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12232 = 3'h4 == state ? valid_0_30 : _GEN_11204; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12233 = 3'h4 == state ? valid_0_31 : _GEN_11205; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12234 = 3'h4 == state ? valid_0_32 : _GEN_11206; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12235 = 3'h4 == state ? valid_0_33 : _GEN_11207; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12236 = 3'h4 == state ? valid_0_34 : _GEN_11208; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12237 = 3'h4 == state ? valid_0_35 : _GEN_11209; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12238 = 3'h4 == state ? valid_0_36 : _GEN_11210; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12239 = 3'h4 == state ? valid_0_37 : _GEN_11211; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12240 = 3'h4 == state ? valid_0_38 : _GEN_11212; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12241 = 3'h4 == state ? valid_0_39 : _GEN_11213; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12242 = 3'h4 == state ? valid_0_40 : _GEN_11214; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12243 = 3'h4 == state ? valid_0_41 : _GEN_11215; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12244 = 3'h4 == state ? valid_0_42 : _GEN_11216; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12245 = 3'h4 == state ? valid_0_43 : _GEN_11217; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12246 = 3'h4 == state ? valid_0_44 : _GEN_11218; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12247 = 3'h4 == state ? valid_0_45 : _GEN_11219; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12248 = 3'h4 == state ? valid_0_46 : _GEN_11220; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12249 = 3'h4 == state ? valid_0_47 : _GEN_11221; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12250 = 3'h4 == state ? valid_0_48 : _GEN_11222; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12251 = 3'h4 == state ? valid_0_49 : _GEN_11223; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12252 = 3'h4 == state ? valid_0_50 : _GEN_11224; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12253 = 3'h4 == state ? valid_0_51 : _GEN_11225; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12254 = 3'h4 == state ? valid_0_52 : _GEN_11226; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12255 = 3'h4 == state ? valid_0_53 : _GEN_11227; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12256 = 3'h4 == state ? valid_0_54 : _GEN_11228; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12257 = 3'h4 == state ? valid_0_55 : _GEN_11229; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12258 = 3'h4 == state ? valid_0_56 : _GEN_11230; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12259 = 3'h4 == state ? valid_0_57 : _GEN_11231; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12260 = 3'h4 == state ? valid_0_58 : _GEN_11232; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12261 = 3'h4 == state ? valid_0_59 : _GEN_11233; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12262 = 3'h4 == state ? valid_0_60 : _GEN_11234; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12263 = 3'h4 == state ? valid_0_61 : _GEN_11235; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12264 = 3'h4 == state ? valid_0_62 : _GEN_11236; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12265 = 3'h4 == state ? valid_0_63 : _GEN_11237; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12266 = 3'h4 == state ? valid_0_64 : _GEN_11238; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12267 = 3'h4 == state ? valid_0_65 : _GEN_11239; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12268 = 3'h4 == state ? valid_0_66 : _GEN_11240; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12269 = 3'h4 == state ? valid_0_67 : _GEN_11241; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12270 = 3'h4 == state ? valid_0_68 : _GEN_11242; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12271 = 3'h4 == state ? valid_0_69 : _GEN_11243; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12272 = 3'h4 == state ? valid_0_70 : _GEN_11244; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12273 = 3'h4 == state ? valid_0_71 : _GEN_11245; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12274 = 3'h4 == state ? valid_0_72 : _GEN_11246; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12275 = 3'h4 == state ? valid_0_73 : _GEN_11247; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12276 = 3'h4 == state ? valid_0_74 : _GEN_11248; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12277 = 3'h4 == state ? valid_0_75 : _GEN_11249; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12278 = 3'h4 == state ? valid_0_76 : _GEN_11250; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12279 = 3'h4 == state ? valid_0_77 : _GEN_11251; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12280 = 3'h4 == state ? valid_0_78 : _GEN_11252; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12281 = 3'h4 == state ? valid_0_79 : _GEN_11253; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12282 = 3'h4 == state ? valid_0_80 : _GEN_11254; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12283 = 3'h4 == state ? valid_0_81 : _GEN_11255; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12284 = 3'h4 == state ? valid_0_82 : _GEN_11256; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12285 = 3'h4 == state ? valid_0_83 : _GEN_11257; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12286 = 3'h4 == state ? valid_0_84 : _GEN_11258; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12287 = 3'h4 == state ? valid_0_85 : _GEN_11259; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12288 = 3'h4 == state ? valid_0_86 : _GEN_11260; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12289 = 3'h4 == state ? valid_0_87 : _GEN_11261; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12290 = 3'h4 == state ? valid_0_88 : _GEN_11262; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12291 = 3'h4 == state ? valid_0_89 : _GEN_11263; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12292 = 3'h4 == state ? valid_0_90 : _GEN_11264; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12293 = 3'h4 == state ? valid_0_91 : _GEN_11265; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12294 = 3'h4 == state ? valid_0_92 : _GEN_11266; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12295 = 3'h4 == state ? valid_0_93 : _GEN_11267; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12296 = 3'h4 == state ? valid_0_94 : _GEN_11268; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12297 = 3'h4 == state ? valid_0_95 : _GEN_11269; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12298 = 3'h4 == state ? valid_0_96 : _GEN_11270; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12299 = 3'h4 == state ? valid_0_97 : _GEN_11271; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12300 = 3'h4 == state ? valid_0_98 : _GEN_11272; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12301 = 3'h4 == state ? valid_0_99 : _GEN_11273; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12302 = 3'h4 == state ? valid_0_100 : _GEN_11274; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12303 = 3'h4 == state ? valid_0_101 : _GEN_11275; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12304 = 3'h4 == state ? valid_0_102 : _GEN_11276; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12305 = 3'h4 == state ? valid_0_103 : _GEN_11277; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12306 = 3'h4 == state ? valid_0_104 : _GEN_11278; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12307 = 3'h4 == state ? valid_0_105 : _GEN_11279; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12308 = 3'h4 == state ? valid_0_106 : _GEN_11280; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12309 = 3'h4 == state ? valid_0_107 : _GEN_11281; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12310 = 3'h4 == state ? valid_0_108 : _GEN_11282; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12311 = 3'h4 == state ? valid_0_109 : _GEN_11283; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12312 = 3'h4 == state ? valid_0_110 : _GEN_11284; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12313 = 3'h4 == state ? valid_0_111 : _GEN_11285; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12314 = 3'h4 == state ? valid_0_112 : _GEN_11286; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12315 = 3'h4 == state ? valid_0_113 : _GEN_11287; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12316 = 3'h4 == state ? valid_0_114 : _GEN_11288; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12317 = 3'h4 == state ? valid_0_115 : _GEN_11289; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12318 = 3'h4 == state ? valid_0_116 : _GEN_11290; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12319 = 3'h4 == state ? valid_0_117 : _GEN_11291; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12320 = 3'h4 == state ? valid_0_118 : _GEN_11292; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12321 = 3'h4 == state ? valid_0_119 : _GEN_11293; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12322 = 3'h4 == state ? valid_0_120 : _GEN_11294; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12323 = 3'h4 == state ? valid_0_121 : _GEN_11295; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12324 = 3'h4 == state ? valid_0_122 : _GEN_11296; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12325 = 3'h4 == state ? valid_0_123 : _GEN_11297; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12326 = 3'h4 == state ? valid_0_124 : _GEN_11298; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12327 = 3'h4 == state ? valid_0_125 : _GEN_11299; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12328 = 3'h4 == state ? valid_0_126 : _GEN_11300; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12329 = 3'h4 == state ? valid_0_127 : _GEN_11301; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_12330 = 3'h4 == state ? quene : _GEN_11302; // @[d_cache.scala 87:18 43:24]
  wire [63:0] _GEN_12331 = 3'h4 == state ? ram_1_0 : _GEN_11303; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12332 = 3'h4 == state ? ram_1_1 : _GEN_11304; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12333 = 3'h4 == state ? ram_1_2 : _GEN_11305; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12334 = 3'h4 == state ? ram_1_3 : _GEN_11306; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12335 = 3'h4 == state ? ram_1_4 : _GEN_11307; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12336 = 3'h4 == state ? ram_1_5 : _GEN_11308; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12337 = 3'h4 == state ? ram_1_6 : _GEN_11309; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12338 = 3'h4 == state ? ram_1_7 : _GEN_11310; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12339 = 3'h4 == state ? ram_1_8 : _GEN_11311; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12340 = 3'h4 == state ? ram_1_9 : _GEN_11312; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12341 = 3'h4 == state ? ram_1_10 : _GEN_11313; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12342 = 3'h4 == state ? ram_1_11 : _GEN_11314; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12343 = 3'h4 == state ? ram_1_12 : _GEN_11315; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12344 = 3'h4 == state ? ram_1_13 : _GEN_11316; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12345 = 3'h4 == state ? ram_1_14 : _GEN_11317; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12346 = 3'h4 == state ? ram_1_15 : _GEN_11318; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12347 = 3'h4 == state ? ram_1_16 : _GEN_11319; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12348 = 3'h4 == state ? ram_1_17 : _GEN_11320; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12349 = 3'h4 == state ? ram_1_18 : _GEN_11321; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12350 = 3'h4 == state ? ram_1_19 : _GEN_11322; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12351 = 3'h4 == state ? ram_1_20 : _GEN_11323; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12352 = 3'h4 == state ? ram_1_21 : _GEN_11324; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12353 = 3'h4 == state ? ram_1_22 : _GEN_11325; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12354 = 3'h4 == state ? ram_1_23 : _GEN_11326; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12355 = 3'h4 == state ? ram_1_24 : _GEN_11327; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12356 = 3'h4 == state ? ram_1_25 : _GEN_11328; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12357 = 3'h4 == state ? ram_1_26 : _GEN_11329; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12358 = 3'h4 == state ? ram_1_27 : _GEN_11330; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12359 = 3'h4 == state ? ram_1_28 : _GEN_11331; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12360 = 3'h4 == state ? ram_1_29 : _GEN_11332; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12361 = 3'h4 == state ? ram_1_30 : _GEN_11333; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12362 = 3'h4 == state ? ram_1_31 : _GEN_11334; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12363 = 3'h4 == state ? ram_1_32 : _GEN_11335; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12364 = 3'h4 == state ? ram_1_33 : _GEN_11336; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12365 = 3'h4 == state ? ram_1_34 : _GEN_11337; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12366 = 3'h4 == state ? ram_1_35 : _GEN_11338; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12367 = 3'h4 == state ? ram_1_36 : _GEN_11339; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12368 = 3'h4 == state ? ram_1_37 : _GEN_11340; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12369 = 3'h4 == state ? ram_1_38 : _GEN_11341; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12370 = 3'h4 == state ? ram_1_39 : _GEN_11342; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12371 = 3'h4 == state ? ram_1_40 : _GEN_11343; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12372 = 3'h4 == state ? ram_1_41 : _GEN_11344; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12373 = 3'h4 == state ? ram_1_42 : _GEN_11345; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12374 = 3'h4 == state ? ram_1_43 : _GEN_11346; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12375 = 3'h4 == state ? ram_1_44 : _GEN_11347; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12376 = 3'h4 == state ? ram_1_45 : _GEN_11348; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12377 = 3'h4 == state ? ram_1_46 : _GEN_11349; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12378 = 3'h4 == state ? ram_1_47 : _GEN_11350; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12379 = 3'h4 == state ? ram_1_48 : _GEN_11351; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12380 = 3'h4 == state ? ram_1_49 : _GEN_11352; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12381 = 3'h4 == state ? ram_1_50 : _GEN_11353; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12382 = 3'h4 == state ? ram_1_51 : _GEN_11354; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12383 = 3'h4 == state ? ram_1_52 : _GEN_11355; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12384 = 3'h4 == state ? ram_1_53 : _GEN_11356; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12385 = 3'h4 == state ? ram_1_54 : _GEN_11357; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12386 = 3'h4 == state ? ram_1_55 : _GEN_11358; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12387 = 3'h4 == state ? ram_1_56 : _GEN_11359; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12388 = 3'h4 == state ? ram_1_57 : _GEN_11360; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12389 = 3'h4 == state ? ram_1_58 : _GEN_11361; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12390 = 3'h4 == state ? ram_1_59 : _GEN_11362; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12391 = 3'h4 == state ? ram_1_60 : _GEN_11363; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12392 = 3'h4 == state ? ram_1_61 : _GEN_11364; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12393 = 3'h4 == state ? ram_1_62 : _GEN_11365; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12394 = 3'h4 == state ? ram_1_63 : _GEN_11366; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12395 = 3'h4 == state ? ram_1_64 : _GEN_11367; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12396 = 3'h4 == state ? ram_1_65 : _GEN_11368; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12397 = 3'h4 == state ? ram_1_66 : _GEN_11369; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12398 = 3'h4 == state ? ram_1_67 : _GEN_11370; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12399 = 3'h4 == state ? ram_1_68 : _GEN_11371; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12400 = 3'h4 == state ? ram_1_69 : _GEN_11372; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12401 = 3'h4 == state ? ram_1_70 : _GEN_11373; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12402 = 3'h4 == state ? ram_1_71 : _GEN_11374; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12403 = 3'h4 == state ? ram_1_72 : _GEN_11375; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12404 = 3'h4 == state ? ram_1_73 : _GEN_11376; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12405 = 3'h4 == state ? ram_1_74 : _GEN_11377; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12406 = 3'h4 == state ? ram_1_75 : _GEN_11378; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12407 = 3'h4 == state ? ram_1_76 : _GEN_11379; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12408 = 3'h4 == state ? ram_1_77 : _GEN_11380; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12409 = 3'h4 == state ? ram_1_78 : _GEN_11381; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12410 = 3'h4 == state ? ram_1_79 : _GEN_11382; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12411 = 3'h4 == state ? ram_1_80 : _GEN_11383; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12412 = 3'h4 == state ? ram_1_81 : _GEN_11384; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12413 = 3'h4 == state ? ram_1_82 : _GEN_11385; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12414 = 3'h4 == state ? ram_1_83 : _GEN_11386; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12415 = 3'h4 == state ? ram_1_84 : _GEN_11387; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12416 = 3'h4 == state ? ram_1_85 : _GEN_11388; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12417 = 3'h4 == state ? ram_1_86 : _GEN_11389; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12418 = 3'h4 == state ? ram_1_87 : _GEN_11390; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12419 = 3'h4 == state ? ram_1_88 : _GEN_11391; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12420 = 3'h4 == state ? ram_1_89 : _GEN_11392; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12421 = 3'h4 == state ? ram_1_90 : _GEN_11393; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12422 = 3'h4 == state ? ram_1_91 : _GEN_11394; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12423 = 3'h4 == state ? ram_1_92 : _GEN_11395; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12424 = 3'h4 == state ? ram_1_93 : _GEN_11396; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12425 = 3'h4 == state ? ram_1_94 : _GEN_11397; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12426 = 3'h4 == state ? ram_1_95 : _GEN_11398; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12427 = 3'h4 == state ? ram_1_96 : _GEN_11399; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12428 = 3'h4 == state ? ram_1_97 : _GEN_11400; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12429 = 3'h4 == state ? ram_1_98 : _GEN_11401; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12430 = 3'h4 == state ? ram_1_99 : _GEN_11402; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12431 = 3'h4 == state ? ram_1_100 : _GEN_11403; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12432 = 3'h4 == state ? ram_1_101 : _GEN_11404; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12433 = 3'h4 == state ? ram_1_102 : _GEN_11405; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12434 = 3'h4 == state ? ram_1_103 : _GEN_11406; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12435 = 3'h4 == state ? ram_1_104 : _GEN_11407; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12436 = 3'h4 == state ? ram_1_105 : _GEN_11408; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12437 = 3'h4 == state ? ram_1_106 : _GEN_11409; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12438 = 3'h4 == state ? ram_1_107 : _GEN_11410; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12439 = 3'h4 == state ? ram_1_108 : _GEN_11411; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12440 = 3'h4 == state ? ram_1_109 : _GEN_11412; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12441 = 3'h4 == state ? ram_1_110 : _GEN_11413; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12442 = 3'h4 == state ? ram_1_111 : _GEN_11414; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12443 = 3'h4 == state ? ram_1_112 : _GEN_11415; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12444 = 3'h4 == state ? ram_1_113 : _GEN_11416; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12445 = 3'h4 == state ? ram_1_114 : _GEN_11417; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12446 = 3'h4 == state ? ram_1_115 : _GEN_11418; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12447 = 3'h4 == state ? ram_1_116 : _GEN_11419; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12448 = 3'h4 == state ? ram_1_117 : _GEN_11420; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12449 = 3'h4 == state ? ram_1_118 : _GEN_11421; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12450 = 3'h4 == state ? ram_1_119 : _GEN_11422; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12451 = 3'h4 == state ? ram_1_120 : _GEN_11423; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12452 = 3'h4 == state ? ram_1_121 : _GEN_11424; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12453 = 3'h4 == state ? ram_1_122 : _GEN_11425; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12454 = 3'h4 == state ? ram_1_123 : _GEN_11426; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12455 = 3'h4 == state ? ram_1_124 : _GEN_11427; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12456 = 3'h4 == state ? ram_1_125 : _GEN_11428; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12457 = 3'h4 == state ? ram_1_126 : _GEN_11429; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_12458 = 3'h4 == state ? ram_1_127 : _GEN_11430; // @[d_cache.scala 87:18 20:24]
  wire [31:0] _GEN_12459 = 3'h4 == state ? tag_1_0 : _GEN_11431; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12460 = 3'h4 == state ? tag_1_1 : _GEN_11432; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12461 = 3'h4 == state ? tag_1_2 : _GEN_11433; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12462 = 3'h4 == state ? tag_1_3 : _GEN_11434; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12463 = 3'h4 == state ? tag_1_4 : _GEN_11435; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12464 = 3'h4 == state ? tag_1_5 : _GEN_11436; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12465 = 3'h4 == state ? tag_1_6 : _GEN_11437; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12466 = 3'h4 == state ? tag_1_7 : _GEN_11438; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12467 = 3'h4 == state ? tag_1_8 : _GEN_11439; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12468 = 3'h4 == state ? tag_1_9 : _GEN_11440; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12469 = 3'h4 == state ? tag_1_10 : _GEN_11441; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12470 = 3'h4 == state ? tag_1_11 : _GEN_11442; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12471 = 3'h4 == state ? tag_1_12 : _GEN_11443; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12472 = 3'h4 == state ? tag_1_13 : _GEN_11444; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12473 = 3'h4 == state ? tag_1_14 : _GEN_11445; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12474 = 3'h4 == state ? tag_1_15 : _GEN_11446; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12475 = 3'h4 == state ? tag_1_16 : _GEN_11447; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12476 = 3'h4 == state ? tag_1_17 : _GEN_11448; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12477 = 3'h4 == state ? tag_1_18 : _GEN_11449; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12478 = 3'h4 == state ? tag_1_19 : _GEN_11450; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12479 = 3'h4 == state ? tag_1_20 : _GEN_11451; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12480 = 3'h4 == state ? tag_1_21 : _GEN_11452; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12481 = 3'h4 == state ? tag_1_22 : _GEN_11453; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12482 = 3'h4 == state ? tag_1_23 : _GEN_11454; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12483 = 3'h4 == state ? tag_1_24 : _GEN_11455; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12484 = 3'h4 == state ? tag_1_25 : _GEN_11456; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12485 = 3'h4 == state ? tag_1_26 : _GEN_11457; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12486 = 3'h4 == state ? tag_1_27 : _GEN_11458; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12487 = 3'h4 == state ? tag_1_28 : _GEN_11459; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12488 = 3'h4 == state ? tag_1_29 : _GEN_11460; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12489 = 3'h4 == state ? tag_1_30 : _GEN_11461; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12490 = 3'h4 == state ? tag_1_31 : _GEN_11462; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12491 = 3'h4 == state ? tag_1_32 : _GEN_11463; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12492 = 3'h4 == state ? tag_1_33 : _GEN_11464; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12493 = 3'h4 == state ? tag_1_34 : _GEN_11465; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12494 = 3'h4 == state ? tag_1_35 : _GEN_11466; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12495 = 3'h4 == state ? tag_1_36 : _GEN_11467; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12496 = 3'h4 == state ? tag_1_37 : _GEN_11468; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12497 = 3'h4 == state ? tag_1_38 : _GEN_11469; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12498 = 3'h4 == state ? tag_1_39 : _GEN_11470; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12499 = 3'h4 == state ? tag_1_40 : _GEN_11471; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12500 = 3'h4 == state ? tag_1_41 : _GEN_11472; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12501 = 3'h4 == state ? tag_1_42 : _GEN_11473; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12502 = 3'h4 == state ? tag_1_43 : _GEN_11474; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12503 = 3'h4 == state ? tag_1_44 : _GEN_11475; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12504 = 3'h4 == state ? tag_1_45 : _GEN_11476; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12505 = 3'h4 == state ? tag_1_46 : _GEN_11477; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12506 = 3'h4 == state ? tag_1_47 : _GEN_11478; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12507 = 3'h4 == state ? tag_1_48 : _GEN_11479; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12508 = 3'h4 == state ? tag_1_49 : _GEN_11480; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12509 = 3'h4 == state ? tag_1_50 : _GEN_11481; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12510 = 3'h4 == state ? tag_1_51 : _GEN_11482; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12511 = 3'h4 == state ? tag_1_52 : _GEN_11483; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12512 = 3'h4 == state ? tag_1_53 : _GEN_11484; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12513 = 3'h4 == state ? tag_1_54 : _GEN_11485; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12514 = 3'h4 == state ? tag_1_55 : _GEN_11486; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12515 = 3'h4 == state ? tag_1_56 : _GEN_11487; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12516 = 3'h4 == state ? tag_1_57 : _GEN_11488; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12517 = 3'h4 == state ? tag_1_58 : _GEN_11489; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12518 = 3'h4 == state ? tag_1_59 : _GEN_11490; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12519 = 3'h4 == state ? tag_1_60 : _GEN_11491; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12520 = 3'h4 == state ? tag_1_61 : _GEN_11492; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12521 = 3'h4 == state ? tag_1_62 : _GEN_11493; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12522 = 3'h4 == state ? tag_1_63 : _GEN_11494; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12523 = 3'h4 == state ? tag_1_64 : _GEN_11495; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12524 = 3'h4 == state ? tag_1_65 : _GEN_11496; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12525 = 3'h4 == state ? tag_1_66 : _GEN_11497; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12526 = 3'h4 == state ? tag_1_67 : _GEN_11498; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12527 = 3'h4 == state ? tag_1_68 : _GEN_11499; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12528 = 3'h4 == state ? tag_1_69 : _GEN_11500; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12529 = 3'h4 == state ? tag_1_70 : _GEN_11501; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12530 = 3'h4 == state ? tag_1_71 : _GEN_11502; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12531 = 3'h4 == state ? tag_1_72 : _GEN_11503; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12532 = 3'h4 == state ? tag_1_73 : _GEN_11504; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12533 = 3'h4 == state ? tag_1_74 : _GEN_11505; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12534 = 3'h4 == state ? tag_1_75 : _GEN_11506; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12535 = 3'h4 == state ? tag_1_76 : _GEN_11507; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12536 = 3'h4 == state ? tag_1_77 : _GEN_11508; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12537 = 3'h4 == state ? tag_1_78 : _GEN_11509; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12538 = 3'h4 == state ? tag_1_79 : _GEN_11510; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12539 = 3'h4 == state ? tag_1_80 : _GEN_11511; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12540 = 3'h4 == state ? tag_1_81 : _GEN_11512; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12541 = 3'h4 == state ? tag_1_82 : _GEN_11513; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12542 = 3'h4 == state ? tag_1_83 : _GEN_11514; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12543 = 3'h4 == state ? tag_1_84 : _GEN_11515; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12544 = 3'h4 == state ? tag_1_85 : _GEN_11516; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12545 = 3'h4 == state ? tag_1_86 : _GEN_11517; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12546 = 3'h4 == state ? tag_1_87 : _GEN_11518; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12547 = 3'h4 == state ? tag_1_88 : _GEN_11519; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12548 = 3'h4 == state ? tag_1_89 : _GEN_11520; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12549 = 3'h4 == state ? tag_1_90 : _GEN_11521; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12550 = 3'h4 == state ? tag_1_91 : _GEN_11522; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12551 = 3'h4 == state ? tag_1_92 : _GEN_11523; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12552 = 3'h4 == state ? tag_1_93 : _GEN_11524; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12553 = 3'h4 == state ? tag_1_94 : _GEN_11525; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12554 = 3'h4 == state ? tag_1_95 : _GEN_11526; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12555 = 3'h4 == state ? tag_1_96 : _GEN_11527; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12556 = 3'h4 == state ? tag_1_97 : _GEN_11528; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12557 = 3'h4 == state ? tag_1_98 : _GEN_11529; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12558 = 3'h4 == state ? tag_1_99 : _GEN_11530; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12559 = 3'h4 == state ? tag_1_100 : _GEN_11531; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12560 = 3'h4 == state ? tag_1_101 : _GEN_11532; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12561 = 3'h4 == state ? tag_1_102 : _GEN_11533; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12562 = 3'h4 == state ? tag_1_103 : _GEN_11534; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12563 = 3'h4 == state ? tag_1_104 : _GEN_11535; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12564 = 3'h4 == state ? tag_1_105 : _GEN_11536; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12565 = 3'h4 == state ? tag_1_106 : _GEN_11537; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12566 = 3'h4 == state ? tag_1_107 : _GEN_11538; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12567 = 3'h4 == state ? tag_1_108 : _GEN_11539; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12568 = 3'h4 == state ? tag_1_109 : _GEN_11540; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12569 = 3'h4 == state ? tag_1_110 : _GEN_11541; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12570 = 3'h4 == state ? tag_1_111 : _GEN_11542; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12571 = 3'h4 == state ? tag_1_112 : _GEN_11543; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12572 = 3'h4 == state ? tag_1_113 : _GEN_11544; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12573 = 3'h4 == state ? tag_1_114 : _GEN_11545; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12574 = 3'h4 == state ? tag_1_115 : _GEN_11546; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12575 = 3'h4 == state ? tag_1_116 : _GEN_11547; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12576 = 3'h4 == state ? tag_1_117 : _GEN_11548; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12577 = 3'h4 == state ? tag_1_118 : _GEN_11549; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12578 = 3'h4 == state ? tag_1_119 : _GEN_11550; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12579 = 3'h4 == state ? tag_1_120 : _GEN_11551; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12580 = 3'h4 == state ? tag_1_121 : _GEN_11552; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12581 = 3'h4 == state ? tag_1_122 : _GEN_11553; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12582 = 3'h4 == state ? tag_1_123 : _GEN_11554; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12583 = 3'h4 == state ? tag_1_124 : _GEN_11555; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12584 = 3'h4 == state ? tag_1_125 : _GEN_11556; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12585 = 3'h4 == state ? tag_1_126 : _GEN_11557; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_12586 = 3'h4 == state ? tag_1_127 : _GEN_11558; // @[d_cache.scala 87:18 29:24]
  wire  _GEN_12587 = 3'h4 == state ? valid_1_0 : _GEN_11559; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12588 = 3'h4 == state ? valid_1_1 : _GEN_11560; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12589 = 3'h4 == state ? valid_1_2 : _GEN_11561; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12590 = 3'h4 == state ? valid_1_3 : _GEN_11562; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12591 = 3'h4 == state ? valid_1_4 : _GEN_11563; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12592 = 3'h4 == state ? valid_1_5 : _GEN_11564; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12593 = 3'h4 == state ? valid_1_6 : _GEN_11565; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12594 = 3'h4 == state ? valid_1_7 : _GEN_11566; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12595 = 3'h4 == state ? valid_1_8 : _GEN_11567; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12596 = 3'h4 == state ? valid_1_9 : _GEN_11568; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12597 = 3'h4 == state ? valid_1_10 : _GEN_11569; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12598 = 3'h4 == state ? valid_1_11 : _GEN_11570; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12599 = 3'h4 == state ? valid_1_12 : _GEN_11571; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12600 = 3'h4 == state ? valid_1_13 : _GEN_11572; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12601 = 3'h4 == state ? valid_1_14 : _GEN_11573; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12602 = 3'h4 == state ? valid_1_15 : _GEN_11574; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12603 = 3'h4 == state ? valid_1_16 : _GEN_11575; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12604 = 3'h4 == state ? valid_1_17 : _GEN_11576; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12605 = 3'h4 == state ? valid_1_18 : _GEN_11577; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12606 = 3'h4 == state ? valid_1_19 : _GEN_11578; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12607 = 3'h4 == state ? valid_1_20 : _GEN_11579; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12608 = 3'h4 == state ? valid_1_21 : _GEN_11580; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12609 = 3'h4 == state ? valid_1_22 : _GEN_11581; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12610 = 3'h4 == state ? valid_1_23 : _GEN_11582; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12611 = 3'h4 == state ? valid_1_24 : _GEN_11583; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12612 = 3'h4 == state ? valid_1_25 : _GEN_11584; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12613 = 3'h4 == state ? valid_1_26 : _GEN_11585; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12614 = 3'h4 == state ? valid_1_27 : _GEN_11586; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12615 = 3'h4 == state ? valid_1_28 : _GEN_11587; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12616 = 3'h4 == state ? valid_1_29 : _GEN_11588; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12617 = 3'h4 == state ? valid_1_30 : _GEN_11589; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12618 = 3'h4 == state ? valid_1_31 : _GEN_11590; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12619 = 3'h4 == state ? valid_1_32 : _GEN_11591; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12620 = 3'h4 == state ? valid_1_33 : _GEN_11592; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12621 = 3'h4 == state ? valid_1_34 : _GEN_11593; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12622 = 3'h4 == state ? valid_1_35 : _GEN_11594; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12623 = 3'h4 == state ? valid_1_36 : _GEN_11595; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12624 = 3'h4 == state ? valid_1_37 : _GEN_11596; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12625 = 3'h4 == state ? valid_1_38 : _GEN_11597; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12626 = 3'h4 == state ? valid_1_39 : _GEN_11598; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12627 = 3'h4 == state ? valid_1_40 : _GEN_11599; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12628 = 3'h4 == state ? valid_1_41 : _GEN_11600; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12629 = 3'h4 == state ? valid_1_42 : _GEN_11601; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12630 = 3'h4 == state ? valid_1_43 : _GEN_11602; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12631 = 3'h4 == state ? valid_1_44 : _GEN_11603; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12632 = 3'h4 == state ? valid_1_45 : _GEN_11604; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12633 = 3'h4 == state ? valid_1_46 : _GEN_11605; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12634 = 3'h4 == state ? valid_1_47 : _GEN_11606; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12635 = 3'h4 == state ? valid_1_48 : _GEN_11607; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12636 = 3'h4 == state ? valid_1_49 : _GEN_11608; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12637 = 3'h4 == state ? valid_1_50 : _GEN_11609; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12638 = 3'h4 == state ? valid_1_51 : _GEN_11610; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12639 = 3'h4 == state ? valid_1_52 : _GEN_11611; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12640 = 3'h4 == state ? valid_1_53 : _GEN_11612; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12641 = 3'h4 == state ? valid_1_54 : _GEN_11613; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12642 = 3'h4 == state ? valid_1_55 : _GEN_11614; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12643 = 3'h4 == state ? valid_1_56 : _GEN_11615; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12644 = 3'h4 == state ? valid_1_57 : _GEN_11616; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12645 = 3'h4 == state ? valid_1_58 : _GEN_11617; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12646 = 3'h4 == state ? valid_1_59 : _GEN_11618; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12647 = 3'h4 == state ? valid_1_60 : _GEN_11619; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12648 = 3'h4 == state ? valid_1_61 : _GEN_11620; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12649 = 3'h4 == state ? valid_1_62 : _GEN_11621; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12650 = 3'h4 == state ? valid_1_63 : _GEN_11622; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12651 = 3'h4 == state ? valid_1_64 : _GEN_11623; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12652 = 3'h4 == state ? valid_1_65 : _GEN_11624; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12653 = 3'h4 == state ? valid_1_66 : _GEN_11625; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12654 = 3'h4 == state ? valid_1_67 : _GEN_11626; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12655 = 3'h4 == state ? valid_1_68 : _GEN_11627; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12656 = 3'h4 == state ? valid_1_69 : _GEN_11628; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12657 = 3'h4 == state ? valid_1_70 : _GEN_11629; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12658 = 3'h4 == state ? valid_1_71 : _GEN_11630; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12659 = 3'h4 == state ? valid_1_72 : _GEN_11631; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12660 = 3'h4 == state ? valid_1_73 : _GEN_11632; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12661 = 3'h4 == state ? valid_1_74 : _GEN_11633; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12662 = 3'h4 == state ? valid_1_75 : _GEN_11634; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12663 = 3'h4 == state ? valid_1_76 : _GEN_11635; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12664 = 3'h4 == state ? valid_1_77 : _GEN_11636; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12665 = 3'h4 == state ? valid_1_78 : _GEN_11637; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12666 = 3'h4 == state ? valid_1_79 : _GEN_11638; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12667 = 3'h4 == state ? valid_1_80 : _GEN_11639; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12668 = 3'h4 == state ? valid_1_81 : _GEN_11640; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12669 = 3'h4 == state ? valid_1_82 : _GEN_11641; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12670 = 3'h4 == state ? valid_1_83 : _GEN_11642; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12671 = 3'h4 == state ? valid_1_84 : _GEN_11643; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12672 = 3'h4 == state ? valid_1_85 : _GEN_11644; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12673 = 3'h4 == state ? valid_1_86 : _GEN_11645; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12674 = 3'h4 == state ? valid_1_87 : _GEN_11646; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12675 = 3'h4 == state ? valid_1_88 : _GEN_11647; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12676 = 3'h4 == state ? valid_1_89 : _GEN_11648; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12677 = 3'h4 == state ? valid_1_90 : _GEN_11649; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12678 = 3'h4 == state ? valid_1_91 : _GEN_11650; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12679 = 3'h4 == state ? valid_1_92 : _GEN_11651; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12680 = 3'h4 == state ? valid_1_93 : _GEN_11652; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12681 = 3'h4 == state ? valid_1_94 : _GEN_11653; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12682 = 3'h4 == state ? valid_1_95 : _GEN_11654; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12683 = 3'h4 == state ? valid_1_96 : _GEN_11655; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12684 = 3'h4 == state ? valid_1_97 : _GEN_11656; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12685 = 3'h4 == state ? valid_1_98 : _GEN_11657; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12686 = 3'h4 == state ? valid_1_99 : _GEN_11658; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12687 = 3'h4 == state ? valid_1_100 : _GEN_11659; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12688 = 3'h4 == state ? valid_1_101 : _GEN_11660; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12689 = 3'h4 == state ? valid_1_102 : _GEN_11661; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12690 = 3'h4 == state ? valid_1_103 : _GEN_11662; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12691 = 3'h4 == state ? valid_1_104 : _GEN_11663; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12692 = 3'h4 == state ? valid_1_105 : _GEN_11664; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12693 = 3'h4 == state ? valid_1_106 : _GEN_11665; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12694 = 3'h4 == state ? valid_1_107 : _GEN_11666; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12695 = 3'h4 == state ? valid_1_108 : _GEN_11667; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12696 = 3'h4 == state ? valid_1_109 : _GEN_11668; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12697 = 3'h4 == state ? valid_1_110 : _GEN_11669; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12698 = 3'h4 == state ? valid_1_111 : _GEN_11670; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12699 = 3'h4 == state ? valid_1_112 : _GEN_11671; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12700 = 3'h4 == state ? valid_1_113 : _GEN_11672; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12701 = 3'h4 == state ? valid_1_114 : _GEN_11673; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12702 = 3'h4 == state ? valid_1_115 : _GEN_11674; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12703 = 3'h4 == state ? valid_1_116 : _GEN_11675; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12704 = 3'h4 == state ? valid_1_117 : _GEN_11676; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12705 = 3'h4 == state ? valid_1_118 : _GEN_11677; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12706 = 3'h4 == state ? valid_1_119 : _GEN_11678; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12707 = 3'h4 == state ? valid_1_120 : _GEN_11679; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12708 = 3'h4 == state ? valid_1_121 : _GEN_11680; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12709 = 3'h4 == state ? valid_1_122 : _GEN_11681; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12710 = 3'h4 == state ? valid_1_123 : _GEN_11682; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12711 = 3'h4 == state ? valid_1_124 : _GEN_11683; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12712 = 3'h4 == state ? valid_1_125 : _GEN_11684; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12713 = 3'h4 == state ? valid_1_126 : _GEN_11685; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_12714 = 3'h4 == state ? valid_1_127 : _GEN_11686; // @[d_cache.scala 87:18 31:26]
  wire [63:0] _GEN_12715 = 3'h4 == state ? write_back_data : _GEN_11687; // @[d_cache.scala 87:18 37:34]
  wire [41:0] _GEN_12716 = 3'h4 == state ? {{10'd0}, write_back_addr} : _GEN_11688; // @[d_cache.scala 87:18 38:34]
  wire  _GEN_12717 = 3'h4 == state ? dirty_0_0 : _GEN_11689; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12718 = 3'h4 == state ? dirty_0_1 : _GEN_11690; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12719 = 3'h4 == state ? dirty_0_2 : _GEN_11691; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12720 = 3'h4 == state ? dirty_0_3 : _GEN_11692; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12721 = 3'h4 == state ? dirty_0_4 : _GEN_11693; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12722 = 3'h4 == state ? dirty_0_5 : _GEN_11694; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12723 = 3'h4 == state ? dirty_0_6 : _GEN_11695; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12724 = 3'h4 == state ? dirty_0_7 : _GEN_11696; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12725 = 3'h4 == state ? dirty_0_8 : _GEN_11697; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12726 = 3'h4 == state ? dirty_0_9 : _GEN_11698; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12727 = 3'h4 == state ? dirty_0_10 : _GEN_11699; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12728 = 3'h4 == state ? dirty_0_11 : _GEN_11700; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12729 = 3'h4 == state ? dirty_0_12 : _GEN_11701; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12730 = 3'h4 == state ? dirty_0_13 : _GEN_11702; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12731 = 3'h4 == state ? dirty_0_14 : _GEN_11703; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12732 = 3'h4 == state ? dirty_0_15 : _GEN_11704; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12733 = 3'h4 == state ? dirty_0_16 : _GEN_11705; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12734 = 3'h4 == state ? dirty_0_17 : _GEN_11706; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12735 = 3'h4 == state ? dirty_0_18 : _GEN_11707; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12736 = 3'h4 == state ? dirty_0_19 : _GEN_11708; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12737 = 3'h4 == state ? dirty_0_20 : _GEN_11709; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12738 = 3'h4 == state ? dirty_0_21 : _GEN_11710; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12739 = 3'h4 == state ? dirty_0_22 : _GEN_11711; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12740 = 3'h4 == state ? dirty_0_23 : _GEN_11712; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12741 = 3'h4 == state ? dirty_0_24 : _GEN_11713; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12742 = 3'h4 == state ? dirty_0_25 : _GEN_11714; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12743 = 3'h4 == state ? dirty_0_26 : _GEN_11715; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12744 = 3'h4 == state ? dirty_0_27 : _GEN_11716; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12745 = 3'h4 == state ? dirty_0_28 : _GEN_11717; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12746 = 3'h4 == state ? dirty_0_29 : _GEN_11718; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12747 = 3'h4 == state ? dirty_0_30 : _GEN_11719; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12748 = 3'h4 == state ? dirty_0_31 : _GEN_11720; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12749 = 3'h4 == state ? dirty_0_32 : _GEN_11721; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12750 = 3'h4 == state ? dirty_0_33 : _GEN_11722; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12751 = 3'h4 == state ? dirty_0_34 : _GEN_11723; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12752 = 3'h4 == state ? dirty_0_35 : _GEN_11724; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12753 = 3'h4 == state ? dirty_0_36 : _GEN_11725; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12754 = 3'h4 == state ? dirty_0_37 : _GEN_11726; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12755 = 3'h4 == state ? dirty_0_38 : _GEN_11727; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12756 = 3'h4 == state ? dirty_0_39 : _GEN_11728; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12757 = 3'h4 == state ? dirty_0_40 : _GEN_11729; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12758 = 3'h4 == state ? dirty_0_41 : _GEN_11730; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12759 = 3'h4 == state ? dirty_0_42 : _GEN_11731; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12760 = 3'h4 == state ? dirty_0_43 : _GEN_11732; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12761 = 3'h4 == state ? dirty_0_44 : _GEN_11733; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12762 = 3'h4 == state ? dirty_0_45 : _GEN_11734; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12763 = 3'h4 == state ? dirty_0_46 : _GEN_11735; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12764 = 3'h4 == state ? dirty_0_47 : _GEN_11736; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12765 = 3'h4 == state ? dirty_0_48 : _GEN_11737; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12766 = 3'h4 == state ? dirty_0_49 : _GEN_11738; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12767 = 3'h4 == state ? dirty_0_50 : _GEN_11739; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12768 = 3'h4 == state ? dirty_0_51 : _GEN_11740; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12769 = 3'h4 == state ? dirty_0_52 : _GEN_11741; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12770 = 3'h4 == state ? dirty_0_53 : _GEN_11742; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12771 = 3'h4 == state ? dirty_0_54 : _GEN_11743; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12772 = 3'h4 == state ? dirty_0_55 : _GEN_11744; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12773 = 3'h4 == state ? dirty_0_56 : _GEN_11745; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12774 = 3'h4 == state ? dirty_0_57 : _GEN_11746; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12775 = 3'h4 == state ? dirty_0_58 : _GEN_11747; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12776 = 3'h4 == state ? dirty_0_59 : _GEN_11748; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12777 = 3'h4 == state ? dirty_0_60 : _GEN_11749; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12778 = 3'h4 == state ? dirty_0_61 : _GEN_11750; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12779 = 3'h4 == state ? dirty_0_62 : _GEN_11751; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12780 = 3'h4 == state ? dirty_0_63 : _GEN_11752; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12781 = 3'h4 == state ? dirty_0_64 : _GEN_11753; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12782 = 3'h4 == state ? dirty_0_65 : _GEN_11754; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12783 = 3'h4 == state ? dirty_0_66 : _GEN_11755; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12784 = 3'h4 == state ? dirty_0_67 : _GEN_11756; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12785 = 3'h4 == state ? dirty_0_68 : _GEN_11757; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12786 = 3'h4 == state ? dirty_0_69 : _GEN_11758; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12787 = 3'h4 == state ? dirty_0_70 : _GEN_11759; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12788 = 3'h4 == state ? dirty_0_71 : _GEN_11760; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12789 = 3'h4 == state ? dirty_0_72 : _GEN_11761; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12790 = 3'h4 == state ? dirty_0_73 : _GEN_11762; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12791 = 3'h4 == state ? dirty_0_74 : _GEN_11763; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12792 = 3'h4 == state ? dirty_0_75 : _GEN_11764; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12793 = 3'h4 == state ? dirty_0_76 : _GEN_11765; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12794 = 3'h4 == state ? dirty_0_77 : _GEN_11766; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12795 = 3'h4 == state ? dirty_0_78 : _GEN_11767; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12796 = 3'h4 == state ? dirty_0_79 : _GEN_11768; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12797 = 3'h4 == state ? dirty_0_80 : _GEN_11769; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12798 = 3'h4 == state ? dirty_0_81 : _GEN_11770; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12799 = 3'h4 == state ? dirty_0_82 : _GEN_11771; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12800 = 3'h4 == state ? dirty_0_83 : _GEN_11772; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12801 = 3'h4 == state ? dirty_0_84 : _GEN_11773; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12802 = 3'h4 == state ? dirty_0_85 : _GEN_11774; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12803 = 3'h4 == state ? dirty_0_86 : _GEN_11775; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12804 = 3'h4 == state ? dirty_0_87 : _GEN_11776; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12805 = 3'h4 == state ? dirty_0_88 : _GEN_11777; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12806 = 3'h4 == state ? dirty_0_89 : _GEN_11778; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12807 = 3'h4 == state ? dirty_0_90 : _GEN_11779; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12808 = 3'h4 == state ? dirty_0_91 : _GEN_11780; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12809 = 3'h4 == state ? dirty_0_92 : _GEN_11781; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12810 = 3'h4 == state ? dirty_0_93 : _GEN_11782; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12811 = 3'h4 == state ? dirty_0_94 : _GEN_11783; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12812 = 3'h4 == state ? dirty_0_95 : _GEN_11784; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12813 = 3'h4 == state ? dirty_0_96 : _GEN_11785; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12814 = 3'h4 == state ? dirty_0_97 : _GEN_11786; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12815 = 3'h4 == state ? dirty_0_98 : _GEN_11787; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12816 = 3'h4 == state ? dirty_0_99 : _GEN_11788; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12817 = 3'h4 == state ? dirty_0_100 : _GEN_11789; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12818 = 3'h4 == state ? dirty_0_101 : _GEN_11790; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12819 = 3'h4 == state ? dirty_0_102 : _GEN_11791; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12820 = 3'h4 == state ? dirty_0_103 : _GEN_11792; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12821 = 3'h4 == state ? dirty_0_104 : _GEN_11793; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12822 = 3'h4 == state ? dirty_0_105 : _GEN_11794; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12823 = 3'h4 == state ? dirty_0_106 : _GEN_11795; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12824 = 3'h4 == state ? dirty_0_107 : _GEN_11796; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12825 = 3'h4 == state ? dirty_0_108 : _GEN_11797; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12826 = 3'h4 == state ? dirty_0_109 : _GEN_11798; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12827 = 3'h4 == state ? dirty_0_110 : _GEN_11799; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12828 = 3'h4 == state ? dirty_0_111 : _GEN_11800; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12829 = 3'h4 == state ? dirty_0_112 : _GEN_11801; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12830 = 3'h4 == state ? dirty_0_113 : _GEN_11802; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12831 = 3'h4 == state ? dirty_0_114 : _GEN_11803; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12832 = 3'h4 == state ? dirty_0_115 : _GEN_11804; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12833 = 3'h4 == state ? dirty_0_116 : _GEN_11805; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12834 = 3'h4 == state ? dirty_0_117 : _GEN_11806; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12835 = 3'h4 == state ? dirty_0_118 : _GEN_11807; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12836 = 3'h4 == state ? dirty_0_119 : _GEN_11808; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12837 = 3'h4 == state ? dirty_0_120 : _GEN_11809; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12838 = 3'h4 == state ? dirty_0_121 : _GEN_11810; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12839 = 3'h4 == state ? dirty_0_122 : _GEN_11811; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12840 = 3'h4 == state ? dirty_0_123 : _GEN_11812; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12841 = 3'h4 == state ? dirty_0_124 : _GEN_11813; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12842 = 3'h4 == state ? dirty_0_125 : _GEN_11814; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12843 = 3'h4 == state ? dirty_0_126 : _GEN_11815; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12844 = 3'h4 == state ? dirty_0_127 : _GEN_11816; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_12845 = 3'h4 == state ? dirty_1_0 : _GEN_11817; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12846 = 3'h4 == state ? dirty_1_1 : _GEN_11818; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12847 = 3'h4 == state ? dirty_1_2 : _GEN_11819; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12848 = 3'h4 == state ? dirty_1_3 : _GEN_11820; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12849 = 3'h4 == state ? dirty_1_4 : _GEN_11821; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12850 = 3'h4 == state ? dirty_1_5 : _GEN_11822; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12851 = 3'h4 == state ? dirty_1_6 : _GEN_11823; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12852 = 3'h4 == state ? dirty_1_7 : _GEN_11824; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12853 = 3'h4 == state ? dirty_1_8 : _GEN_11825; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12854 = 3'h4 == state ? dirty_1_9 : _GEN_11826; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12855 = 3'h4 == state ? dirty_1_10 : _GEN_11827; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12856 = 3'h4 == state ? dirty_1_11 : _GEN_11828; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12857 = 3'h4 == state ? dirty_1_12 : _GEN_11829; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12858 = 3'h4 == state ? dirty_1_13 : _GEN_11830; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12859 = 3'h4 == state ? dirty_1_14 : _GEN_11831; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12860 = 3'h4 == state ? dirty_1_15 : _GEN_11832; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12861 = 3'h4 == state ? dirty_1_16 : _GEN_11833; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12862 = 3'h4 == state ? dirty_1_17 : _GEN_11834; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12863 = 3'h4 == state ? dirty_1_18 : _GEN_11835; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12864 = 3'h4 == state ? dirty_1_19 : _GEN_11836; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12865 = 3'h4 == state ? dirty_1_20 : _GEN_11837; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12866 = 3'h4 == state ? dirty_1_21 : _GEN_11838; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12867 = 3'h4 == state ? dirty_1_22 : _GEN_11839; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12868 = 3'h4 == state ? dirty_1_23 : _GEN_11840; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12869 = 3'h4 == state ? dirty_1_24 : _GEN_11841; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12870 = 3'h4 == state ? dirty_1_25 : _GEN_11842; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12871 = 3'h4 == state ? dirty_1_26 : _GEN_11843; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12872 = 3'h4 == state ? dirty_1_27 : _GEN_11844; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12873 = 3'h4 == state ? dirty_1_28 : _GEN_11845; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12874 = 3'h4 == state ? dirty_1_29 : _GEN_11846; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12875 = 3'h4 == state ? dirty_1_30 : _GEN_11847; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12876 = 3'h4 == state ? dirty_1_31 : _GEN_11848; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12877 = 3'h4 == state ? dirty_1_32 : _GEN_11849; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12878 = 3'h4 == state ? dirty_1_33 : _GEN_11850; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12879 = 3'h4 == state ? dirty_1_34 : _GEN_11851; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12880 = 3'h4 == state ? dirty_1_35 : _GEN_11852; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12881 = 3'h4 == state ? dirty_1_36 : _GEN_11853; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12882 = 3'h4 == state ? dirty_1_37 : _GEN_11854; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12883 = 3'h4 == state ? dirty_1_38 : _GEN_11855; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12884 = 3'h4 == state ? dirty_1_39 : _GEN_11856; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12885 = 3'h4 == state ? dirty_1_40 : _GEN_11857; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12886 = 3'h4 == state ? dirty_1_41 : _GEN_11858; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12887 = 3'h4 == state ? dirty_1_42 : _GEN_11859; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12888 = 3'h4 == state ? dirty_1_43 : _GEN_11860; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12889 = 3'h4 == state ? dirty_1_44 : _GEN_11861; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12890 = 3'h4 == state ? dirty_1_45 : _GEN_11862; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12891 = 3'h4 == state ? dirty_1_46 : _GEN_11863; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12892 = 3'h4 == state ? dirty_1_47 : _GEN_11864; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12893 = 3'h4 == state ? dirty_1_48 : _GEN_11865; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12894 = 3'h4 == state ? dirty_1_49 : _GEN_11866; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12895 = 3'h4 == state ? dirty_1_50 : _GEN_11867; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12896 = 3'h4 == state ? dirty_1_51 : _GEN_11868; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12897 = 3'h4 == state ? dirty_1_52 : _GEN_11869; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12898 = 3'h4 == state ? dirty_1_53 : _GEN_11870; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12899 = 3'h4 == state ? dirty_1_54 : _GEN_11871; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12900 = 3'h4 == state ? dirty_1_55 : _GEN_11872; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12901 = 3'h4 == state ? dirty_1_56 : _GEN_11873; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12902 = 3'h4 == state ? dirty_1_57 : _GEN_11874; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12903 = 3'h4 == state ? dirty_1_58 : _GEN_11875; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12904 = 3'h4 == state ? dirty_1_59 : _GEN_11876; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12905 = 3'h4 == state ? dirty_1_60 : _GEN_11877; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12906 = 3'h4 == state ? dirty_1_61 : _GEN_11878; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12907 = 3'h4 == state ? dirty_1_62 : _GEN_11879; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12908 = 3'h4 == state ? dirty_1_63 : _GEN_11880; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12909 = 3'h4 == state ? dirty_1_64 : _GEN_11881; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12910 = 3'h4 == state ? dirty_1_65 : _GEN_11882; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12911 = 3'h4 == state ? dirty_1_66 : _GEN_11883; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12912 = 3'h4 == state ? dirty_1_67 : _GEN_11884; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12913 = 3'h4 == state ? dirty_1_68 : _GEN_11885; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12914 = 3'h4 == state ? dirty_1_69 : _GEN_11886; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12915 = 3'h4 == state ? dirty_1_70 : _GEN_11887; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12916 = 3'h4 == state ? dirty_1_71 : _GEN_11888; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12917 = 3'h4 == state ? dirty_1_72 : _GEN_11889; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12918 = 3'h4 == state ? dirty_1_73 : _GEN_11890; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12919 = 3'h4 == state ? dirty_1_74 : _GEN_11891; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12920 = 3'h4 == state ? dirty_1_75 : _GEN_11892; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12921 = 3'h4 == state ? dirty_1_76 : _GEN_11893; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12922 = 3'h4 == state ? dirty_1_77 : _GEN_11894; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12923 = 3'h4 == state ? dirty_1_78 : _GEN_11895; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12924 = 3'h4 == state ? dirty_1_79 : _GEN_11896; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12925 = 3'h4 == state ? dirty_1_80 : _GEN_11897; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12926 = 3'h4 == state ? dirty_1_81 : _GEN_11898; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12927 = 3'h4 == state ? dirty_1_82 : _GEN_11899; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12928 = 3'h4 == state ? dirty_1_83 : _GEN_11900; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12929 = 3'h4 == state ? dirty_1_84 : _GEN_11901; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12930 = 3'h4 == state ? dirty_1_85 : _GEN_11902; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12931 = 3'h4 == state ? dirty_1_86 : _GEN_11903; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12932 = 3'h4 == state ? dirty_1_87 : _GEN_11904; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12933 = 3'h4 == state ? dirty_1_88 : _GEN_11905; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12934 = 3'h4 == state ? dirty_1_89 : _GEN_11906; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12935 = 3'h4 == state ? dirty_1_90 : _GEN_11907; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12936 = 3'h4 == state ? dirty_1_91 : _GEN_11908; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12937 = 3'h4 == state ? dirty_1_92 : _GEN_11909; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12938 = 3'h4 == state ? dirty_1_93 : _GEN_11910; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12939 = 3'h4 == state ? dirty_1_94 : _GEN_11911; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12940 = 3'h4 == state ? dirty_1_95 : _GEN_11912; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12941 = 3'h4 == state ? dirty_1_96 : _GEN_11913; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12942 = 3'h4 == state ? dirty_1_97 : _GEN_11914; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12943 = 3'h4 == state ? dirty_1_98 : _GEN_11915; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12944 = 3'h4 == state ? dirty_1_99 : _GEN_11916; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12945 = 3'h4 == state ? dirty_1_100 : _GEN_11917; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12946 = 3'h4 == state ? dirty_1_101 : _GEN_11918; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12947 = 3'h4 == state ? dirty_1_102 : _GEN_11919; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12948 = 3'h4 == state ? dirty_1_103 : _GEN_11920; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12949 = 3'h4 == state ? dirty_1_104 : _GEN_11921; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12950 = 3'h4 == state ? dirty_1_105 : _GEN_11922; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12951 = 3'h4 == state ? dirty_1_106 : _GEN_11923; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12952 = 3'h4 == state ? dirty_1_107 : _GEN_11924; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12953 = 3'h4 == state ? dirty_1_108 : _GEN_11925; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12954 = 3'h4 == state ? dirty_1_109 : _GEN_11926; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12955 = 3'h4 == state ? dirty_1_110 : _GEN_11927; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12956 = 3'h4 == state ? dirty_1_111 : _GEN_11928; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12957 = 3'h4 == state ? dirty_1_112 : _GEN_11929; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12958 = 3'h4 == state ? dirty_1_113 : _GEN_11930; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12959 = 3'h4 == state ? dirty_1_114 : _GEN_11931; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12960 = 3'h4 == state ? dirty_1_115 : _GEN_11932; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12961 = 3'h4 == state ? dirty_1_116 : _GEN_11933; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12962 = 3'h4 == state ? dirty_1_117 : _GEN_11934; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12963 = 3'h4 == state ? dirty_1_118 : _GEN_11935; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12964 = 3'h4 == state ? dirty_1_119 : _GEN_11936; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12965 = 3'h4 == state ? dirty_1_120 : _GEN_11937; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12966 = 3'h4 == state ? dirty_1_121 : _GEN_11938; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12967 = 3'h4 == state ? dirty_1_122 : _GEN_11939; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12968 = 3'h4 == state ? dirty_1_123 : _GEN_11940; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12969 = 3'h4 == state ? dirty_1_124 : _GEN_11941; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12970 = 3'h4 == state ? dirty_1_125 : _GEN_11942; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12971 = 3'h4 == state ? dirty_1_126 : _GEN_11943; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_12972 = 3'h4 == state ? dirty_1_127 : _GEN_11944; // @[d_cache.scala 87:18 33:26]
  wire [2:0] _GEN_12973 = 3'h3 == state ? _GEN_4235 : _GEN_11945; // @[d_cache.scala 87:18]
  wire [63:0] _GEN_12974 = 3'h3 == state ? _GEN_4236 : receive_data; // @[d_cache.scala 87:18 42:31]
  wire [63:0] _GEN_12975 = 3'h3 == state ? ram_0_0 : _GEN_11946; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12976 = 3'h3 == state ? ram_0_1 : _GEN_11947; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12977 = 3'h3 == state ? ram_0_2 : _GEN_11948; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12978 = 3'h3 == state ? ram_0_3 : _GEN_11949; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12979 = 3'h3 == state ? ram_0_4 : _GEN_11950; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12980 = 3'h3 == state ? ram_0_5 : _GEN_11951; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12981 = 3'h3 == state ? ram_0_6 : _GEN_11952; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12982 = 3'h3 == state ? ram_0_7 : _GEN_11953; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12983 = 3'h3 == state ? ram_0_8 : _GEN_11954; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12984 = 3'h3 == state ? ram_0_9 : _GEN_11955; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12985 = 3'h3 == state ? ram_0_10 : _GEN_11956; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12986 = 3'h3 == state ? ram_0_11 : _GEN_11957; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12987 = 3'h3 == state ? ram_0_12 : _GEN_11958; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12988 = 3'h3 == state ? ram_0_13 : _GEN_11959; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12989 = 3'h3 == state ? ram_0_14 : _GEN_11960; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12990 = 3'h3 == state ? ram_0_15 : _GEN_11961; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12991 = 3'h3 == state ? ram_0_16 : _GEN_11962; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12992 = 3'h3 == state ? ram_0_17 : _GEN_11963; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12993 = 3'h3 == state ? ram_0_18 : _GEN_11964; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12994 = 3'h3 == state ? ram_0_19 : _GEN_11965; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12995 = 3'h3 == state ? ram_0_20 : _GEN_11966; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12996 = 3'h3 == state ? ram_0_21 : _GEN_11967; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12997 = 3'h3 == state ? ram_0_22 : _GEN_11968; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12998 = 3'h3 == state ? ram_0_23 : _GEN_11969; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_12999 = 3'h3 == state ? ram_0_24 : _GEN_11970; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13000 = 3'h3 == state ? ram_0_25 : _GEN_11971; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13001 = 3'h3 == state ? ram_0_26 : _GEN_11972; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13002 = 3'h3 == state ? ram_0_27 : _GEN_11973; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13003 = 3'h3 == state ? ram_0_28 : _GEN_11974; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13004 = 3'h3 == state ? ram_0_29 : _GEN_11975; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13005 = 3'h3 == state ? ram_0_30 : _GEN_11976; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13006 = 3'h3 == state ? ram_0_31 : _GEN_11977; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13007 = 3'h3 == state ? ram_0_32 : _GEN_11978; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13008 = 3'h3 == state ? ram_0_33 : _GEN_11979; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13009 = 3'h3 == state ? ram_0_34 : _GEN_11980; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13010 = 3'h3 == state ? ram_0_35 : _GEN_11981; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13011 = 3'h3 == state ? ram_0_36 : _GEN_11982; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13012 = 3'h3 == state ? ram_0_37 : _GEN_11983; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13013 = 3'h3 == state ? ram_0_38 : _GEN_11984; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13014 = 3'h3 == state ? ram_0_39 : _GEN_11985; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13015 = 3'h3 == state ? ram_0_40 : _GEN_11986; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13016 = 3'h3 == state ? ram_0_41 : _GEN_11987; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13017 = 3'h3 == state ? ram_0_42 : _GEN_11988; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13018 = 3'h3 == state ? ram_0_43 : _GEN_11989; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13019 = 3'h3 == state ? ram_0_44 : _GEN_11990; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13020 = 3'h3 == state ? ram_0_45 : _GEN_11991; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13021 = 3'h3 == state ? ram_0_46 : _GEN_11992; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13022 = 3'h3 == state ? ram_0_47 : _GEN_11993; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13023 = 3'h3 == state ? ram_0_48 : _GEN_11994; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13024 = 3'h3 == state ? ram_0_49 : _GEN_11995; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13025 = 3'h3 == state ? ram_0_50 : _GEN_11996; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13026 = 3'h3 == state ? ram_0_51 : _GEN_11997; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13027 = 3'h3 == state ? ram_0_52 : _GEN_11998; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13028 = 3'h3 == state ? ram_0_53 : _GEN_11999; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13029 = 3'h3 == state ? ram_0_54 : _GEN_12000; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13030 = 3'h3 == state ? ram_0_55 : _GEN_12001; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13031 = 3'h3 == state ? ram_0_56 : _GEN_12002; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13032 = 3'h3 == state ? ram_0_57 : _GEN_12003; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13033 = 3'h3 == state ? ram_0_58 : _GEN_12004; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13034 = 3'h3 == state ? ram_0_59 : _GEN_12005; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13035 = 3'h3 == state ? ram_0_60 : _GEN_12006; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13036 = 3'h3 == state ? ram_0_61 : _GEN_12007; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13037 = 3'h3 == state ? ram_0_62 : _GEN_12008; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13038 = 3'h3 == state ? ram_0_63 : _GEN_12009; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13039 = 3'h3 == state ? ram_0_64 : _GEN_12010; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13040 = 3'h3 == state ? ram_0_65 : _GEN_12011; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13041 = 3'h3 == state ? ram_0_66 : _GEN_12012; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13042 = 3'h3 == state ? ram_0_67 : _GEN_12013; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13043 = 3'h3 == state ? ram_0_68 : _GEN_12014; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13044 = 3'h3 == state ? ram_0_69 : _GEN_12015; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13045 = 3'h3 == state ? ram_0_70 : _GEN_12016; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13046 = 3'h3 == state ? ram_0_71 : _GEN_12017; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13047 = 3'h3 == state ? ram_0_72 : _GEN_12018; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13048 = 3'h3 == state ? ram_0_73 : _GEN_12019; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13049 = 3'h3 == state ? ram_0_74 : _GEN_12020; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13050 = 3'h3 == state ? ram_0_75 : _GEN_12021; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13051 = 3'h3 == state ? ram_0_76 : _GEN_12022; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13052 = 3'h3 == state ? ram_0_77 : _GEN_12023; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13053 = 3'h3 == state ? ram_0_78 : _GEN_12024; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13054 = 3'h3 == state ? ram_0_79 : _GEN_12025; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13055 = 3'h3 == state ? ram_0_80 : _GEN_12026; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13056 = 3'h3 == state ? ram_0_81 : _GEN_12027; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13057 = 3'h3 == state ? ram_0_82 : _GEN_12028; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13058 = 3'h3 == state ? ram_0_83 : _GEN_12029; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13059 = 3'h3 == state ? ram_0_84 : _GEN_12030; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13060 = 3'h3 == state ? ram_0_85 : _GEN_12031; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13061 = 3'h3 == state ? ram_0_86 : _GEN_12032; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13062 = 3'h3 == state ? ram_0_87 : _GEN_12033; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13063 = 3'h3 == state ? ram_0_88 : _GEN_12034; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13064 = 3'h3 == state ? ram_0_89 : _GEN_12035; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13065 = 3'h3 == state ? ram_0_90 : _GEN_12036; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13066 = 3'h3 == state ? ram_0_91 : _GEN_12037; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13067 = 3'h3 == state ? ram_0_92 : _GEN_12038; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13068 = 3'h3 == state ? ram_0_93 : _GEN_12039; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13069 = 3'h3 == state ? ram_0_94 : _GEN_12040; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13070 = 3'h3 == state ? ram_0_95 : _GEN_12041; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13071 = 3'h3 == state ? ram_0_96 : _GEN_12042; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13072 = 3'h3 == state ? ram_0_97 : _GEN_12043; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13073 = 3'h3 == state ? ram_0_98 : _GEN_12044; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13074 = 3'h3 == state ? ram_0_99 : _GEN_12045; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13075 = 3'h3 == state ? ram_0_100 : _GEN_12046; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13076 = 3'h3 == state ? ram_0_101 : _GEN_12047; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13077 = 3'h3 == state ? ram_0_102 : _GEN_12048; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13078 = 3'h3 == state ? ram_0_103 : _GEN_12049; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13079 = 3'h3 == state ? ram_0_104 : _GEN_12050; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13080 = 3'h3 == state ? ram_0_105 : _GEN_12051; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13081 = 3'h3 == state ? ram_0_106 : _GEN_12052; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13082 = 3'h3 == state ? ram_0_107 : _GEN_12053; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13083 = 3'h3 == state ? ram_0_108 : _GEN_12054; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13084 = 3'h3 == state ? ram_0_109 : _GEN_12055; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13085 = 3'h3 == state ? ram_0_110 : _GEN_12056; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13086 = 3'h3 == state ? ram_0_111 : _GEN_12057; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13087 = 3'h3 == state ? ram_0_112 : _GEN_12058; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13088 = 3'h3 == state ? ram_0_113 : _GEN_12059; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13089 = 3'h3 == state ? ram_0_114 : _GEN_12060; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13090 = 3'h3 == state ? ram_0_115 : _GEN_12061; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13091 = 3'h3 == state ? ram_0_116 : _GEN_12062; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13092 = 3'h3 == state ? ram_0_117 : _GEN_12063; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13093 = 3'h3 == state ? ram_0_118 : _GEN_12064; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13094 = 3'h3 == state ? ram_0_119 : _GEN_12065; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13095 = 3'h3 == state ? ram_0_120 : _GEN_12066; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13096 = 3'h3 == state ? ram_0_121 : _GEN_12067; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13097 = 3'h3 == state ? ram_0_122 : _GEN_12068; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13098 = 3'h3 == state ? ram_0_123 : _GEN_12069; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13099 = 3'h3 == state ? ram_0_124 : _GEN_12070; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13100 = 3'h3 == state ? ram_0_125 : _GEN_12071; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13101 = 3'h3 == state ? ram_0_126 : _GEN_12072; // @[d_cache.scala 87:18 19:24]
  wire [63:0] _GEN_13102 = 3'h3 == state ? ram_0_127 : _GEN_12073; // @[d_cache.scala 87:18 19:24]
  wire [31:0] _GEN_13103 = 3'h3 == state ? tag_0_0 : _GEN_12074; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13104 = 3'h3 == state ? tag_0_1 : _GEN_12075; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13105 = 3'h3 == state ? tag_0_2 : _GEN_12076; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13106 = 3'h3 == state ? tag_0_3 : _GEN_12077; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13107 = 3'h3 == state ? tag_0_4 : _GEN_12078; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13108 = 3'h3 == state ? tag_0_5 : _GEN_12079; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13109 = 3'h3 == state ? tag_0_6 : _GEN_12080; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13110 = 3'h3 == state ? tag_0_7 : _GEN_12081; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13111 = 3'h3 == state ? tag_0_8 : _GEN_12082; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13112 = 3'h3 == state ? tag_0_9 : _GEN_12083; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13113 = 3'h3 == state ? tag_0_10 : _GEN_12084; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13114 = 3'h3 == state ? tag_0_11 : _GEN_12085; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13115 = 3'h3 == state ? tag_0_12 : _GEN_12086; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13116 = 3'h3 == state ? tag_0_13 : _GEN_12087; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13117 = 3'h3 == state ? tag_0_14 : _GEN_12088; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13118 = 3'h3 == state ? tag_0_15 : _GEN_12089; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13119 = 3'h3 == state ? tag_0_16 : _GEN_12090; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13120 = 3'h3 == state ? tag_0_17 : _GEN_12091; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13121 = 3'h3 == state ? tag_0_18 : _GEN_12092; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13122 = 3'h3 == state ? tag_0_19 : _GEN_12093; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13123 = 3'h3 == state ? tag_0_20 : _GEN_12094; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13124 = 3'h3 == state ? tag_0_21 : _GEN_12095; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13125 = 3'h3 == state ? tag_0_22 : _GEN_12096; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13126 = 3'h3 == state ? tag_0_23 : _GEN_12097; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13127 = 3'h3 == state ? tag_0_24 : _GEN_12098; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13128 = 3'h3 == state ? tag_0_25 : _GEN_12099; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13129 = 3'h3 == state ? tag_0_26 : _GEN_12100; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13130 = 3'h3 == state ? tag_0_27 : _GEN_12101; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13131 = 3'h3 == state ? tag_0_28 : _GEN_12102; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13132 = 3'h3 == state ? tag_0_29 : _GEN_12103; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13133 = 3'h3 == state ? tag_0_30 : _GEN_12104; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13134 = 3'h3 == state ? tag_0_31 : _GEN_12105; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13135 = 3'h3 == state ? tag_0_32 : _GEN_12106; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13136 = 3'h3 == state ? tag_0_33 : _GEN_12107; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13137 = 3'h3 == state ? tag_0_34 : _GEN_12108; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13138 = 3'h3 == state ? tag_0_35 : _GEN_12109; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13139 = 3'h3 == state ? tag_0_36 : _GEN_12110; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13140 = 3'h3 == state ? tag_0_37 : _GEN_12111; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13141 = 3'h3 == state ? tag_0_38 : _GEN_12112; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13142 = 3'h3 == state ? tag_0_39 : _GEN_12113; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13143 = 3'h3 == state ? tag_0_40 : _GEN_12114; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13144 = 3'h3 == state ? tag_0_41 : _GEN_12115; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13145 = 3'h3 == state ? tag_0_42 : _GEN_12116; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13146 = 3'h3 == state ? tag_0_43 : _GEN_12117; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13147 = 3'h3 == state ? tag_0_44 : _GEN_12118; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13148 = 3'h3 == state ? tag_0_45 : _GEN_12119; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13149 = 3'h3 == state ? tag_0_46 : _GEN_12120; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13150 = 3'h3 == state ? tag_0_47 : _GEN_12121; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13151 = 3'h3 == state ? tag_0_48 : _GEN_12122; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13152 = 3'h3 == state ? tag_0_49 : _GEN_12123; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13153 = 3'h3 == state ? tag_0_50 : _GEN_12124; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13154 = 3'h3 == state ? tag_0_51 : _GEN_12125; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13155 = 3'h3 == state ? tag_0_52 : _GEN_12126; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13156 = 3'h3 == state ? tag_0_53 : _GEN_12127; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13157 = 3'h3 == state ? tag_0_54 : _GEN_12128; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13158 = 3'h3 == state ? tag_0_55 : _GEN_12129; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13159 = 3'h3 == state ? tag_0_56 : _GEN_12130; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13160 = 3'h3 == state ? tag_0_57 : _GEN_12131; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13161 = 3'h3 == state ? tag_0_58 : _GEN_12132; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13162 = 3'h3 == state ? tag_0_59 : _GEN_12133; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13163 = 3'h3 == state ? tag_0_60 : _GEN_12134; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13164 = 3'h3 == state ? tag_0_61 : _GEN_12135; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13165 = 3'h3 == state ? tag_0_62 : _GEN_12136; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13166 = 3'h3 == state ? tag_0_63 : _GEN_12137; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13167 = 3'h3 == state ? tag_0_64 : _GEN_12138; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13168 = 3'h3 == state ? tag_0_65 : _GEN_12139; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13169 = 3'h3 == state ? tag_0_66 : _GEN_12140; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13170 = 3'h3 == state ? tag_0_67 : _GEN_12141; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13171 = 3'h3 == state ? tag_0_68 : _GEN_12142; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13172 = 3'h3 == state ? tag_0_69 : _GEN_12143; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13173 = 3'h3 == state ? tag_0_70 : _GEN_12144; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13174 = 3'h3 == state ? tag_0_71 : _GEN_12145; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13175 = 3'h3 == state ? tag_0_72 : _GEN_12146; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13176 = 3'h3 == state ? tag_0_73 : _GEN_12147; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13177 = 3'h3 == state ? tag_0_74 : _GEN_12148; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13178 = 3'h3 == state ? tag_0_75 : _GEN_12149; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13179 = 3'h3 == state ? tag_0_76 : _GEN_12150; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13180 = 3'h3 == state ? tag_0_77 : _GEN_12151; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13181 = 3'h3 == state ? tag_0_78 : _GEN_12152; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13182 = 3'h3 == state ? tag_0_79 : _GEN_12153; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13183 = 3'h3 == state ? tag_0_80 : _GEN_12154; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13184 = 3'h3 == state ? tag_0_81 : _GEN_12155; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13185 = 3'h3 == state ? tag_0_82 : _GEN_12156; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13186 = 3'h3 == state ? tag_0_83 : _GEN_12157; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13187 = 3'h3 == state ? tag_0_84 : _GEN_12158; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13188 = 3'h3 == state ? tag_0_85 : _GEN_12159; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13189 = 3'h3 == state ? tag_0_86 : _GEN_12160; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13190 = 3'h3 == state ? tag_0_87 : _GEN_12161; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13191 = 3'h3 == state ? tag_0_88 : _GEN_12162; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13192 = 3'h3 == state ? tag_0_89 : _GEN_12163; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13193 = 3'h3 == state ? tag_0_90 : _GEN_12164; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13194 = 3'h3 == state ? tag_0_91 : _GEN_12165; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13195 = 3'h3 == state ? tag_0_92 : _GEN_12166; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13196 = 3'h3 == state ? tag_0_93 : _GEN_12167; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13197 = 3'h3 == state ? tag_0_94 : _GEN_12168; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13198 = 3'h3 == state ? tag_0_95 : _GEN_12169; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13199 = 3'h3 == state ? tag_0_96 : _GEN_12170; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13200 = 3'h3 == state ? tag_0_97 : _GEN_12171; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13201 = 3'h3 == state ? tag_0_98 : _GEN_12172; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13202 = 3'h3 == state ? tag_0_99 : _GEN_12173; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13203 = 3'h3 == state ? tag_0_100 : _GEN_12174; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13204 = 3'h3 == state ? tag_0_101 : _GEN_12175; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13205 = 3'h3 == state ? tag_0_102 : _GEN_12176; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13206 = 3'h3 == state ? tag_0_103 : _GEN_12177; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13207 = 3'h3 == state ? tag_0_104 : _GEN_12178; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13208 = 3'h3 == state ? tag_0_105 : _GEN_12179; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13209 = 3'h3 == state ? tag_0_106 : _GEN_12180; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13210 = 3'h3 == state ? tag_0_107 : _GEN_12181; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13211 = 3'h3 == state ? tag_0_108 : _GEN_12182; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13212 = 3'h3 == state ? tag_0_109 : _GEN_12183; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13213 = 3'h3 == state ? tag_0_110 : _GEN_12184; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13214 = 3'h3 == state ? tag_0_111 : _GEN_12185; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13215 = 3'h3 == state ? tag_0_112 : _GEN_12186; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13216 = 3'h3 == state ? tag_0_113 : _GEN_12187; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13217 = 3'h3 == state ? tag_0_114 : _GEN_12188; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13218 = 3'h3 == state ? tag_0_115 : _GEN_12189; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13219 = 3'h3 == state ? tag_0_116 : _GEN_12190; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13220 = 3'h3 == state ? tag_0_117 : _GEN_12191; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13221 = 3'h3 == state ? tag_0_118 : _GEN_12192; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13222 = 3'h3 == state ? tag_0_119 : _GEN_12193; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13223 = 3'h3 == state ? tag_0_120 : _GEN_12194; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13224 = 3'h3 == state ? tag_0_121 : _GEN_12195; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13225 = 3'h3 == state ? tag_0_122 : _GEN_12196; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13226 = 3'h3 == state ? tag_0_123 : _GEN_12197; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13227 = 3'h3 == state ? tag_0_124 : _GEN_12198; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13228 = 3'h3 == state ? tag_0_125 : _GEN_12199; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13229 = 3'h3 == state ? tag_0_126 : _GEN_12200; // @[d_cache.scala 87:18 28:24]
  wire [31:0] _GEN_13230 = 3'h3 == state ? tag_0_127 : _GEN_12201; // @[d_cache.scala 87:18 28:24]
  wire  _GEN_13231 = 3'h3 == state ? valid_0_0 : _GEN_12202; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13232 = 3'h3 == state ? valid_0_1 : _GEN_12203; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13233 = 3'h3 == state ? valid_0_2 : _GEN_12204; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13234 = 3'h3 == state ? valid_0_3 : _GEN_12205; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13235 = 3'h3 == state ? valid_0_4 : _GEN_12206; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13236 = 3'h3 == state ? valid_0_5 : _GEN_12207; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13237 = 3'h3 == state ? valid_0_6 : _GEN_12208; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13238 = 3'h3 == state ? valid_0_7 : _GEN_12209; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13239 = 3'h3 == state ? valid_0_8 : _GEN_12210; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13240 = 3'h3 == state ? valid_0_9 : _GEN_12211; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13241 = 3'h3 == state ? valid_0_10 : _GEN_12212; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13242 = 3'h3 == state ? valid_0_11 : _GEN_12213; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13243 = 3'h3 == state ? valid_0_12 : _GEN_12214; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13244 = 3'h3 == state ? valid_0_13 : _GEN_12215; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13245 = 3'h3 == state ? valid_0_14 : _GEN_12216; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13246 = 3'h3 == state ? valid_0_15 : _GEN_12217; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13247 = 3'h3 == state ? valid_0_16 : _GEN_12218; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13248 = 3'h3 == state ? valid_0_17 : _GEN_12219; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13249 = 3'h3 == state ? valid_0_18 : _GEN_12220; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13250 = 3'h3 == state ? valid_0_19 : _GEN_12221; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13251 = 3'h3 == state ? valid_0_20 : _GEN_12222; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13252 = 3'h3 == state ? valid_0_21 : _GEN_12223; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13253 = 3'h3 == state ? valid_0_22 : _GEN_12224; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13254 = 3'h3 == state ? valid_0_23 : _GEN_12225; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13255 = 3'h3 == state ? valid_0_24 : _GEN_12226; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13256 = 3'h3 == state ? valid_0_25 : _GEN_12227; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13257 = 3'h3 == state ? valid_0_26 : _GEN_12228; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13258 = 3'h3 == state ? valid_0_27 : _GEN_12229; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13259 = 3'h3 == state ? valid_0_28 : _GEN_12230; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13260 = 3'h3 == state ? valid_0_29 : _GEN_12231; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13261 = 3'h3 == state ? valid_0_30 : _GEN_12232; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13262 = 3'h3 == state ? valid_0_31 : _GEN_12233; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13263 = 3'h3 == state ? valid_0_32 : _GEN_12234; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13264 = 3'h3 == state ? valid_0_33 : _GEN_12235; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13265 = 3'h3 == state ? valid_0_34 : _GEN_12236; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13266 = 3'h3 == state ? valid_0_35 : _GEN_12237; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13267 = 3'h3 == state ? valid_0_36 : _GEN_12238; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13268 = 3'h3 == state ? valid_0_37 : _GEN_12239; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13269 = 3'h3 == state ? valid_0_38 : _GEN_12240; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13270 = 3'h3 == state ? valid_0_39 : _GEN_12241; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13271 = 3'h3 == state ? valid_0_40 : _GEN_12242; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13272 = 3'h3 == state ? valid_0_41 : _GEN_12243; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13273 = 3'h3 == state ? valid_0_42 : _GEN_12244; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13274 = 3'h3 == state ? valid_0_43 : _GEN_12245; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13275 = 3'h3 == state ? valid_0_44 : _GEN_12246; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13276 = 3'h3 == state ? valid_0_45 : _GEN_12247; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13277 = 3'h3 == state ? valid_0_46 : _GEN_12248; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13278 = 3'h3 == state ? valid_0_47 : _GEN_12249; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13279 = 3'h3 == state ? valid_0_48 : _GEN_12250; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13280 = 3'h3 == state ? valid_0_49 : _GEN_12251; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13281 = 3'h3 == state ? valid_0_50 : _GEN_12252; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13282 = 3'h3 == state ? valid_0_51 : _GEN_12253; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13283 = 3'h3 == state ? valid_0_52 : _GEN_12254; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13284 = 3'h3 == state ? valid_0_53 : _GEN_12255; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13285 = 3'h3 == state ? valid_0_54 : _GEN_12256; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13286 = 3'h3 == state ? valid_0_55 : _GEN_12257; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13287 = 3'h3 == state ? valid_0_56 : _GEN_12258; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13288 = 3'h3 == state ? valid_0_57 : _GEN_12259; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13289 = 3'h3 == state ? valid_0_58 : _GEN_12260; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13290 = 3'h3 == state ? valid_0_59 : _GEN_12261; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13291 = 3'h3 == state ? valid_0_60 : _GEN_12262; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13292 = 3'h3 == state ? valid_0_61 : _GEN_12263; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13293 = 3'h3 == state ? valid_0_62 : _GEN_12264; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13294 = 3'h3 == state ? valid_0_63 : _GEN_12265; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13295 = 3'h3 == state ? valid_0_64 : _GEN_12266; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13296 = 3'h3 == state ? valid_0_65 : _GEN_12267; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13297 = 3'h3 == state ? valid_0_66 : _GEN_12268; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13298 = 3'h3 == state ? valid_0_67 : _GEN_12269; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13299 = 3'h3 == state ? valid_0_68 : _GEN_12270; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13300 = 3'h3 == state ? valid_0_69 : _GEN_12271; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13301 = 3'h3 == state ? valid_0_70 : _GEN_12272; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13302 = 3'h3 == state ? valid_0_71 : _GEN_12273; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13303 = 3'h3 == state ? valid_0_72 : _GEN_12274; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13304 = 3'h3 == state ? valid_0_73 : _GEN_12275; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13305 = 3'h3 == state ? valid_0_74 : _GEN_12276; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13306 = 3'h3 == state ? valid_0_75 : _GEN_12277; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13307 = 3'h3 == state ? valid_0_76 : _GEN_12278; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13308 = 3'h3 == state ? valid_0_77 : _GEN_12279; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13309 = 3'h3 == state ? valid_0_78 : _GEN_12280; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13310 = 3'h3 == state ? valid_0_79 : _GEN_12281; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13311 = 3'h3 == state ? valid_0_80 : _GEN_12282; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13312 = 3'h3 == state ? valid_0_81 : _GEN_12283; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13313 = 3'h3 == state ? valid_0_82 : _GEN_12284; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13314 = 3'h3 == state ? valid_0_83 : _GEN_12285; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13315 = 3'h3 == state ? valid_0_84 : _GEN_12286; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13316 = 3'h3 == state ? valid_0_85 : _GEN_12287; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13317 = 3'h3 == state ? valid_0_86 : _GEN_12288; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13318 = 3'h3 == state ? valid_0_87 : _GEN_12289; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13319 = 3'h3 == state ? valid_0_88 : _GEN_12290; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13320 = 3'h3 == state ? valid_0_89 : _GEN_12291; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13321 = 3'h3 == state ? valid_0_90 : _GEN_12292; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13322 = 3'h3 == state ? valid_0_91 : _GEN_12293; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13323 = 3'h3 == state ? valid_0_92 : _GEN_12294; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13324 = 3'h3 == state ? valid_0_93 : _GEN_12295; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13325 = 3'h3 == state ? valid_0_94 : _GEN_12296; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13326 = 3'h3 == state ? valid_0_95 : _GEN_12297; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13327 = 3'h3 == state ? valid_0_96 : _GEN_12298; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13328 = 3'h3 == state ? valid_0_97 : _GEN_12299; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13329 = 3'h3 == state ? valid_0_98 : _GEN_12300; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13330 = 3'h3 == state ? valid_0_99 : _GEN_12301; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13331 = 3'h3 == state ? valid_0_100 : _GEN_12302; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13332 = 3'h3 == state ? valid_0_101 : _GEN_12303; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13333 = 3'h3 == state ? valid_0_102 : _GEN_12304; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13334 = 3'h3 == state ? valid_0_103 : _GEN_12305; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13335 = 3'h3 == state ? valid_0_104 : _GEN_12306; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13336 = 3'h3 == state ? valid_0_105 : _GEN_12307; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13337 = 3'h3 == state ? valid_0_106 : _GEN_12308; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13338 = 3'h3 == state ? valid_0_107 : _GEN_12309; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13339 = 3'h3 == state ? valid_0_108 : _GEN_12310; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13340 = 3'h3 == state ? valid_0_109 : _GEN_12311; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13341 = 3'h3 == state ? valid_0_110 : _GEN_12312; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13342 = 3'h3 == state ? valid_0_111 : _GEN_12313; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13343 = 3'h3 == state ? valid_0_112 : _GEN_12314; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13344 = 3'h3 == state ? valid_0_113 : _GEN_12315; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13345 = 3'h3 == state ? valid_0_114 : _GEN_12316; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13346 = 3'h3 == state ? valid_0_115 : _GEN_12317; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13347 = 3'h3 == state ? valid_0_116 : _GEN_12318; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13348 = 3'h3 == state ? valid_0_117 : _GEN_12319; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13349 = 3'h3 == state ? valid_0_118 : _GEN_12320; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13350 = 3'h3 == state ? valid_0_119 : _GEN_12321; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13351 = 3'h3 == state ? valid_0_120 : _GEN_12322; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13352 = 3'h3 == state ? valid_0_121 : _GEN_12323; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13353 = 3'h3 == state ? valid_0_122 : _GEN_12324; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13354 = 3'h3 == state ? valid_0_123 : _GEN_12325; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13355 = 3'h3 == state ? valid_0_124 : _GEN_12326; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13356 = 3'h3 == state ? valid_0_125 : _GEN_12327; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13357 = 3'h3 == state ? valid_0_126 : _GEN_12328; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13358 = 3'h3 == state ? valid_0_127 : _GEN_12329; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_13359 = 3'h3 == state ? quene : _GEN_12330; // @[d_cache.scala 87:18 43:24]
  wire [63:0] _GEN_13360 = 3'h3 == state ? ram_1_0 : _GEN_12331; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13361 = 3'h3 == state ? ram_1_1 : _GEN_12332; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13362 = 3'h3 == state ? ram_1_2 : _GEN_12333; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13363 = 3'h3 == state ? ram_1_3 : _GEN_12334; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13364 = 3'h3 == state ? ram_1_4 : _GEN_12335; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13365 = 3'h3 == state ? ram_1_5 : _GEN_12336; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13366 = 3'h3 == state ? ram_1_6 : _GEN_12337; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13367 = 3'h3 == state ? ram_1_7 : _GEN_12338; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13368 = 3'h3 == state ? ram_1_8 : _GEN_12339; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13369 = 3'h3 == state ? ram_1_9 : _GEN_12340; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13370 = 3'h3 == state ? ram_1_10 : _GEN_12341; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13371 = 3'h3 == state ? ram_1_11 : _GEN_12342; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13372 = 3'h3 == state ? ram_1_12 : _GEN_12343; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13373 = 3'h3 == state ? ram_1_13 : _GEN_12344; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13374 = 3'h3 == state ? ram_1_14 : _GEN_12345; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13375 = 3'h3 == state ? ram_1_15 : _GEN_12346; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13376 = 3'h3 == state ? ram_1_16 : _GEN_12347; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13377 = 3'h3 == state ? ram_1_17 : _GEN_12348; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13378 = 3'h3 == state ? ram_1_18 : _GEN_12349; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13379 = 3'h3 == state ? ram_1_19 : _GEN_12350; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13380 = 3'h3 == state ? ram_1_20 : _GEN_12351; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13381 = 3'h3 == state ? ram_1_21 : _GEN_12352; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13382 = 3'h3 == state ? ram_1_22 : _GEN_12353; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13383 = 3'h3 == state ? ram_1_23 : _GEN_12354; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13384 = 3'h3 == state ? ram_1_24 : _GEN_12355; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13385 = 3'h3 == state ? ram_1_25 : _GEN_12356; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13386 = 3'h3 == state ? ram_1_26 : _GEN_12357; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13387 = 3'h3 == state ? ram_1_27 : _GEN_12358; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13388 = 3'h3 == state ? ram_1_28 : _GEN_12359; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13389 = 3'h3 == state ? ram_1_29 : _GEN_12360; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13390 = 3'h3 == state ? ram_1_30 : _GEN_12361; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13391 = 3'h3 == state ? ram_1_31 : _GEN_12362; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13392 = 3'h3 == state ? ram_1_32 : _GEN_12363; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13393 = 3'h3 == state ? ram_1_33 : _GEN_12364; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13394 = 3'h3 == state ? ram_1_34 : _GEN_12365; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13395 = 3'h3 == state ? ram_1_35 : _GEN_12366; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13396 = 3'h3 == state ? ram_1_36 : _GEN_12367; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13397 = 3'h3 == state ? ram_1_37 : _GEN_12368; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13398 = 3'h3 == state ? ram_1_38 : _GEN_12369; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13399 = 3'h3 == state ? ram_1_39 : _GEN_12370; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13400 = 3'h3 == state ? ram_1_40 : _GEN_12371; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13401 = 3'h3 == state ? ram_1_41 : _GEN_12372; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13402 = 3'h3 == state ? ram_1_42 : _GEN_12373; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13403 = 3'h3 == state ? ram_1_43 : _GEN_12374; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13404 = 3'h3 == state ? ram_1_44 : _GEN_12375; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13405 = 3'h3 == state ? ram_1_45 : _GEN_12376; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13406 = 3'h3 == state ? ram_1_46 : _GEN_12377; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13407 = 3'h3 == state ? ram_1_47 : _GEN_12378; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13408 = 3'h3 == state ? ram_1_48 : _GEN_12379; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13409 = 3'h3 == state ? ram_1_49 : _GEN_12380; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13410 = 3'h3 == state ? ram_1_50 : _GEN_12381; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13411 = 3'h3 == state ? ram_1_51 : _GEN_12382; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13412 = 3'h3 == state ? ram_1_52 : _GEN_12383; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13413 = 3'h3 == state ? ram_1_53 : _GEN_12384; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13414 = 3'h3 == state ? ram_1_54 : _GEN_12385; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13415 = 3'h3 == state ? ram_1_55 : _GEN_12386; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13416 = 3'h3 == state ? ram_1_56 : _GEN_12387; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13417 = 3'h3 == state ? ram_1_57 : _GEN_12388; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13418 = 3'h3 == state ? ram_1_58 : _GEN_12389; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13419 = 3'h3 == state ? ram_1_59 : _GEN_12390; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13420 = 3'h3 == state ? ram_1_60 : _GEN_12391; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13421 = 3'h3 == state ? ram_1_61 : _GEN_12392; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13422 = 3'h3 == state ? ram_1_62 : _GEN_12393; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13423 = 3'h3 == state ? ram_1_63 : _GEN_12394; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13424 = 3'h3 == state ? ram_1_64 : _GEN_12395; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13425 = 3'h3 == state ? ram_1_65 : _GEN_12396; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13426 = 3'h3 == state ? ram_1_66 : _GEN_12397; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13427 = 3'h3 == state ? ram_1_67 : _GEN_12398; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13428 = 3'h3 == state ? ram_1_68 : _GEN_12399; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13429 = 3'h3 == state ? ram_1_69 : _GEN_12400; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13430 = 3'h3 == state ? ram_1_70 : _GEN_12401; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13431 = 3'h3 == state ? ram_1_71 : _GEN_12402; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13432 = 3'h3 == state ? ram_1_72 : _GEN_12403; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13433 = 3'h3 == state ? ram_1_73 : _GEN_12404; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13434 = 3'h3 == state ? ram_1_74 : _GEN_12405; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13435 = 3'h3 == state ? ram_1_75 : _GEN_12406; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13436 = 3'h3 == state ? ram_1_76 : _GEN_12407; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13437 = 3'h3 == state ? ram_1_77 : _GEN_12408; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13438 = 3'h3 == state ? ram_1_78 : _GEN_12409; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13439 = 3'h3 == state ? ram_1_79 : _GEN_12410; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13440 = 3'h3 == state ? ram_1_80 : _GEN_12411; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13441 = 3'h3 == state ? ram_1_81 : _GEN_12412; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13442 = 3'h3 == state ? ram_1_82 : _GEN_12413; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13443 = 3'h3 == state ? ram_1_83 : _GEN_12414; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13444 = 3'h3 == state ? ram_1_84 : _GEN_12415; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13445 = 3'h3 == state ? ram_1_85 : _GEN_12416; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13446 = 3'h3 == state ? ram_1_86 : _GEN_12417; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13447 = 3'h3 == state ? ram_1_87 : _GEN_12418; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13448 = 3'h3 == state ? ram_1_88 : _GEN_12419; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13449 = 3'h3 == state ? ram_1_89 : _GEN_12420; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13450 = 3'h3 == state ? ram_1_90 : _GEN_12421; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13451 = 3'h3 == state ? ram_1_91 : _GEN_12422; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13452 = 3'h3 == state ? ram_1_92 : _GEN_12423; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13453 = 3'h3 == state ? ram_1_93 : _GEN_12424; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13454 = 3'h3 == state ? ram_1_94 : _GEN_12425; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13455 = 3'h3 == state ? ram_1_95 : _GEN_12426; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13456 = 3'h3 == state ? ram_1_96 : _GEN_12427; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13457 = 3'h3 == state ? ram_1_97 : _GEN_12428; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13458 = 3'h3 == state ? ram_1_98 : _GEN_12429; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13459 = 3'h3 == state ? ram_1_99 : _GEN_12430; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13460 = 3'h3 == state ? ram_1_100 : _GEN_12431; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13461 = 3'h3 == state ? ram_1_101 : _GEN_12432; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13462 = 3'h3 == state ? ram_1_102 : _GEN_12433; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13463 = 3'h3 == state ? ram_1_103 : _GEN_12434; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13464 = 3'h3 == state ? ram_1_104 : _GEN_12435; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13465 = 3'h3 == state ? ram_1_105 : _GEN_12436; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13466 = 3'h3 == state ? ram_1_106 : _GEN_12437; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13467 = 3'h3 == state ? ram_1_107 : _GEN_12438; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13468 = 3'h3 == state ? ram_1_108 : _GEN_12439; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13469 = 3'h3 == state ? ram_1_109 : _GEN_12440; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13470 = 3'h3 == state ? ram_1_110 : _GEN_12441; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13471 = 3'h3 == state ? ram_1_111 : _GEN_12442; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13472 = 3'h3 == state ? ram_1_112 : _GEN_12443; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13473 = 3'h3 == state ? ram_1_113 : _GEN_12444; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13474 = 3'h3 == state ? ram_1_114 : _GEN_12445; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13475 = 3'h3 == state ? ram_1_115 : _GEN_12446; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13476 = 3'h3 == state ? ram_1_116 : _GEN_12447; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13477 = 3'h3 == state ? ram_1_117 : _GEN_12448; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13478 = 3'h3 == state ? ram_1_118 : _GEN_12449; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13479 = 3'h3 == state ? ram_1_119 : _GEN_12450; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13480 = 3'h3 == state ? ram_1_120 : _GEN_12451; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13481 = 3'h3 == state ? ram_1_121 : _GEN_12452; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13482 = 3'h3 == state ? ram_1_122 : _GEN_12453; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13483 = 3'h3 == state ? ram_1_123 : _GEN_12454; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13484 = 3'h3 == state ? ram_1_124 : _GEN_12455; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13485 = 3'h3 == state ? ram_1_125 : _GEN_12456; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13486 = 3'h3 == state ? ram_1_126 : _GEN_12457; // @[d_cache.scala 87:18 20:24]
  wire [63:0] _GEN_13487 = 3'h3 == state ? ram_1_127 : _GEN_12458; // @[d_cache.scala 87:18 20:24]
  wire [31:0] _GEN_13488 = 3'h3 == state ? tag_1_0 : _GEN_12459; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13489 = 3'h3 == state ? tag_1_1 : _GEN_12460; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13490 = 3'h3 == state ? tag_1_2 : _GEN_12461; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13491 = 3'h3 == state ? tag_1_3 : _GEN_12462; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13492 = 3'h3 == state ? tag_1_4 : _GEN_12463; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13493 = 3'h3 == state ? tag_1_5 : _GEN_12464; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13494 = 3'h3 == state ? tag_1_6 : _GEN_12465; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13495 = 3'h3 == state ? tag_1_7 : _GEN_12466; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13496 = 3'h3 == state ? tag_1_8 : _GEN_12467; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13497 = 3'h3 == state ? tag_1_9 : _GEN_12468; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13498 = 3'h3 == state ? tag_1_10 : _GEN_12469; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13499 = 3'h3 == state ? tag_1_11 : _GEN_12470; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13500 = 3'h3 == state ? tag_1_12 : _GEN_12471; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13501 = 3'h3 == state ? tag_1_13 : _GEN_12472; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13502 = 3'h3 == state ? tag_1_14 : _GEN_12473; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13503 = 3'h3 == state ? tag_1_15 : _GEN_12474; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13504 = 3'h3 == state ? tag_1_16 : _GEN_12475; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13505 = 3'h3 == state ? tag_1_17 : _GEN_12476; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13506 = 3'h3 == state ? tag_1_18 : _GEN_12477; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13507 = 3'h3 == state ? tag_1_19 : _GEN_12478; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13508 = 3'h3 == state ? tag_1_20 : _GEN_12479; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13509 = 3'h3 == state ? tag_1_21 : _GEN_12480; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13510 = 3'h3 == state ? tag_1_22 : _GEN_12481; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13511 = 3'h3 == state ? tag_1_23 : _GEN_12482; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13512 = 3'h3 == state ? tag_1_24 : _GEN_12483; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13513 = 3'h3 == state ? tag_1_25 : _GEN_12484; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13514 = 3'h3 == state ? tag_1_26 : _GEN_12485; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13515 = 3'h3 == state ? tag_1_27 : _GEN_12486; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13516 = 3'h3 == state ? tag_1_28 : _GEN_12487; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13517 = 3'h3 == state ? tag_1_29 : _GEN_12488; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13518 = 3'h3 == state ? tag_1_30 : _GEN_12489; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13519 = 3'h3 == state ? tag_1_31 : _GEN_12490; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13520 = 3'h3 == state ? tag_1_32 : _GEN_12491; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13521 = 3'h3 == state ? tag_1_33 : _GEN_12492; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13522 = 3'h3 == state ? tag_1_34 : _GEN_12493; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13523 = 3'h3 == state ? tag_1_35 : _GEN_12494; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13524 = 3'h3 == state ? tag_1_36 : _GEN_12495; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13525 = 3'h3 == state ? tag_1_37 : _GEN_12496; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13526 = 3'h3 == state ? tag_1_38 : _GEN_12497; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13527 = 3'h3 == state ? tag_1_39 : _GEN_12498; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13528 = 3'h3 == state ? tag_1_40 : _GEN_12499; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13529 = 3'h3 == state ? tag_1_41 : _GEN_12500; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13530 = 3'h3 == state ? tag_1_42 : _GEN_12501; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13531 = 3'h3 == state ? tag_1_43 : _GEN_12502; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13532 = 3'h3 == state ? tag_1_44 : _GEN_12503; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13533 = 3'h3 == state ? tag_1_45 : _GEN_12504; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13534 = 3'h3 == state ? tag_1_46 : _GEN_12505; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13535 = 3'h3 == state ? tag_1_47 : _GEN_12506; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13536 = 3'h3 == state ? tag_1_48 : _GEN_12507; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13537 = 3'h3 == state ? tag_1_49 : _GEN_12508; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13538 = 3'h3 == state ? tag_1_50 : _GEN_12509; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13539 = 3'h3 == state ? tag_1_51 : _GEN_12510; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13540 = 3'h3 == state ? tag_1_52 : _GEN_12511; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13541 = 3'h3 == state ? tag_1_53 : _GEN_12512; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13542 = 3'h3 == state ? tag_1_54 : _GEN_12513; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13543 = 3'h3 == state ? tag_1_55 : _GEN_12514; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13544 = 3'h3 == state ? tag_1_56 : _GEN_12515; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13545 = 3'h3 == state ? tag_1_57 : _GEN_12516; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13546 = 3'h3 == state ? tag_1_58 : _GEN_12517; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13547 = 3'h3 == state ? tag_1_59 : _GEN_12518; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13548 = 3'h3 == state ? tag_1_60 : _GEN_12519; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13549 = 3'h3 == state ? tag_1_61 : _GEN_12520; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13550 = 3'h3 == state ? tag_1_62 : _GEN_12521; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13551 = 3'h3 == state ? tag_1_63 : _GEN_12522; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13552 = 3'h3 == state ? tag_1_64 : _GEN_12523; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13553 = 3'h3 == state ? tag_1_65 : _GEN_12524; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13554 = 3'h3 == state ? tag_1_66 : _GEN_12525; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13555 = 3'h3 == state ? tag_1_67 : _GEN_12526; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13556 = 3'h3 == state ? tag_1_68 : _GEN_12527; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13557 = 3'h3 == state ? tag_1_69 : _GEN_12528; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13558 = 3'h3 == state ? tag_1_70 : _GEN_12529; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13559 = 3'h3 == state ? tag_1_71 : _GEN_12530; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13560 = 3'h3 == state ? tag_1_72 : _GEN_12531; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13561 = 3'h3 == state ? tag_1_73 : _GEN_12532; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13562 = 3'h3 == state ? tag_1_74 : _GEN_12533; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13563 = 3'h3 == state ? tag_1_75 : _GEN_12534; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13564 = 3'h3 == state ? tag_1_76 : _GEN_12535; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13565 = 3'h3 == state ? tag_1_77 : _GEN_12536; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13566 = 3'h3 == state ? tag_1_78 : _GEN_12537; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13567 = 3'h3 == state ? tag_1_79 : _GEN_12538; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13568 = 3'h3 == state ? tag_1_80 : _GEN_12539; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13569 = 3'h3 == state ? tag_1_81 : _GEN_12540; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13570 = 3'h3 == state ? tag_1_82 : _GEN_12541; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13571 = 3'h3 == state ? tag_1_83 : _GEN_12542; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13572 = 3'h3 == state ? tag_1_84 : _GEN_12543; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13573 = 3'h3 == state ? tag_1_85 : _GEN_12544; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13574 = 3'h3 == state ? tag_1_86 : _GEN_12545; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13575 = 3'h3 == state ? tag_1_87 : _GEN_12546; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13576 = 3'h3 == state ? tag_1_88 : _GEN_12547; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13577 = 3'h3 == state ? tag_1_89 : _GEN_12548; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13578 = 3'h3 == state ? tag_1_90 : _GEN_12549; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13579 = 3'h3 == state ? tag_1_91 : _GEN_12550; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13580 = 3'h3 == state ? tag_1_92 : _GEN_12551; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13581 = 3'h3 == state ? tag_1_93 : _GEN_12552; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13582 = 3'h3 == state ? tag_1_94 : _GEN_12553; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13583 = 3'h3 == state ? tag_1_95 : _GEN_12554; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13584 = 3'h3 == state ? tag_1_96 : _GEN_12555; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13585 = 3'h3 == state ? tag_1_97 : _GEN_12556; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13586 = 3'h3 == state ? tag_1_98 : _GEN_12557; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13587 = 3'h3 == state ? tag_1_99 : _GEN_12558; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13588 = 3'h3 == state ? tag_1_100 : _GEN_12559; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13589 = 3'h3 == state ? tag_1_101 : _GEN_12560; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13590 = 3'h3 == state ? tag_1_102 : _GEN_12561; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13591 = 3'h3 == state ? tag_1_103 : _GEN_12562; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13592 = 3'h3 == state ? tag_1_104 : _GEN_12563; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13593 = 3'h3 == state ? tag_1_105 : _GEN_12564; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13594 = 3'h3 == state ? tag_1_106 : _GEN_12565; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13595 = 3'h3 == state ? tag_1_107 : _GEN_12566; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13596 = 3'h3 == state ? tag_1_108 : _GEN_12567; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13597 = 3'h3 == state ? tag_1_109 : _GEN_12568; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13598 = 3'h3 == state ? tag_1_110 : _GEN_12569; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13599 = 3'h3 == state ? tag_1_111 : _GEN_12570; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13600 = 3'h3 == state ? tag_1_112 : _GEN_12571; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13601 = 3'h3 == state ? tag_1_113 : _GEN_12572; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13602 = 3'h3 == state ? tag_1_114 : _GEN_12573; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13603 = 3'h3 == state ? tag_1_115 : _GEN_12574; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13604 = 3'h3 == state ? tag_1_116 : _GEN_12575; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13605 = 3'h3 == state ? tag_1_117 : _GEN_12576; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13606 = 3'h3 == state ? tag_1_118 : _GEN_12577; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13607 = 3'h3 == state ? tag_1_119 : _GEN_12578; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13608 = 3'h3 == state ? tag_1_120 : _GEN_12579; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13609 = 3'h3 == state ? tag_1_121 : _GEN_12580; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13610 = 3'h3 == state ? tag_1_122 : _GEN_12581; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13611 = 3'h3 == state ? tag_1_123 : _GEN_12582; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13612 = 3'h3 == state ? tag_1_124 : _GEN_12583; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13613 = 3'h3 == state ? tag_1_125 : _GEN_12584; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13614 = 3'h3 == state ? tag_1_126 : _GEN_12585; // @[d_cache.scala 87:18 29:24]
  wire [31:0] _GEN_13615 = 3'h3 == state ? tag_1_127 : _GEN_12586; // @[d_cache.scala 87:18 29:24]
  wire  _GEN_13616 = 3'h3 == state ? valid_1_0 : _GEN_12587; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13617 = 3'h3 == state ? valid_1_1 : _GEN_12588; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13618 = 3'h3 == state ? valid_1_2 : _GEN_12589; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13619 = 3'h3 == state ? valid_1_3 : _GEN_12590; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13620 = 3'h3 == state ? valid_1_4 : _GEN_12591; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13621 = 3'h3 == state ? valid_1_5 : _GEN_12592; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13622 = 3'h3 == state ? valid_1_6 : _GEN_12593; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13623 = 3'h3 == state ? valid_1_7 : _GEN_12594; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13624 = 3'h3 == state ? valid_1_8 : _GEN_12595; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13625 = 3'h3 == state ? valid_1_9 : _GEN_12596; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13626 = 3'h3 == state ? valid_1_10 : _GEN_12597; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13627 = 3'h3 == state ? valid_1_11 : _GEN_12598; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13628 = 3'h3 == state ? valid_1_12 : _GEN_12599; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13629 = 3'h3 == state ? valid_1_13 : _GEN_12600; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13630 = 3'h3 == state ? valid_1_14 : _GEN_12601; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13631 = 3'h3 == state ? valid_1_15 : _GEN_12602; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13632 = 3'h3 == state ? valid_1_16 : _GEN_12603; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13633 = 3'h3 == state ? valid_1_17 : _GEN_12604; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13634 = 3'h3 == state ? valid_1_18 : _GEN_12605; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13635 = 3'h3 == state ? valid_1_19 : _GEN_12606; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13636 = 3'h3 == state ? valid_1_20 : _GEN_12607; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13637 = 3'h3 == state ? valid_1_21 : _GEN_12608; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13638 = 3'h3 == state ? valid_1_22 : _GEN_12609; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13639 = 3'h3 == state ? valid_1_23 : _GEN_12610; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13640 = 3'h3 == state ? valid_1_24 : _GEN_12611; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13641 = 3'h3 == state ? valid_1_25 : _GEN_12612; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13642 = 3'h3 == state ? valid_1_26 : _GEN_12613; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13643 = 3'h3 == state ? valid_1_27 : _GEN_12614; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13644 = 3'h3 == state ? valid_1_28 : _GEN_12615; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13645 = 3'h3 == state ? valid_1_29 : _GEN_12616; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13646 = 3'h3 == state ? valid_1_30 : _GEN_12617; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13647 = 3'h3 == state ? valid_1_31 : _GEN_12618; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13648 = 3'h3 == state ? valid_1_32 : _GEN_12619; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13649 = 3'h3 == state ? valid_1_33 : _GEN_12620; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13650 = 3'h3 == state ? valid_1_34 : _GEN_12621; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13651 = 3'h3 == state ? valid_1_35 : _GEN_12622; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13652 = 3'h3 == state ? valid_1_36 : _GEN_12623; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13653 = 3'h3 == state ? valid_1_37 : _GEN_12624; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13654 = 3'h3 == state ? valid_1_38 : _GEN_12625; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13655 = 3'h3 == state ? valid_1_39 : _GEN_12626; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13656 = 3'h3 == state ? valid_1_40 : _GEN_12627; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13657 = 3'h3 == state ? valid_1_41 : _GEN_12628; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13658 = 3'h3 == state ? valid_1_42 : _GEN_12629; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13659 = 3'h3 == state ? valid_1_43 : _GEN_12630; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13660 = 3'h3 == state ? valid_1_44 : _GEN_12631; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13661 = 3'h3 == state ? valid_1_45 : _GEN_12632; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13662 = 3'h3 == state ? valid_1_46 : _GEN_12633; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13663 = 3'h3 == state ? valid_1_47 : _GEN_12634; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13664 = 3'h3 == state ? valid_1_48 : _GEN_12635; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13665 = 3'h3 == state ? valid_1_49 : _GEN_12636; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13666 = 3'h3 == state ? valid_1_50 : _GEN_12637; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13667 = 3'h3 == state ? valid_1_51 : _GEN_12638; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13668 = 3'h3 == state ? valid_1_52 : _GEN_12639; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13669 = 3'h3 == state ? valid_1_53 : _GEN_12640; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13670 = 3'h3 == state ? valid_1_54 : _GEN_12641; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13671 = 3'h3 == state ? valid_1_55 : _GEN_12642; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13672 = 3'h3 == state ? valid_1_56 : _GEN_12643; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13673 = 3'h3 == state ? valid_1_57 : _GEN_12644; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13674 = 3'h3 == state ? valid_1_58 : _GEN_12645; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13675 = 3'h3 == state ? valid_1_59 : _GEN_12646; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13676 = 3'h3 == state ? valid_1_60 : _GEN_12647; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13677 = 3'h3 == state ? valid_1_61 : _GEN_12648; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13678 = 3'h3 == state ? valid_1_62 : _GEN_12649; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13679 = 3'h3 == state ? valid_1_63 : _GEN_12650; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13680 = 3'h3 == state ? valid_1_64 : _GEN_12651; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13681 = 3'h3 == state ? valid_1_65 : _GEN_12652; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13682 = 3'h3 == state ? valid_1_66 : _GEN_12653; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13683 = 3'h3 == state ? valid_1_67 : _GEN_12654; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13684 = 3'h3 == state ? valid_1_68 : _GEN_12655; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13685 = 3'h3 == state ? valid_1_69 : _GEN_12656; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13686 = 3'h3 == state ? valid_1_70 : _GEN_12657; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13687 = 3'h3 == state ? valid_1_71 : _GEN_12658; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13688 = 3'h3 == state ? valid_1_72 : _GEN_12659; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13689 = 3'h3 == state ? valid_1_73 : _GEN_12660; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13690 = 3'h3 == state ? valid_1_74 : _GEN_12661; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13691 = 3'h3 == state ? valid_1_75 : _GEN_12662; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13692 = 3'h3 == state ? valid_1_76 : _GEN_12663; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13693 = 3'h3 == state ? valid_1_77 : _GEN_12664; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13694 = 3'h3 == state ? valid_1_78 : _GEN_12665; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13695 = 3'h3 == state ? valid_1_79 : _GEN_12666; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13696 = 3'h3 == state ? valid_1_80 : _GEN_12667; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13697 = 3'h3 == state ? valid_1_81 : _GEN_12668; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13698 = 3'h3 == state ? valid_1_82 : _GEN_12669; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13699 = 3'h3 == state ? valid_1_83 : _GEN_12670; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13700 = 3'h3 == state ? valid_1_84 : _GEN_12671; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13701 = 3'h3 == state ? valid_1_85 : _GEN_12672; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13702 = 3'h3 == state ? valid_1_86 : _GEN_12673; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13703 = 3'h3 == state ? valid_1_87 : _GEN_12674; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13704 = 3'h3 == state ? valid_1_88 : _GEN_12675; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13705 = 3'h3 == state ? valid_1_89 : _GEN_12676; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13706 = 3'h3 == state ? valid_1_90 : _GEN_12677; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13707 = 3'h3 == state ? valid_1_91 : _GEN_12678; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13708 = 3'h3 == state ? valid_1_92 : _GEN_12679; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13709 = 3'h3 == state ? valid_1_93 : _GEN_12680; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13710 = 3'h3 == state ? valid_1_94 : _GEN_12681; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13711 = 3'h3 == state ? valid_1_95 : _GEN_12682; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13712 = 3'h3 == state ? valid_1_96 : _GEN_12683; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13713 = 3'h3 == state ? valid_1_97 : _GEN_12684; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13714 = 3'h3 == state ? valid_1_98 : _GEN_12685; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13715 = 3'h3 == state ? valid_1_99 : _GEN_12686; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13716 = 3'h3 == state ? valid_1_100 : _GEN_12687; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13717 = 3'h3 == state ? valid_1_101 : _GEN_12688; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13718 = 3'h3 == state ? valid_1_102 : _GEN_12689; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13719 = 3'h3 == state ? valid_1_103 : _GEN_12690; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13720 = 3'h3 == state ? valid_1_104 : _GEN_12691; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13721 = 3'h3 == state ? valid_1_105 : _GEN_12692; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13722 = 3'h3 == state ? valid_1_106 : _GEN_12693; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13723 = 3'h3 == state ? valid_1_107 : _GEN_12694; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13724 = 3'h3 == state ? valid_1_108 : _GEN_12695; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13725 = 3'h3 == state ? valid_1_109 : _GEN_12696; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13726 = 3'h3 == state ? valid_1_110 : _GEN_12697; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13727 = 3'h3 == state ? valid_1_111 : _GEN_12698; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13728 = 3'h3 == state ? valid_1_112 : _GEN_12699; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13729 = 3'h3 == state ? valid_1_113 : _GEN_12700; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13730 = 3'h3 == state ? valid_1_114 : _GEN_12701; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13731 = 3'h3 == state ? valid_1_115 : _GEN_12702; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13732 = 3'h3 == state ? valid_1_116 : _GEN_12703; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13733 = 3'h3 == state ? valid_1_117 : _GEN_12704; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13734 = 3'h3 == state ? valid_1_118 : _GEN_12705; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13735 = 3'h3 == state ? valid_1_119 : _GEN_12706; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13736 = 3'h3 == state ? valid_1_120 : _GEN_12707; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13737 = 3'h3 == state ? valid_1_121 : _GEN_12708; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13738 = 3'h3 == state ? valid_1_122 : _GEN_12709; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13739 = 3'h3 == state ? valid_1_123 : _GEN_12710; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13740 = 3'h3 == state ? valid_1_124 : _GEN_12711; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13741 = 3'h3 == state ? valid_1_125 : _GEN_12712; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13742 = 3'h3 == state ? valid_1_126 : _GEN_12713; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_13743 = 3'h3 == state ? valid_1_127 : _GEN_12714; // @[d_cache.scala 87:18 31:26]
  wire [63:0] _GEN_13744 = 3'h3 == state ? write_back_data : _GEN_12715; // @[d_cache.scala 87:18 37:34]
  wire [41:0] _GEN_13745 = 3'h3 == state ? {{10'd0}, write_back_addr} : _GEN_12716; // @[d_cache.scala 87:18 38:34]
  wire  _GEN_13746 = 3'h3 == state ? dirty_0_0 : _GEN_12717; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13747 = 3'h3 == state ? dirty_0_1 : _GEN_12718; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13748 = 3'h3 == state ? dirty_0_2 : _GEN_12719; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13749 = 3'h3 == state ? dirty_0_3 : _GEN_12720; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13750 = 3'h3 == state ? dirty_0_4 : _GEN_12721; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13751 = 3'h3 == state ? dirty_0_5 : _GEN_12722; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13752 = 3'h3 == state ? dirty_0_6 : _GEN_12723; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13753 = 3'h3 == state ? dirty_0_7 : _GEN_12724; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13754 = 3'h3 == state ? dirty_0_8 : _GEN_12725; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13755 = 3'h3 == state ? dirty_0_9 : _GEN_12726; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13756 = 3'h3 == state ? dirty_0_10 : _GEN_12727; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13757 = 3'h3 == state ? dirty_0_11 : _GEN_12728; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13758 = 3'h3 == state ? dirty_0_12 : _GEN_12729; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13759 = 3'h3 == state ? dirty_0_13 : _GEN_12730; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13760 = 3'h3 == state ? dirty_0_14 : _GEN_12731; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13761 = 3'h3 == state ? dirty_0_15 : _GEN_12732; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13762 = 3'h3 == state ? dirty_0_16 : _GEN_12733; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13763 = 3'h3 == state ? dirty_0_17 : _GEN_12734; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13764 = 3'h3 == state ? dirty_0_18 : _GEN_12735; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13765 = 3'h3 == state ? dirty_0_19 : _GEN_12736; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13766 = 3'h3 == state ? dirty_0_20 : _GEN_12737; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13767 = 3'h3 == state ? dirty_0_21 : _GEN_12738; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13768 = 3'h3 == state ? dirty_0_22 : _GEN_12739; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13769 = 3'h3 == state ? dirty_0_23 : _GEN_12740; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13770 = 3'h3 == state ? dirty_0_24 : _GEN_12741; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13771 = 3'h3 == state ? dirty_0_25 : _GEN_12742; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13772 = 3'h3 == state ? dirty_0_26 : _GEN_12743; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13773 = 3'h3 == state ? dirty_0_27 : _GEN_12744; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13774 = 3'h3 == state ? dirty_0_28 : _GEN_12745; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13775 = 3'h3 == state ? dirty_0_29 : _GEN_12746; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13776 = 3'h3 == state ? dirty_0_30 : _GEN_12747; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13777 = 3'h3 == state ? dirty_0_31 : _GEN_12748; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13778 = 3'h3 == state ? dirty_0_32 : _GEN_12749; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13779 = 3'h3 == state ? dirty_0_33 : _GEN_12750; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13780 = 3'h3 == state ? dirty_0_34 : _GEN_12751; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13781 = 3'h3 == state ? dirty_0_35 : _GEN_12752; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13782 = 3'h3 == state ? dirty_0_36 : _GEN_12753; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13783 = 3'h3 == state ? dirty_0_37 : _GEN_12754; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13784 = 3'h3 == state ? dirty_0_38 : _GEN_12755; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13785 = 3'h3 == state ? dirty_0_39 : _GEN_12756; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13786 = 3'h3 == state ? dirty_0_40 : _GEN_12757; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13787 = 3'h3 == state ? dirty_0_41 : _GEN_12758; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13788 = 3'h3 == state ? dirty_0_42 : _GEN_12759; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13789 = 3'h3 == state ? dirty_0_43 : _GEN_12760; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13790 = 3'h3 == state ? dirty_0_44 : _GEN_12761; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13791 = 3'h3 == state ? dirty_0_45 : _GEN_12762; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13792 = 3'h3 == state ? dirty_0_46 : _GEN_12763; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13793 = 3'h3 == state ? dirty_0_47 : _GEN_12764; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13794 = 3'h3 == state ? dirty_0_48 : _GEN_12765; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13795 = 3'h3 == state ? dirty_0_49 : _GEN_12766; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13796 = 3'h3 == state ? dirty_0_50 : _GEN_12767; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13797 = 3'h3 == state ? dirty_0_51 : _GEN_12768; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13798 = 3'h3 == state ? dirty_0_52 : _GEN_12769; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13799 = 3'h3 == state ? dirty_0_53 : _GEN_12770; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13800 = 3'h3 == state ? dirty_0_54 : _GEN_12771; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13801 = 3'h3 == state ? dirty_0_55 : _GEN_12772; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13802 = 3'h3 == state ? dirty_0_56 : _GEN_12773; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13803 = 3'h3 == state ? dirty_0_57 : _GEN_12774; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13804 = 3'h3 == state ? dirty_0_58 : _GEN_12775; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13805 = 3'h3 == state ? dirty_0_59 : _GEN_12776; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13806 = 3'h3 == state ? dirty_0_60 : _GEN_12777; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13807 = 3'h3 == state ? dirty_0_61 : _GEN_12778; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13808 = 3'h3 == state ? dirty_0_62 : _GEN_12779; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13809 = 3'h3 == state ? dirty_0_63 : _GEN_12780; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13810 = 3'h3 == state ? dirty_0_64 : _GEN_12781; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13811 = 3'h3 == state ? dirty_0_65 : _GEN_12782; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13812 = 3'h3 == state ? dirty_0_66 : _GEN_12783; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13813 = 3'h3 == state ? dirty_0_67 : _GEN_12784; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13814 = 3'h3 == state ? dirty_0_68 : _GEN_12785; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13815 = 3'h3 == state ? dirty_0_69 : _GEN_12786; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13816 = 3'h3 == state ? dirty_0_70 : _GEN_12787; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13817 = 3'h3 == state ? dirty_0_71 : _GEN_12788; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13818 = 3'h3 == state ? dirty_0_72 : _GEN_12789; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13819 = 3'h3 == state ? dirty_0_73 : _GEN_12790; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13820 = 3'h3 == state ? dirty_0_74 : _GEN_12791; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13821 = 3'h3 == state ? dirty_0_75 : _GEN_12792; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13822 = 3'h3 == state ? dirty_0_76 : _GEN_12793; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13823 = 3'h3 == state ? dirty_0_77 : _GEN_12794; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13824 = 3'h3 == state ? dirty_0_78 : _GEN_12795; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13825 = 3'h3 == state ? dirty_0_79 : _GEN_12796; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13826 = 3'h3 == state ? dirty_0_80 : _GEN_12797; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13827 = 3'h3 == state ? dirty_0_81 : _GEN_12798; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13828 = 3'h3 == state ? dirty_0_82 : _GEN_12799; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13829 = 3'h3 == state ? dirty_0_83 : _GEN_12800; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13830 = 3'h3 == state ? dirty_0_84 : _GEN_12801; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13831 = 3'h3 == state ? dirty_0_85 : _GEN_12802; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13832 = 3'h3 == state ? dirty_0_86 : _GEN_12803; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13833 = 3'h3 == state ? dirty_0_87 : _GEN_12804; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13834 = 3'h3 == state ? dirty_0_88 : _GEN_12805; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13835 = 3'h3 == state ? dirty_0_89 : _GEN_12806; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13836 = 3'h3 == state ? dirty_0_90 : _GEN_12807; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13837 = 3'h3 == state ? dirty_0_91 : _GEN_12808; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13838 = 3'h3 == state ? dirty_0_92 : _GEN_12809; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13839 = 3'h3 == state ? dirty_0_93 : _GEN_12810; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13840 = 3'h3 == state ? dirty_0_94 : _GEN_12811; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13841 = 3'h3 == state ? dirty_0_95 : _GEN_12812; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13842 = 3'h3 == state ? dirty_0_96 : _GEN_12813; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13843 = 3'h3 == state ? dirty_0_97 : _GEN_12814; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13844 = 3'h3 == state ? dirty_0_98 : _GEN_12815; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13845 = 3'h3 == state ? dirty_0_99 : _GEN_12816; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13846 = 3'h3 == state ? dirty_0_100 : _GEN_12817; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13847 = 3'h3 == state ? dirty_0_101 : _GEN_12818; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13848 = 3'h3 == state ? dirty_0_102 : _GEN_12819; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13849 = 3'h3 == state ? dirty_0_103 : _GEN_12820; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13850 = 3'h3 == state ? dirty_0_104 : _GEN_12821; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13851 = 3'h3 == state ? dirty_0_105 : _GEN_12822; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13852 = 3'h3 == state ? dirty_0_106 : _GEN_12823; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13853 = 3'h3 == state ? dirty_0_107 : _GEN_12824; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13854 = 3'h3 == state ? dirty_0_108 : _GEN_12825; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13855 = 3'h3 == state ? dirty_0_109 : _GEN_12826; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13856 = 3'h3 == state ? dirty_0_110 : _GEN_12827; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13857 = 3'h3 == state ? dirty_0_111 : _GEN_12828; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13858 = 3'h3 == state ? dirty_0_112 : _GEN_12829; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13859 = 3'h3 == state ? dirty_0_113 : _GEN_12830; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13860 = 3'h3 == state ? dirty_0_114 : _GEN_12831; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13861 = 3'h3 == state ? dirty_0_115 : _GEN_12832; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13862 = 3'h3 == state ? dirty_0_116 : _GEN_12833; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13863 = 3'h3 == state ? dirty_0_117 : _GEN_12834; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13864 = 3'h3 == state ? dirty_0_118 : _GEN_12835; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13865 = 3'h3 == state ? dirty_0_119 : _GEN_12836; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13866 = 3'h3 == state ? dirty_0_120 : _GEN_12837; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13867 = 3'h3 == state ? dirty_0_121 : _GEN_12838; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13868 = 3'h3 == state ? dirty_0_122 : _GEN_12839; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13869 = 3'h3 == state ? dirty_0_123 : _GEN_12840; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13870 = 3'h3 == state ? dirty_0_124 : _GEN_12841; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13871 = 3'h3 == state ? dirty_0_125 : _GEN_12842; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13872 = 3'h3 == state ? dirty_0_126 : _GEN_12843; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13873 = 3'h3 == state ? dirty_0_127 : _GEN_12844; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_13874 = 3'h3 == state ? dirty_1_0 : _GEN_12845; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13875 = 3'h3 == state ? dirty_1_1 : _GEN_12846; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13876 = 3'h3 == state ? dirty_1_2 : _GEN_12847; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13877 = 3'h3 == state ? dirty_1_3 : _GEN_12848; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13878 = 3'h3 == state ? dirty_1_4 : _GEN_12849; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13879 = 3'h3 == state ? dirty_1_5 : _GEN_12850; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13880 = 3'h3 == state ? dirty_1_6 : _GEN_12851; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13881 = 3'h3 == state ? dirty_1_7 : _GEN_12852; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13882 = 3'h3 == state ? dirty_1_8 : _GEN_12853; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13883 = 3'h3 == state ? dirty_1_9 : _GEN_12854; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13884 = 3'h3 == state ? dirty_1_10 : _GEN_12855; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13885 = 3'h3 == state ? dirty_1_11 : _GEN_12856; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13886 = 3'h3 == state ? dirty_1_12 : _GEN_12857; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13887 = 3'h3 == state ? dirty_1_13 : _GEN_12858; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13888 = 3'h3 == state ? dirty_1_14 : _GEN_12859; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13889 = 3'h3 == state ? dirty_1_15 : _GEN_12860; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13890 = 3'h3 == state ? dirty_1_16 : _GEN_12861; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13891 = 3'h3 == state ? dirty_1_17 : _GEN_12862; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13892 = 3'h3 == state ? dirty_1_18 : _GEN_12863; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13893 = 3'h3 == state ? dirty_1_19 : _GEN_12864; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13894 = 3'h3 == state ? dirty_1_20 : _GEN_12865; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13895 = 3'h3 == state ? dirty_1_21 : _GEN_12866; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13896 = 3'h3 == state ? dirty_1_22 : _GEN_12867; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13897 = 3'h3 == state ? dirty_1_23 : _GEN_12868; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13898 = 3'h3 == state ? dirty_1_24 : _GEN_12869; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13899 = 3'h3 == state ? dirty_1_25 : _GEN_12870; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13900 = 3'h3 == state ? dirty_1_26 : _GEN_12871; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13901 = 3'h3 == state ? dirty_1_27 : _GEN_12872; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13902 = 3'h3 == state ? dirty_1_28 : _GEN_12873; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13903 = 3'h3 == state ? dirty_1_29 : _GEN_12874; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13904 = 3'h3 == state ? dirty_1_30 : _GEN_12875; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13905 = 3'h3 == state ? dirty_1_31 : _GEN_12876; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13906 = 3'h3 == state ? dirty_1_32 : _GEN_12877; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13907 = 3'h3 == state ? dirty_1_33 : _GEN_12878; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13908 = 3'h3 == state ? dirty_1_34 : _GEN_12879; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13909 = 3'h3 == state ? dirty_1_35 : _GEN_12880; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13910 = 3'h3 == state ? dirty_1_36 : _GEN_12881; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13911 = 3'h3 == state ? dirty_1_37 : _GEN_12882; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13912 = 3'h3 == state ? dirty_1_38 : _GEN_12883; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13913 = 3'h3 == state ? dirty_1_39 : _GEN_12884; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13914 = 3'h3 == state ? dirty_1_40 : _GEN_12885; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13915 = 3'h3 == state ? dirty_1_41 : _GEN_12886; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13916 = 3'h3 == state ? dirty_1_42 : _GEN_12887; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13917 = 3'h3 == state ? dirty_1_43 : _GEN_12888; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13918 = 3'h3 == state ? dirty_1_44 : _GEN_12889; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13919 = 3'h3 == state ? dirty_1_45 : _GEN_12890; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13920 = 3'h3 == state ? dirty_1_46 : _GEN_12891; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13921 = 3'h3 == state ? dirty_1_47 : _GEN_12892; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13922 = 3'h3 == state ? dirty_1_48 : _GEN_12893; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13923 = 3'h3 == state ? dirty_1_49 : _GEN_12894; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13924 = 3'h3 == state ? dirty_1_50 : _GEN_12895; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13925 = 3'h3 == state ? dirty_1_51 : _GEN_12896; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13926 = 3'h3 == state ? dirty_1_52 : _GEN_12897; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13927 = 3'h3 == state ? dirty_1_53 : _GEN_12898; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13928 = 3'h3 == state ? dirty_1_54 : _GEN_12899; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13929 = 3'h3 == state ? dirty_1_55 : _GEN_12900; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13930 = 3'h3 == state ? dirty_1_56 : _GEN_12901; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13931 = 3'h3 == state ? dirty_1_57 : _GEN_12902; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13932 = 3'h3 == state ? dirty_1_58 : _GEN_12903; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13933 = 3'h3 == state ? dirty_1_59 : _GEN_12904; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13934 = 3'h3 == state ? dirty_1_60 : _GEN_12905; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13935 = 3'h3 == state ? dirty_1_61 : _GEN_12906; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13936 = 3'h3 == state ? dirty_1_62 : _GEN_12907; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13937 = 3'h3 == state ? dirty_1_63 : _GEN_12908; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13938 = 3'h3 == state ? dirty_1_64 : _GEN_12909; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13939 = 3'h3 == state ? dirty_1_65 : _GEN_12910; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13940 = 3'h3 == state ? dirty_1_66 : _GEN_12911; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13941 = 3'h3 == state ? dirty_1_67 : _GEN_12912; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13942 = 3'h3 == state ? dirty_1_68 : _GEN_12913; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13943 = 3'h3 == state ? dirty_1_69 : _GEN_12914; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13944 = 3'h3 == state ? dirty_1_70 : _GEN_12915; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13945 = 3'h3 == state ? dirty_1_71 : _GEN_12916; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13946 = 3'h3 == state ? dirty_1_72 : _GEN_12917; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13947 = 3'h3 == state ? dirty_1_73 : _GEN_12918; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13948 = 3'h3 == state ? dirty_1_74 : _GEN_12919; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13949 = 3'h3 == state ? dirty_1_75 : _GEN_12920; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13950 = 3'h3 == state ? dirty_1_76 : _GEN_12921; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13951 = 3'h3 == state ? dirty_1_77 : _GEN_12922; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13952 = 3'h3 == state ? dirty_1_78 : _GEN_12923; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13953 = 3'h3 == state ? dirty_1_79 : _GEN_12924; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13954 = 3'h3 == state ? dirty_1_80 : _GEN_12925; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13955 = 3'h3 == state ? dirty_1_81 : _GEN_12926; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13956 = 3'h3 == state ? dirty_1_82 : _GEN_12927; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13957 = 3'h3 == state ? dirty_1_83 : _GEN_12928; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13958 = 3'h3 == state ? dirty_1_84 : _GEN_12929; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13959 = 3'h3 == state ? dirty_1_85 : _GEN_12930; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13960 = 3'h3 == state ? dirty_1_86 : _GEN_12931; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13961 = 3'h3 == state ? dirty_1_87 : _GEN_12932; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13962 = 3'h3 == state ? dirty_1_88 : _GEN_12933; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13963 = 3'h3 == state ? dirty_1_89 : _GEN_12934; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13964 = 3'h3 == state ? dirty_1_90 : _GEN_12935; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13965 = 3'h3 == state ? dirty_1_91 : _GEN_12936; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13966 = 3'h3 == state ? dirty_1_92 : _GEN_12937; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13967 = 3'h3 == state ? dirty_1_93 : _GEN_12938; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13968 = 3'h3 == state ? dirty_1_94 : _GEN_12939; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13969 = 3'h3 == state ? dirty_1_95 : _GEN_12940; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13970 = 3'h3 == state ? dirty_1_96 : _GEN_12941; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13971 = 3'h3 == state ? dirty_1_97 : _GEN_12942; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13972 = 3'h3 == state ? dirty_1_98 : _GEN_12943; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13973 = 3'h3 == state ? dirty_1_99 : _GEN_12944; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13974 = 3'h3 == state ? dirty_1_100 : _GEN_12945; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13975 = 3'h3 == state ? dirty_1_101 : _GEN_12946; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13976 = 3'h3 == state ? dirty_1_102 : _GEN_12947; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13977 = 3'h3 == state ? dirty_1_103 : _GEN_12948; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13978 = 3'h3 == state ? dirty_1_104 : _GEN_12949; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13979 = 3'h3 == state ? dirty_1_105 : _GEN_12950; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13980 = 3'h3 == state ? dirty_1_106 : _GEN_12951; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13981 = 3'h3 == state ? dirty_1_107 : _GEN_12952; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13982 = 3'h3 == state ? dirty_1_108 : _GEN_12953; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13983 = 3'h3 == state ? dirty_1_109 : _GEN_12954; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13984 = 3'h3 == state ? dirty_1_110 : _GEN_12955; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13985 = 3'h3 == state ? dirty_1_111 : _GEN_12956; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13986 = 3'h3 == state ? dirty_1_112 : _GEN_12957; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13987 = 3'h3 == state ? dirty_1_113 : _GEN_12958; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13988 = 3'h3 == state ? dirty_1_114 : _GEN_12959; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13989 = 3'h3 == state ? dirty_1_115 : _GEN_12960; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13990 = 3'h3 == state ? dirty_1_116 : _GEN_12961; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13991 = 3'h3 == state ? dirty_1_117 : _GEN_12962; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13992 = 3'h3 == state ? dirty_1_118 : _GEN_12963; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13993 = 3'h3 == state ? dirty_1_119 : _GEN_12964; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13994 = 3'h3 == state ? dirty_1_120 : _GEN_12965; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13995 = 3'h3 == state ? dirty_1_121 : _GEN_12966; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13996 = 3'h3 == state ? dirty_1_122 : _GEN_12967; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13997 = 3'h3 == state ? dirty_1_123 : _GEN_12968; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13998 = 3'h3 == state ? dirty_1_124 : _GEN_12969; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_13999 = 3'h3 == state ? dirty_1_125 : _GEN_12970; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_14000 = 3'h3 == state ? dirty_1_126 : _GEN_12971; // @[d_cache.scala 87:18 33:26]
  wire  _GEN_14001 = 3'h3 == state ? dirty_1_127 : _GEN_12972; // @[d_cache.scala 87:18 33:26]
  wire [41:0] _GEN_15670 = 3'h2 == state ? {{10'd0}, write_back_addr} : _GEN_13745; // @[d_cache.scala 87:18 38:34]
  wire [41:0] _GEN_17339 = 3'h1 == state ? {{10'd0}, write_back_addr} : _GEN_15670; // @[d_cache.scala 87:18 38:34]
  wire [41:0] _GEN_19008 = 3'h0 == state ? {{10'd0}, write_back_addr} : _GEN_17339; // @[d_cache.scala 87:18 38:34]
  wire [63:0] _io_to_lsu_rdata_T = _GEN_904 >> shift_bit; // @[d_cache.scala 237:49]
  wire [63:0] _io_to_lsu_rdata_T_1 = _GEN_1416 >> shift_bit; // @[d_cache.scala 244:49]
  wire [63:0] _GEN_19009 = way1_hit ? _io_to_lsu_rdata_T_1 : 64'h0; // @[d_cache.scala 243:33 244:33 251:33]
  wire [63:0] _GEN_19013 = way0_hit ? _io_to_lsu_rdata_T : _GEN_19009; // @[d_cache.scala 236:23 237:33]
  wire  _GEN_19015 = way0_hit | way1_hit; // @[d_cache.scala 236:23 239:34]
  wire  _GEN_19017 = way1_hit ? 1'h0 : 1'h1; // @[d_cache.scala 275:33 277:35 284:35]
  wire  _GEN_19018 = way0_hit ? 1'h0 : _GEN_19017; // @[d_cache.scala 268:23 270:35]
  wire  _T_34 = state == 3'h3; // @[d_cache.scala 290:21]
  wire [63:0] _GEN_20773 = {{32'd0}, io_from_lsu_araddr}; // @[d_cache.scala 298:48]
  wire [63:0] _io_to_axi_araddr_T = _GEN_20773 & 64'hfffffffffffffff8; // @[d_cache.scala 298:48]
  wire  _T_37 = state == 3'h6; // @[d_cache.scala 339:21]
  wire [31:0] _GEN_19021 = state == 3'h6 ? 32'h0 : io_from_lsu_araddr; // @[d_cache.scala 339:35 347:26 363:26]
  wire  _GEN_19022 = state == 3'h6 ? 1'h0 : io_from_lsu_rready; // @[d_cache.scala 339:35 348:26 364:26]
  wire [31:0] _GEN_19023 = state == 3'h6 ? write_back_addr : 32'h0; // @[d_cache.scala 339:35 349:26 365:26]
  wire [63:0] _GEN_19024 = state == 3'h6 ? write_back_data : 64'h0; // @[d_cache.scala 339:35 351:25 367:25]
  wire [7:0] _GEN_19025 = state == 3'h6 ? 8'hff : 8'h0; // @[d_cache.scala 339:35 352:25 368:25]
  wire  _GEN_19027 = state == 3'h5 | _T_37; // @[d_cache.scala 323:31 325:27]
  wire [31:0] _GEN_19028 = state == 3'h5 ? io_from_lsu_araddr : _GEN_19021; // @[d_cache.scala 323:31 331:26]
  wire  _GEN_19029 = state == 3'h5 ? io_from_lsu_rready : _GEN_19022; // @[d_cache.scala 323:31 332:26]
  wire [31:0] _GEN_19030 = state == 3'h5 ? 32'h0 : _GEN_19023; // @[d_cache.scala 323:31 333:26]
  wire  _GEN_19031 = state == 3'h5 ? 1'h0 : _T_37; // @[d_cache.scala 323:31 334:27]
  wire [63:0] _GEN_19032 = state == 3'h5 ? 64'h0 : _GEN_19024; // @[d_cache.scala 323:31 335:25]
  wire [7:0] _GEN_19033 = state == 3'h5 ? 8'h0 : _GEN_19025; // @[d_cache.scala 323:31 336:25]
  wire  _GEN_19035 = state == 3'h4 | _GEN_19027; // @[d_cache.scala 306:31 308:27]
  wire  _GEN_19036 = state == 3'h4 & io_from_axi_wready; // @[d_cache.scala 306:31 310:26]
  wire  _GEN_19037 = state == 3'h4 & io_from_axi_bvalid; // @[d_cache.scala 306:31 311:26]
  wire  _GEN_19038 = state == 3'h4 & io_from_axi_awready; // @[d_cache.scala 306:31 312:27]
  wire [31:0] _GEN_19039 = state == 3'h4 ? 32'h0 : _GEN_19028; // @[d_cache.scala 306:31 314:26]
  wire  _GEN_19040 = state == 3'h4 ? io_from_lsu_rready : _GEN_19029; // @[d_cache.scala 306:31 315:26]
  wire [31:0] _GEN_19041 = state == 3'h4 ? io_from_lsu_awaddr : _GEN_19030; // @[d_cache.scala 306:31 316:26]
  wire  _GEN_19042 = state == 3'h4 ? io_from_lsu_awvalid : _GEN_19031; // @[d_cache.scala 306:31 317:27]
  wire [63:0] _GEN_19043 = state == 3'h4 ? io_from_lsu_wdata : _GEN_19032; // @[d_cache.scala 306:31 318:25]
  wire [7:0] _GEN_19044 = state == 3'h4 ? io_from_lsu_wstrb : _GEN_19033; // @[d_cache.scala 306:31 319:25]
  wire  _GEN_19045 = state == 3'h4 ? io_from_lsu_wvalid : _GEN_19031; // @[d_cache.scala 306:31 320:26]
  wire  _GEN_19046 = state == 3'h4 ? io_from_lsu_bready : _GEN_19031; // @[d_cache.scala 306:31 321:26]
  wire  _GEN_19048 = state == 3'h3 | _GEN_19035; // @[d_cache.scala 290:31 292:27]
  wire  _GEN_19049 = state == 3'h3 ? 1'h0 : _GEN_19036; // @[d_cache.scala 290:31 294:26]
  wire  _GEN_19050 = state == 3'h3 ? 1'h0 : _GEN_19037; // @[d_cache.scala 290:31 295:26]
  wire  _GEN_19051 = state == 3'h3 ? 1'h0 : _GEN_19038; // @[d_cache.scala 290:31 296:27]
  wire [63:0] _GEN_19053 = state == 3'h3 ? _io_to_axi_araddr_T : {{32'd0}, _GEN_19039}; // @[d_cache.scala 290:31 298:26]
  wire  _GEN_19054 = state == 3'h3 ? io_from_lsu_rready : _GEN_19040; // @[d_cache.scala 290:31 299:26]
  wire [31:0] _GEN_19055 = state == 3'h3 ? 32'h0 : _GEN_19041; // @[d_cache.scala 290:31 300:26]
  wire  _GEN_19056 = state == 3'h3 ? 1'h0 : _GEN_19042; // @[d_cache.scala 290:31 301:27]
  wire [63:0] _GEN_19057 = state == 3'h3 ? 64'h0 : _GEN_19043; // @[d_cache.scala 290:31 302:25]
  wire [7:0] _GEN_19058 = state == 3'h3 ? 8'h0 : _GEN_19044; // @[d_cache.scala 290:31 303:25]
  wire  _GEN_19059 = state == 3'h3 ? 1'h0 : _GEN_19045; // @[d_cache.scala 290:31 304:26]
  wire  _GEN_19060 = state == 3'h3 ? 1'h0 : _GEN_19046; // @[d_cache.scala 290:31 305:26]
  wire  _GEN_19061 = state == 3'h2 ? 1'h0 : _T_34; // @[d_cache.scala 258:33 259:27]
  wire [63:0] _GEN_19062 = state == 3'h2 ? {{32'd0}, io_from_lsu_araddr} : _GEN_19053; // @[d_cache.scala 258:33 260:26]
  wire  _GEN_19063 = state == 3'h2 ? 1'h0 : _GEN_19054; // @[d_cache.scala 258:33 261:26]
  wire [31:0] _GEN_19064 = state == 3'h2 ? 32'h0 : _GEN_19055; // @[d_cache.scala 258:33 262:26]
  wire  _GEN_19065 = state == 3'h2 ? 1'h0 : _GEN_19056; // @[d_cache.scala 258:33 263:27]
  wire [63:0] _GEN_19066 = state == 3'h2 ? 64'h0 : _GEN_19057; // @[d_cache.scala 258:33 264:25]
  wire [7:0] _GEN_19067 = state == 3'h2 ? 8'h0 : _GEN_19058; // @[d_cache.scala 258:33 265:25]
  wire  _GEN_19068 = state == 3'h2 ? 1'h0 : _GEN_19059; // @[d_cache.scala 258:33 266:26]
  wire  _GEN_19069 = state == 3'h2 ? 1'h0 : _GEN_19060; // @[d_cache.scala 258:33 267:26]
  wire  _GEN_19071 = state == 3'h2 ? _GEN_19018 : _GEN_19048; // @[d_cache.scala 258:33]
  wire  _GEN_19072 = state == 3'h2 ? _GEN_19015 : _GEN_19049; // @[d_cache.scala 258:33]
  wire  _GEN_19073 = state == 3'h2 ? _GEN_19015 : _GEN_19051; // @[d_cache.scala 258:33]
  wire  _GEN_19074 = state == 3'h2 ? _GEN_19015 : _GEN_19050; // @[d_cache.scala 258:33]
  wire  _GEN_19075 = state == 3'h1 ? 1'h0 : _GEN_19061; // @[d_cache.scala 226:33 227:27]
  wire [63:0] _GEN_19076 = state == 3'h1 ? {{32'd0}, io_from_lsu_araddr} : _GEN_19062; // @[d_cache.scala 226:33 228:26]
  wire  _GEN_19077 = state == 3'h1 ? io_from_lsu_rready : _GEN_19063; // @[d_cache.scala 226:33 229:26]
  wire [31:0] _GEN_19078 = state == 3'h1 ? 32'h0 : _GEN_19064; // @[d_cache.scala 226:33 230:26]
  wire  _GEN_19079 = state == 3'h1 ? 1'h0 : _GEN_19065; // @[d_cache.scala 226:33 231:27]
  wire [63:0] _GEN_19080 = state == 3'h1 ? 64'h0 : _GEN_19066; // @[d_cache.scala 226:33 232:25]
  wire [7:0] _GEN_19081 = state == 3'h1 ? 8'h0 : _GEN_19067; // @[d_cache.scala 226:33 233:25]
  wire  _GEN_19082 = state == 3'h1 ? 1'h0 : _GEN_19068; // @[d_cache.scala 226:33 234:26]
  wire  _GEN_19083 = state == 3'h1 ? io_from_lsu_bready : _GEN_19069; // @[d_cache.scala 226:33 235:26]
  wire [63:0] _GEN_19084 = state == 3'h1 ? _GEN_19013 : 64'h0; // @[d_cache.scala 226:33]
  wire  _GEN_19085 = state == 3'h1 | _GEN_19071; // @[d_cache.scala 226:33]
  wire  _GEN_19086 = state == 3'h1 & _GEN_19015; // @[d_cache.scala 226:33]
  wire  _GEN_19087 = state == 3'h1 ? 1'h0 : _GEN_19072; // @[d_cache.scala 226:33]
  wire  _GEN_19088 = state == 3'h1 ? 1'h0 : _GEN_19073; // @[d_cache.scala 226:33]
  wire  _GEN_19089 = state == 3'h1 ? 1'h0 : _GEN_19074; // @[d_cache.scala 226:33]
  wire [63:0] _GEN_19097 = state == 3'h0 ? {{32'd0}, io_from_lsu_araddr} : _GEN_19076; // @[d_cache.scala 210:23 218:26]
  wire [63:0] _GEN_19106 = 7'h1 == index ? record_wdata1_1 : record_wdata1_0; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19107 = 7'h2 == index ? record_wdata1_2 : _GEN_19106; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19108 = 7'h3 == index ? record_wdata1_3 : _GEN_19107; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19109 = 7'h4 == index ? record_wdata1_4 : _GEN_19108; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19110 = 7'h5 == index ? record_wdata1_5 : _GEN_19109; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19111 = 7'h6 == index ? record_wdata1_6 : _GEN_19110; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19112 = 7'h7 == index ? record_wdata1_7 : _GEN_19111; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19113 = 7'h8 == index ? record_wdata1_8 : _GEN_19112; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19114 = 7'h9 == index ? record_wdata1_9 : _GEN_19113; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19115 = 7'ha == index ? record_wdata1_10 : _GEN_19114; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19116 = 7'hb == index ? record_wdata1_11 : _GEN_19115; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19117 = 7'hc == index ? record_wdata1_12 : _GEN_19116; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19118 = 7'hd == index ? record_wdata1_13 : _GEN_19117; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19119 = 7'he == index ? record_wdata1_14 : _GEN_19118; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19120 = 7'hf == index ? record_wdata1_15 : _GEN_19119; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19121 = 7'h10 == index ? record_wdata1_16 : _GEN_19120; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19122 = 7'h11 == index ? record_wdata1_17 : _GEN_19121; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19123 = 7'h12 == index ? record_wdata1_18 : _GEN_19122; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19124 = 7'h13 == index ? record_wdata1_19 : _GEN_19123; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19125 = 7'h14 == index ? record_wdata1_20 : _GEN_19124; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19126 = 7'h15 == index ? record_wdata1_21 : _GEN_19125; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19127 = 7'h16 == index ? record_wdata1_22 : _GEN_19126; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19128 = 7'h17 == index ? record_wdata1_23 : _GEN_19127; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19129 = 7'h18 == index ? record_wdata1_24 : _GEN_19128; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19130 = 7'h19 == index ? record_wdata1_25 : _GEN_19129; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19131 = 7'h1a == index ? record_wdata1_26 : _GEN_19130; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19132 = 7'h1b == index ? record_wdata1_27 : _GEN_19131; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19133 = 7'h1c == index ? record_wdata1_28 : _GEN_19132; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19134 = 7'h1d == index ? record_wdata1_29 : _GEN_19133; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19135 = 7'h1e == index ? record_wdata1_30 : _GEN_19134; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19136 = 7'h1f == index ? record_wdata1_31 : _GEN_19135; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19137 = 7'h20 == index ? record_wdata1_32 : _GEN_19136; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19138 = 7'h21 == index ? record_wdata1_33 : _GEN_19137; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19139 = 7'h22 == index ? record_wdata1_34 : _GEN_19138; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19140 = 7'h23 == index ? record_wdata1_35 : _GEN_19139; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19141 = 7'h24 == index ? record_wdata1_36 : _GEN_19140; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19142 = 7'h25 == index ? record_wdata1_37 : _GEN_19141; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19143 = 7'h26 == index ? record_wdata1_38 : _GEN_19142; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19144 = 7'h27 == index ? record_wdata1_39 : _GEN_19143; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19145 = 7'h28 == index ? record_wdata1_40 : _GEN_19144; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19146 = 7'h29 == index ? record_wdata1_41 : _GEN_19145; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19147 = 7'h2a == index ? record_wdata1_42 : _GEN_19146; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19148 = 7'h2b == index ? record_wdata1_43 : _GEN_19147; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19149 = 7'h2c == index ? record_wdata1_44 : _GEN_19148; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19150 = 7'h2d == index ? record_wdata1_45 : _GEN_19149; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19151 = 7'h2e == index ? record_wdata1_46 : _GEN_19150; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19152 = 7'h2f == index ? record_wdata1_47 : _GEN_19151; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19153 = 7'h30 == index ? record_wdata1_48 : _GEN_19152; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19154 = 7'h31 == index ? record_wdata1_49 : _GEN_19153; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19155 = 7'h32 == index ? record_wdata1_50 : _GEN_19154; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19156 = 7'h33 == index ? record_wdata1_51 : _GEN_19155; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19157 = 7'h34 == index ? record_wdata1_52 : _GEN_19156; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19158 = 7'h35 == index ? record_wdata1_53 : _GEN_19157; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19159 = 7'h36 == index ? record_wdata1_54 : _GEN_19158; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19160 = 7'h37 == index ? record_wdata1_55 : _GEN_19159; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19161 = 7'h38 == index ? record_wdata1_56 : _GEN_19160; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19162 = 7'h39 == index ? record_wdata1_57 : _GEN_19161; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19163 = 7'h3a == index ? record_wdata1_58 : _GEN_19162; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19164 = 7'h3b == index ? record_wdata1_59 : _GEN_19163; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19165 = 7'h3c == index ? record_wdata1_60 : _GEN_19164; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19166 = 7'h3d == index ? record_wdata1_61 : _GEN_19165; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19167 = 7'h3e == index ? record_wdata1_62 : _GEN_19166; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19168 = 7'h3f == index ? record_wdata1_63 : _GEN_19167; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19169 = 7'h40 == index ? record_wdata1_64 : _GEN_19168; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19170 = 7'h41 == index ? record_wdata1_65 : _GEN_19169; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19171 = 7'h42 == index ? record_wdata1_66 : _GEN_19170; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19172 = 7'h43 == index ? record_wdata1_67 : _GEN_19171; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19173 = 7'h44 == index ? record_wdata1_68 : _GEN_19172; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19174 = 7'h45 == index ? record_wdata1_69 : _GEN_19173; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19175 = 7'h46 == index ? record_wdata1_70 : _GEN_19174; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19176 = 7'h47 == index ? record_wdata1_71 : _GEN_19175; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19177 = 7'h48 == index ? record_wdata1_72 : _GEN_19176; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19178 = 7'h49 == index ? record_wdata1_73 : _GEN_19177; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19179 = 7'h4a == index ? record_wdata1_74 : _GEN_19178; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19180 = 7'h4b == index ? record_wdata1_75 : _GEN_19179; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19181 = 7'h4c == index ? record_wdata1_76 : _GEN_19180; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19182 = 7'h4d == index ? record_wdata1_77 : _GEN_19181; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19183 = 7'h4e == index ? record_wdata1_78 : _GEN_19182; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19184 = 7'h4f == index ? record_wdata1_79 : _GEN_19183; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19185 = 7'h50 == index ? record_wdata1_80 : _GEN_19184; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19186 = 7'h51 == index ? record_wdata1_81 : _GEN_19185; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19187 = 7'h52 == index ? record_wdata1_82 : _GEN_19186; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19188 = 7'h53 == index ? record_wdata1_83 : _GEN_19187; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19189 = 7'h54 == index ? record_wdata1_84 : _GEN_19188; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19190 = 7'h55 == index ? record_wdata1_85 : _GEN_19189; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19191 = 7'h56 == index ? record_wdata1_86 : _GEN_19190; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19192 = 7'h57 == index ? record_wdata1_87 : _GEN_19191; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19193 = 7'h58 == index ? record_wdata1_88 : _GEN_19192; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19194 = 7'h59 == index ? record_wdata1_89 : _GEN_19193; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19195 = 7'h5a == index ? record_wdata1_90 : _GEN_19194; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19196 = 7'h5b == index ? record_wdata1_91 : _GEN_19195; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19197 = 7'h5c == index ? record_wdata1_92 : _GEN_19196; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19198 = 7'h5d == index ? record_wdata1_93 : _GEN_19197; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19199 = 7'h5e == index ? record_wdata1_94 : _GEN_19198; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19200 = 7'h5f == index ? record_wdata1_95 : _GEN_19199; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19201 = 7'h60 == index ? record_wdata1_96 : _GEN_19200; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19202 = 7'h61 == index ? record_wdata1_97 : _GEN_19201; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19203 = 7'h62 == index ? record_wdata1_98 : _GEN_19202; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19204 = 7'h63 == index ? record_wdata1_99 : _GEN_19203; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19205 = 7'h64 == index ? record_wdata1_100 : _GEN_19204; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19206 = 7'h65 == index ? record_wdata1_101 : _GEN_19205; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19207 = 7'h66 == index ? record_wdata1_102 : _GEN_19206; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19208 = 7'h67 == index ? record_wdata1_103 : _GEN_19207; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19209 = 7'h68 == index ? record_wdata1_104 : _GEN_19208; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19210 = 7'h69 == index ? record_wdata1_105 : _GEN_19209; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19211 = 7'h6a == index ? record_wdata1_106 : _GEN_19210; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19212 = 7'h6b == index ? record_wdata1_107 : _GEN_19211; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19213 = 7'h6c == index ? record_wdata1_108 : _GEN_19212; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19214 = 7'h6d == index ? record_wdata1_109 : _GEN_19213; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19215 = 7'h6e == index ? record_wdata1_110 : _GEN_19214; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19216 = 7'h6f == index ? record_wdata1_111 : _GEN_19215; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19217 = 7'h70 == index ? record_wdata1_112 : _GEN_19216; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19218 = 7'h71 == index ? record_wdata1_113 : _GEN_19217; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19219 = 7'h72 == index ? record_wdata1_114 : _GEN_19218; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19220 = 7'h73 == index ? record_wdata1_115 : _GEN_19219; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19221 = 7'h74 == index ? record_wdata1_116 : _GEN_19220; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19222 = 7'h75 == index ? record_wdata1_117 : _GEN_19221; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19223 = 7'h76 == index ? record_wdata1_118 : _GEN_19222; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19224 = 7'h77 == index ? record_wdata1_119 : _GEN_19223; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19225 = 7'h78 == index ? record_wdata1_120 : _GEN_19224; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19226 = 7'h79 == index ? record_wdata1_121 : _GEN_19225; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19227 = 7'h7a == index ? record_wdata1_122 : _GEN_19226; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19228 = 7'h7b == index ? record_wdata1_123 : _GEN_19227; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19229 = 7'h7c == index ? record_wdata1_124 : _GEN_19228; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19230 = 7'h7d == index ? record_wdata1_125 : _GEN_19229; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19231 = 7'h7e == index ? record_wdata1_126 : _GEN_19230; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19234 = 7'h1 == index ? record_wstrb1_1 : record_wstrb1_0; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19235 = 7'h2 == index ? record_wstrb1_2 : _GEN_19234; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19236 = 7'h3 == index ? record_wstrb1_3 : _GEN_19235; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19237 = 7'h4 == index ? record_wstrb1_4 : _GEN_19236; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19238 = 7'h5 == index ? record_wstrb1_5 : _GEN_19237; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19239 = 7'h6 == index ? record_wstrb1_6 : _GEN_19238; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19240 = 7'h7 == index ? record_wstrb1_7 : _GEN_19239; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19241 = 7'h8 == index ? record_wstrb1_8 : _GEN_19240; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19242 = 7'h9 == index ? record_wstrb1_9 : _GEN_19241; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19243 = 7'ha == index ? record_wstrb1_10 : _GEN_19242; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19244 = 7'hb == index ? record_wstrb1_11 : _GEN_19243; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19245 = 7'hc == index ? record_wstrb1_12 : _GEN_19244; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19246 = 7'hd == index ? record_wstrb1_13 : _GEN_19245; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19247 = 7'he == index ? record_wstrb1_14 : _GEN_19246; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19248 = 7'hf == index ? record_wstrb1_15 : _GEN_19247; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19249 = 7'h10 == index ? record_wstrb1_16 : _GEN_19248; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19250 = 7'h11 == index ? record_wstrb1_17 : _GEN_19249; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19251 = 7'h12 == index ? record_wstrb1_18 : _GEN_19250; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19252 = 7'h13 == index ? record_wstrb1_19 : _GEN_19251; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19253 = 7'h14 == index ? record_wstrb1_20 : _GEN_19252; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19254 = 7'h15 == index ? record_wstrb1_21 : _GEN_19253; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19255 = 7'h16 == index ? record_wstrb1_22 : _GEN_19254; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19256 = 7'h17 == index ? record_wstrb1_23 : _GEN_19255; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19257 = 7'h18 == index ? record_wstrb1_24 : _GEN_19256; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19258 = 7'h19 == index ? record_wstrb1_25 : _GEN_19257; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19259 = 7'h1a == index ? record_wstrb1_26 : _GEN_19258; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19260 = 7'h1b == index ? record_wstrb1_27 : _GEN_19259; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19261 = 7'h1c == index ? record_wstrb1_28 : _GEN_19260; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19262 = 7'h1d == index ? record_wstrb1_29 : _GEN_19261; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19263 = 7'h1e == index ? record_wstrb1_30 : _GEN_19262; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19264 = 7'h1f == index ? record_wstrb1_31 : _GEN_19263; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19265 = 7'h20 == index ? record_wstrb1_32 : _GEN_19264; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19266 = 7'h21 == index ? record_wstrb1_33 : _GEN_19265; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19267 = 7'h22 == index ? record_wstrb1_34 : _GEN_19266; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19268 = 7'h23 == index ? record_wstrb1_35 : _GEN_19267; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19269 = 7'h24 == index ? record_wstrb1_36 : _GEN_19268; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19270 = 7'h25 == index ? record_wstrb1_37 : _GEN_19269; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19271 = 7'h26 == index ? record_wstrb1_38 : _GEN_19270; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19272 = 7'h27 == index ? record_wstrb1_39 : _GEN_19271; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19273 = 7'h28 == index ? record_wstrb1_40 : _GEN_19272; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19274 = 7'h29 == index ? record_wstrb1_41 : _GEN_19273; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19275 = 7'h2a == index ? record_wstrb1_42 : _GEN_19274; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19276 = 7'h2b == index ? record_wstrb1_43 : _GEN_19275; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19277 = 7'h2c == index ? record_wstrb1_44 : _GEN_19276; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19278 = 7'h2d == index ? record_wstrb1_45 : _GEN_19277; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19279 = 7'h2e == index ? record_wstrb1_46 : _GEN_19278; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19280 = 7'h2f == index ? record_wstrb1_47 : _GEN_19279; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19281 = 7'h30 == index ? record_wstrb1_48 : _GEN_19280; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19282 = 7'h31 == index ? record_wstrb1_49 : _GEN_19281; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19283 = 7'h32 == index ? record_wstrb1_50 : _GEN_19282; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19284 = 7'h33 == index ? record_wstrb1_51 : _GEN_19283; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19285 = 7'h34 == index ? record_wstrb1_52 : _GEN_19284; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19286 = 7'h35 == index ? record_wstrb1_53 : _GEN_19285; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19287 = 7'h36 == index ? record_wstrb1_54 : _GEN_19286; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19288 = 7'h37 == index ? record_wstrb1_55 : _GEN_19287; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19289 = 7'h38 == index ? record_wstrb1_56 : _GEN_19288; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19290 = 7'h39 == index ? record_wstrb1_57 : _GEN_19289; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19291 = 7'h3a == index ? record_wstrb1_58 : _GEN_19290; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19292 = 7'h3b == index ? record_wstrb1_59 : _GEN_19291; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19293 = 7'h3c == index ? record_wstrb1_60 : _GEN_19292; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19294 = 7'h3d == index ? record_wstrb1_61 : _GEN_19293; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19295 = 7'h3e == index ? record_wstrb1_62 : _GEN_19294; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19296 = 7'h3f == index ? record_wstrb1_63 : _GEN_19295; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19297 = 7'h40 == index ? record_wstrb1_64 : _GEN_19296; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19298 = 7'h41 == index ? record_wstrb1_65 : _GEN_19297; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19299 = 7'h42 == index ? record_wstrb1_66 : _GEN_19298; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19300 = 7'h43 == index ? record_wstrb1_67 : _GEN_19299; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19301 = 7'h44 == index ? record_wstrb1_68 : _GEN_19300; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19302 = 7'h45 == index ? record_wstrb1_69 : _GEN_19301; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19303 = 7'h46 == index ? record_wstrb1_70 : _GEN_19302; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19304 = 7'h47 == index ? record_wstrb1_71 : _GEN_19303; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19305 = 7'h48 == index ? record_wstrb1_72 : _GEN_19304; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19306 = 7'h49 == index ? record_wstrb1_73 : _GEN_19305; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19307 = 7'h4a == index ? record_wstrb1_74 : _GEN_19306; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19308 = 7'h4b == index ? record_wstrb1_75 : _GEN_19307; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19309 = 7'h4c == index ? record_wstrb1_76 : _GEN_19308; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19310 = 7'h4d == index ? record_wstrb1_77 : _GEN_19309; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19311 = 7'h4e == index ? record_wstrb1_78 : _GEN_19310; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19312 = 7'h4f == index ? record_wstrb1_79 : _GEN_19311; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19313 = 7'h50 == index ? record_wstrb1_80 : _GEN_19312; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19314 = 7'h51 == index ? record_wstrb1_81 : _GEN_19313; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19315 = 7'h52 == index ? record_wstrb1_82 : _GEN_19314; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19316 = 7'h53 == index ? record_wstrb1_83 : _GEN_19315; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19317 = 7'h54 == index ? record_wstrb1_84 : _GEN_19316; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19318 = 7'h55 == index ? record_wstrb1_85 : _GEN_19317; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19319 = 7'h56 == index ? record_wstrb1_86 : _GEN_19318; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19320 = 7'h57 == index ? record_wstrb1_87 : _GEN_19319; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19321 = 7'h58 == index ? record_wstrb1_88 : _GEN_19320; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19322 = 7'h59 == index ? record_wstrb1_89 : _GEN_19321; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19323 = 7'h5a == index ? record_wstrb1_90 : _GEN_19322; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19324 = 7'h5b == index ? record_wstrb1_91 : _GEN_19323; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19325 = 7'h5c == index ? record_wstrb1_92 : _GEN_19324; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19326 = 7'h5d == index ? record_wstrb1_93 : _GEN_19325; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19327 = 7'h5e == index ? record_wstrb1_94 : _GEN_19326; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19328 = 7'h5f == index ? record_wstrb1_95 : _GEN_19327; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19329 = 7'h60 == index ? record_wstrb1_96 : _GEN_19328; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19330 = 7'h61 == index ? record_wstrb1_97 : _GEN_19329; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19331 = 7'h62 == index ? record_wstrb1_98 : _GEN_19330; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19332 = 7'h63 == index ? record_wstrb1_99 : _GEN_19331; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19333 = 7'h64 == index ? record_wstrb1_100 : _GEN_19332; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19334 = 7'h65 == index ? record_wstrb1_101 : _GEN_19333; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19335 = 7'h66 == index ? record_wstrb1_102 : _GEN_19334; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19336 = 7'h67 == index ? record_wstrb1_103 : _GEN_19335; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19337 = 7'h68 == index ? record_wstrb1_104 : _GEN_19336; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19338 = 7'h69 == index ? record_wstrb1_105 : _GEN_19337; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19339 = 7'h6a == index ? record_wstrb1_106 : _GEN_19338; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19340 = 7'h6b == index ? record_wstrb1_107 : _GEN_19339; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19341 = 7'h6c == index ? record_wstrb1_108 : _GEN_19340; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19342 = 7'h6d == index ? record_wstrb1_109 : _GEN_19341; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19343 = 7'h6e == index ? record_wstrb1_110 : _GEN_19342; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19344 = 7'h6f == index ? record_wstrb1_111 : _GEN_19343; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19345 = 7'h70 == index ? record_wstrb1_112 : _GEN_19344; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19346 = 7'h71 == index ? record_wstrb1_113 : _GEN_19345; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19347 = 7'h72 == index ? record_wstrb1_114 : _GEN_19346; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19348 = 7'h73 == index ? record_wstrb1_115 : _GEN_19347; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19349 = 7'h74 == index ? record_wstrb1_116 : _GEN_19348; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19350 = 7'h75 == index ? record_wstrb1_117 : _GEN_19349; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19351 = 7'h76 == index ? record_wstrb1_118 : _GEN_19350; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19352 = 7'h77 == index ? record_wstrb1_119 : _GEN_19351; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19353 = 7'h78 == index ? record_wstrb1_120 : _GEN_19352; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19354 = 7'h79 == index ? record_wstrb1_121 : _GEN_19353; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19355 = 7'h7a == index ? record_wstrb1_122 : _GEN_19354; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19356 = 7'h7b == index ? record_wstrb1_123 : _GEN_19355; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19357 = 7'h7c == index ? record_wstrb1_124 : _GEN_19356; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19358 = 7'h7d == index ? record_wstrb1_125 : _GEN_19357; // @[d_cache.scala 374:{11,11}]
  wire [7:0] _GEN_19359 = 7'h7e == index ? record_wstrb1_126 : _GEN_19358; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19362 = 7'h1 == index ? record_pc_1 : record_pc_0; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19363 = 7'h2 == index ? record_pc_2 : _GEN_19362; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19364 = 7'h3 == index ? record_pc_3 : _GEN_19363; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19365 = 7'h4 == index ? record_pc_4 : _GEN_19364; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19366 = 7'h5 == index ? record_pc_5 : _GEN_19365; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19367 = 7'h6 == index ? record_pc_6 : _GEN_19366; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19368 = 7'h7 == index ? record_pc_7 : _GEN_19367; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19369 = 7'h8 == index ? record_pc_8 : _GEN_19368; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19370 = 7'h9 == index ? record_pc_9 : _GEN_19369; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19371 = 7'ha == index ? record_pc_10 : _GEN_19370; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19372 = 7'hb == index ? record_pc_11 : _GEN_19371; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19373 = 7'hc == index ? record_pc_12 : _GEN_19372; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19374 = 7'hd == index ? record_pc_13 : _GEN_19373; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19375 = 7'he == index ? record_pc_14 : _GEN_19374; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19376 = 7'hf == index ? record_pc_15 : _GEN_19375; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19377 = 7'h10 == index ? record_pc_16 : _GEN_19376; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19378 = 7'h11 == index ? record_pc_17 : _GEN_19377; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19379 = 7'h12 == index ? record_pc_18 : _GEN_19378; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19380 = 7'h13 == index ? record_pc_19 : _GEN_19379; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19381 = 7'h14 == index ? record_pc_20 : _GEN_19380; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19382 = 7'h15 == index ? record_pc_21 : _GEN_19381; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19383 = 7'h16 == index ? record_pc_22 : _GEN_19382; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19384 = 7'h17 == index ? record_pc_23 : _GEN_19383; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19385 = 7'h18 == index ? record_pc_24 : _GEN_19384; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19386 = 7'h19 == index ? record_pc_25 : _GEN_19385; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19387 = 7'h1a == index ? record_pc_26 : _GEN_19386; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19388 = 7'h1b == index ? record_pc_27 : _GEN_19387; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19389 = 7'h1c == index ? record_pc_28 : _GEN_19388; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19390 = 7'h1d == index ? record_pc_29 : _GEN_19389; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19391 = 7'h1e == index ? record_pc_30 : _GEN_19390; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19392 = 7'h1f == index ? record_pc_31 : _GEN_19391; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19393 = 7'h20 == index ? record_pc_32 : _GEN_19392; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19394 = 7'h21 == index ? record_pc_33 : _GEN_19393; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19395 = 7'h22 == index ? record_pc_34 : _GEN_19394; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19396 = 7'h23 == index ? record_pc_35 : _GEN_19395; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19397 = 7'h24 == index ? record_pc_36 : _GEN_19396; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19398 = 7'h25 == index ? record_pc_37 : _GEN_19397; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19399 = 7'h26 == index ? record_pc_38 : _GEN_19398; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19400 = 7'h27 == index ? record_pc_39 : _GEN_19399; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19401 = 7'h28 == index ? record_pc_40 : _GEN_19400; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19402 = 7'h29 == index ? record_pc_41 : _GEN_19401; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19403 = 7'h2a == index ? record_pc_42 : _GEN_19402; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19404 = 7'h2b == index ? record_pc_43 : _GEN_19403; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19405 = 7'h2c == index ? record_pc_44 : _GEN_19404; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19406 = 7'h2d == index ? record_pc_45 : _GEN_19405; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19407 = 7'h2e == index ? record_pc_46 : _GEN_19406; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19408 = 7'h2f == index ? record_pc_47 : _GEN_19407; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19409 = 7'h30 == index ? record_pc_48 : _GEN_19408; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19410 = 7'h31 == index ? record_pc_49 : _GEN_19409; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19411 = 7'h32 == index ? record_pc_50 : _GEN_19410; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19412 = 7'h33 == index ? record_pc_51 : _GEN_19411; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19413 = 7'h34 == index ? record_pc_52 : _GEN_19412; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19414 = 7'h35 == index ? record_pc_53 : _GEN_19413; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19415 = 7'h36 == index ? record_pc_54 : _GEN_19414; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19416 = 7'h37 == index ? record_pc_55 : _GEN_19415; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19417 = 7'h38 == index ? record_pc_56 : _GEN_19416; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19418 = 7'h39 == index ? record_pc_57 : _GEN_19417; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19419 = 7'h3a == index ? record_pc_58 : _GEN_19418; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19420 = 7'h3b == index ? record_pc_59 : _GEN_19419; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19421 = 7'h3c == index ? record_pc_60 : _GEN_19420; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19422 = 7'h3d == index ? record_pc_61 : _GEN_19421; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19423 = 7'h3e == index ? record_pc_62 : _GEN_19422; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19424 = 7'h3f == index ? record_pc_63 : _GEN_19423; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19425 = 7'h40 == index ? record_pc_64 : _GEN_19424; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19426 = 7'h41 == index ? record_pc_65 : _GEN_19425; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19427 = 7'h42 == index ? record_pc_66 : _GEN_19426; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19428 = 7'h43 == index ? record_pc_67 : _GEN_19427; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19429 = 7'h44 == index ? record_pc_68 : _GEN_19428; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19430 = 7'h45 == index ? record_pc_69 : _GEN_19429; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19431 = 7'h46 == index ? record_pc_70 : _GEN_19430; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19432 = 7'h47 == index ? record_pc_71 : _GEN_19431; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19433 = 7'h48 == index ? record_pc_72 : _GEN_19432; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19434 = 7'h49 == index ? record_pc_73 : _GEN_19433; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19435 = 7'h4a == index ? record_pc_74 : _GEN_19434; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19436 = 7'h4b == index ? record_pc_75 : _GEN_19435; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19437 = 7'h4c == index ? record_pc_76 : _GEN_19436; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19438 = 7'h4d == index ? record_pc_77 : _GEN_19437; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19439 = 7'h4e == index ? record_pc_78 : _GEN_19438; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19440 = 7'h4f == index ? record_pc_79 : _GEN_19439; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19441 = 7'h50 == index ? record_pc_80 : _GEN_19440; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19442 = 7'h51 == index ? record_pc_81 : _GEN_19441; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19443 = 7'h52 == index ? record_pc_82 : _GEN_19442; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19444 = 7'h53 == index ? record_pc_83 : _GEN_19443; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19445 = 7'h54 == index ? record_pc_84 : _GEN_19444; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19446 = 7'h55 == index ? record_pc_85 : _GEN_19445; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19447 = 7'h56 == index ? record_pc_86 : _GEN_19446; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19448 = 7'h57 == index ? record_pc_87 : _GEN_19447; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19449 = 7'h58 == index ? record_pc_88 : _GEN_19448; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19450 = 7'h59 == index ? record_pc_89 : _GEN_19449; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19451 = 7'h5a == index ? record_pc_90 : _GEN_19450; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19452 = 7'h5b == index ? record_pc_91 : _GEN_19451; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19453 = 7'h5c == index ? record_pc_92 : _GEN_19452; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19454 = 7'h5d == index ? record_pc_93 : _GEN_19453; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19455 = 7'h5e == index ? record_pc_94 : _GEN_19454; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19456 = 7'h5f == index ? record_pc_95 : _GEN_19455; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19457 = 7'h60 == index ? record_pc_96 : _GEN_19456; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19458 = 7'h61 == index ? record_pc_97 : _GEN_19457; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19459 = 7'h62 == index ? record_pc_98 : _GEN_19458; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19460 = 7'h63 == index ? record_pc_99 : _GEN_19459; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19461 = 7'h64 == index ? record_pc_100 : _GEN_19460; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19462 = 7'h65 == index ? record_pc_101 : _GEN_19461; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19463 = 7'h66 == index ? record_pc_102 : _GEN_19462; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19464 = 7'h67 == index ? record_pc_103 : _GEN_19463; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19465 = 7'h68 == index ? record_pc_104 : _GEN_19464; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19466 = 7'h69 == index ? record_pc_105 : _GEN_19465; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19467 = 7'h6a == index ? record_pc_106 : _GEN_19466; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19468 = 7'h6b == index ? record_pc_107 : _GEN_19467; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19469 = 7'h6c == index ? record_pc_108 : _GEN_19468; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19470 = 7'h6d == index ? record_pc_109 : _GEN_19469; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19471 = 7'h6e == index ? record_pc_110 : _GEN_19470; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19472 = 7'h6f == index ? record_pc_111 : _GEN_19471; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19473 = 7'h70 == index ? record_pc_112 : _GEN_19472; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19474 = 7'h71 == index ? record_pc_113 : _GEN_19473; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19475 = 7'h72 == index ? record_pc_114 : _GEN_19474; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19476 = 7'h73 == index ? record_pc_115 : _GEN_19475; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19477 = 7'h74 == index ? record_pc_116 : _GEN_19476; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19478 = 7'h75 == index ? record_pc_117 : _GEN_19477; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19479 = 7'h76 == index ? record_pc_118 : _GEN_19478; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19480 = 7'h77 == index ? record_pc_119 : _GEN_19479; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19481 = 7'h78 == index ? record_pc_120 : _GEN_19480; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19482 = 7'h79 == index ? record_pc_121 : _GEN_19481; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19483 = 7'h7a == index ? record_pc_122 : _GEN_19482; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19484 = 7'h7b == index ? record_pc_123 : _GEN_19483; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19485 = 7'h7c == index ? record_pc_124 : _GEN_19484; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19486 = 7'h7d == index ? record_pc_125 : _GEN_19485; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19487 = 7'h7e == index ? record_pc_126 : _GEN_19486; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19490 = 7'h1 == index ? record_addr_1 : record_addr_0; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19491 = 7'h2 == index ? record_addr_2 : _GEN_19490; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19492 = 7'h3 == index ? record_addr_3 : _GEN_19491; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19493 = 7'h4 == index ? record_addr_4 : _GEN_19492; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19494 = 7'h5 == index ? record_addr_5 : _GEN_19493; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19495 = 7'h6 == index ? record_addr_6 : _GEN_19494; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19496 = 7'h7 == index ? record_addr_7 : _GEN_19495; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19497 = 7'h8 == index ? record_addr_8 : _GEN_19496; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19498 = 7'h9 == index ? record_addr_9 : _GEN_19497; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19499 = 7'ha == index ? record_addr_10 : _GEN_19498; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19500 = 7'hb == index ? record_addr_11 : _GEN_19499; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19501 = 7'hc == index ? record_addr_12 : _GEN_19500; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19502 = 7'hd == index ? record_addr_13 : _GEN_19501; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19503 = 7'he == index ? record_addr_14 : _GEN_19502; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19504 = 7'hf == index ? record_addr_15 : _GEN_19503; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19505 = 7'h10 == index ? record_addr_16 : _GEN_19504; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19506 = 7'h11 == index ? record_addr_17 : _GEN_19505; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19507 = 7'h12 == index ? record_addr_18 : _GEN_19506; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19508 = 7'h13 == index ? record_addr_19 : _GEN_19507; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19509 = 7'h14 == index ? record_addr_20 : _GEN_19508; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19510 = 7'h15 == index ? record_addr_21 : _GEN_19509; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19511 = 7'h16 == index ? record_addr_22 : _GEN_19510; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19512 = 7'h17 == index ? record_addr_23 : _GEN_19511; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19513 = 7'h18 == index ? record_addr_24 : _GEN_19512; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19514 = 7'h19 == index ? record_addr_25 : _GEN_19513; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19515 = 7'h1a == index ? record_addr_26 : _GEN_19514; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19516 = 7'h1b == index ? record_addr_27 : _GEN_19515; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19517 = 7'h1c == index ? record_addr_28 : _GEN_19516; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19518 = 7'h1d == index ? record_addr_29 : _GEN_19517; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19519 = 7'h1e == index ? record_addr_30 : _GEN_19518; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19520 = 7'h1f == index ? record_addr_31 : _GEN_19519; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19521 = 7'h20 == index ? record_addr_32 : _GEN_19520; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19522 = 7'h21 == index ? record_addr_33 : _GEN_19521; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19523 = 7'h22 == index ? record_addr_34 : _GEN_19522; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19524 = 7'h23 == index ? record_addr_35 : _GEN_19523; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19525 = 7'h24 == index ? record_addr_36 : _GEN_19524; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19526 = 7'h25 == index ? record_addr_37 : _GEN_19525; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19527 = 7'h26 == index ? record_addr_38 : _GEN_19526; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19528 = 7'h27 == index ? record_addr_39 : _GEN_19527; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19529 = 7'h28 == index ? record_addr_40 : _GEN_19528; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19530 = 7'h29 == index ? record_addr_41 : _GEN_19529; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19531 = 7'h2a == index ? record_addr_42 : _GEN_19530; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19532 = 7'h2b == index ? record_addr_43 : _GEN_19531; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19533 = 7'h2c == index ? record_addr_44 : _GEN_19532; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19534 = 7'h2d == index ? record_addr_45 : _GEN_19533; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19535 = 7'h2e == index ? record_addr_46 : _GEN_19534; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19536 = 7'h2f == index ? record_addr_47 : _GEN_19535; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19537 = 7'h30 == index ? record_addr_48 : _GEN_19536; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19538 = 7'h31 == index ? record_addr_49 : _GEN_19537; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19539 = 7'h32 == index ? record_addr_50 : _GEN_19538; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19540 = 7'h33 == index ? record_addr_51 : _GEN_19539; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19541 = 7'h34 == index ? record_addr_52 : _GEN_19540; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19542 = 7'h35 == index ? record_addr_53 : _GEN_19541; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19543 = 7'h36 == index ? record_addr_54 : _GEN_19542; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19544 = 7'h37 == index ? record_addr_55 : _GEN_19543; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19545 = 7'h38 == index ? record_addr_56 : _GEN_19544; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19546 = 7'h39 == index ? record_addr_57 : _GEN_19545; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19547 = 7'h3a == index ? record_addr_58 : _GEN_19546; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19548 = 7'h3b == index ? record_addr_59 : _GEN_19547; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19549 = 7'h3c == index ? record_addr_60 : _GEN_19548; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19550 = 7'h3d == index ? record_addr_61 : _GEN_19549; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19551 = 7'h3e == index ? record_addr_62 : _GEN_19550; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19552 = 7'h3f == index ? record_addr_63 : _GEN_19551; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19553 = 7'h40 == index ? record_addr_64 : _GEN_19552; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19554 = 7'h41 == index ? record_addr_65 : _GEN_19553; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19555 = 7'h42 == index ? record_addr_66 : _GEN_19554; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19556 = 7'h43 == index ? record_addr_67 : _GEN_19555; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19557 = 7'h44 == index ? record_addr_68 : _GEN_19556; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19558 = 7'h45 == index ? record_addr_69 : _GEN_19557; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19559 = 7'h46 == index ? record_addr_70 : _GEN_19558; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19560 = 7'h47 == index ? record_addr_71 : _GEN_19559; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19561 = 7'h48 == index ? record_addr_72 : _GEN_19560; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19562 = 7'h49 == index ? record_addr_73 : _GEN_19561; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19563 = 7'h4a == index ? record_addr_74 : _GEN_19562; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19564 = 7'h4b == index ? record_addr_75 : _GEN_19563; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19565 = 7'h4c == index ? record_addr_76 : _GEN_19564; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19566 = 7'h4d == index ? record_addr_77 : _GEN_19565; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19567 = 7'h4e == index ? record_addr_78 : _GEN_19566; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19568 = 7'h4f == index ? record_addr_79 : _GEN_19567; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19569 = 7'h50 == index ? record_addr_80 : _GEN_19568; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19570 = 7'h51 == index ? record_addr_81 : _GEN_19569; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19571 = 7'h52 == index ? record_addr_82 : _GEN_19570; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19572 = 7'h53 == index ? record_addr_83 : _GEN_19571; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19573 = 7'h54 == index ? record_addr_84 : _GEN_19572; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19574 = 7'h55 == index ? record_addr_85 : _GEN_19573; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19575 = 7'h56 == index ? record_addr_86 : _GEN_19574; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19576 = 7'h57 == index ? record_addr_87 : _GEN_19575; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19577 = 7'h58 == index ? record_addr_88 : _GEN_19576; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19578 = 7'h59 == index ? record_addr_89 : _GEN_19577; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19579 = 7'h5a == index ? record_addr_90 : _GEN_19578; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19580 = 7'h5b == index ? record_addr_91 : _GEN_19579; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19581 = 7'h5c == index ? record_addr_92 : _GEN_19580; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19582 = 7'h5d == index ? record_addr_93 : _GEN_19581; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19583 = 7'h5e == index ? record_addr_94 : _GEN_19582; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19584 = 7'h5f == index ? record_addr_95 : _GEN_19583; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19585 = 7'h60 == index ? record_addr_96 : _GEN_19584; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19586 = 7'h61 == index ? record_addr_97 : _GEN_19585; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19587 = 7'h62 == index ? record_addr_98 : _GEN_19586; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19588 = 7'h63 == index ? record_addr_99 : _GEN_19587; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19589 = 7'h64 == index ? record_addr_100 : _GEN_19588; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19590 = 7'h65 == index ? record_addr_101 : _GEN_19589; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19591 = 7'h66 == index ? record_addr_102 : _GEN_19590; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19592 = 7'h67 == index ? record_addr_103 : _GEN_19591; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19593 = 7'h68 == index ? record_addr_104 : _GEN_19592; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19594 = 7'h69 == index ? record_addr_105 : _GEN_19593; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19595 = 7'h6a == index ? record_addr_106 : _GEN_19594; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19596 = 7'h6b == index ? record_addr_107 : _GEN_19595; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19597 = 7'h6c == index ? record_addr_108 : _GEN_19596; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19598 = 7'h6d == index ? record_addr_109 : _GEN_19597; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19599 = 7'h6e == index ? record_addr_110 : _GEN_19598; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19600 = 7'h6f == index ? record_addr_111 : _GEN_19599; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19601 = 7'h70 == index ? record_addr_112 : _GEN_19600; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19602 = 7'h71 == index ? record_addr_113 : _GEN_19601; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19603 = 7'h72 == index ? record_addr_114 : _GEN_19602; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19604 = 7'h73 == index ? record_addr_115 : _GEN_19603; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19605 = 7'h74 == index ? record_addr_116 : _GEN_19604; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19606 = 7'h75 == index ? record_addr_117 : _GEN_19605; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19607 = 7'h76 == index ? record_addr_118 : _GEN_19606; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19608 = 7'h77 == index ? record_addr_119 : _GEN_19607; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19609 = 7'h78 == index ? record_addr_120 : _GEN_19608; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19610 = 7'h79 == index ? record_addr_121 : _GEN_19609; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19611 = 7'h7a == index ? record_addr_122 : _GEN_19610; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19612 = 7'h7b == index ? record_addr_123 : _GEN_19611; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19613 = 7'h7c == index ? record_addr_124 : _GEN_19612; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19614 = 7'h7d == index ? record_addr_125 : _GEN_19613; // @[d_cache.scala 374:{11,11}]
  wire [31:0] _GEN_19615 = 7'h7e == index ? record_addr_126 : _GEN_19614; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19618 = 7'h1 == index ? record_olddata_1 : record_olddata_0; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19619 = 7'h2 == index ? record_olddata_2 : _GEN_19618; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19620 = 7'h3 == index ? record_olddata_3 : _GEN_19619; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19621 = 7'h4 == index ? record_olddata_4 : _GEN_19620; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19622 = 7'h5 == index ? record_olddata_5 : _GEN_19621; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19623 = 7'h6 == index ? record_olddata_6 : _GEN_19622; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19624 = 7'h7 == index ? record_olddata_7 : _GEN_19623; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19625 = 7'h8 == index ? record_olddata_8 : _GEN_19624; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19626 = 7'h9 == index ? record_olddata_9 : _GEN_19625; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19627 = 7'ha == index ? record_olddata_10 : _GEN_19626; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19628 = 7'hb == index ? record_olddata_11 : _GEN_19627; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19629 = 7'hc == index ? record_olddata_12 : _GEN_19628; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19630 = 7'hd == index ? record_olddata_13 : _GEN_19629; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19631 = 7'he == index ? record_olddata_14 : _GEN_19630; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19632 = 7'hf == index ? record_olddata_15 : _GEN_19631; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19633 = 7'h10 == index ? record_olddata_16 : _GEN_19632; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19634 = 7'h11 == index ? record_olddata_17 : _GEN_19633; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19635 = 7'h12 == index ? record_olddata_18 : _GEN_19634; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19636 = 7'h13 == index ? record_olddata_19 : _GEN_19635; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19637 = 7'h14 == index ? record_olddata_20 : _GEN_19636; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19638 = 7'h15 == index ? record_olddata_21 : _GEN_19637; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19639 = 7'h16 == index ? record_olddata_22 : _GEN_19638; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19640 = 7'h17 == index ? record_olddata_23 : _GEN_19639; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19641 = 7'h18 == index ? record_olddata_24 : _GEN_19640; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19642 = 7'h19 == index ? record_olddata_25 : _GEN_19641; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19643 = 7'h1a == index ? record_olddata_26 : _GEN_19642; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19644 = 7'h1b == index ? record_olddata_27 : _GEN_19643; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19645 = 7'h1c == index ? record_olddata_28 : _GEN_19644; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19646 = 7'h1d == index ? record_olddata_29 : _GEN_19645; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19647 = 7'h1e == index ? record_olddata_30 : _GEN_19646; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19648 = 7'h1f == index ? record_olddata_31 : _GEN_19647; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19649 = 7'h20 == index ? record_olddata_32 : _GEN_19648; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19650 = 7'h21 == index ? record_olddata_33 : _GEN_19649; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19651 = 7'h22 == index ? record_olddata_34 : _GEN_19650; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19652 = 7'h23 == index ? record_olddata_35 : _GEN_19651; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19653 = 7'h24 == index ? record_olddata_36 : _GEN_19652; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19654 = 7'h25 == index ? record_olddata_37 : _GEN_19653; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19655 = 7'h26 == index ? record_olddata_38 : _GEN_19654; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19656 = 7'h27 == index ? record_olddata_39 : _GEN_19655; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19657 = 7'h28 == index ? record_olddata_40 : _GEN_19656; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19658 = 7'h29 == index ? record_olddata_41 : _GEN_19657; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19659 = 7'h2a == index ? record_olddata_42 : _GEN_19658; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19660 = 7'h2b == index ? record_olddata_43 : _GEN_19659; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19661 = 7'h2c == index ? record_olddata_44 : _GEN_19660; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19662 = 7'h2d == index ? record_olddata_45 : _GEN_19661; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19663 = 7'h2e == index ? record_olddata_46 : _GEN_19662; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19664 = 7'h2f == index ? record_olddata_47 : _GEN_19663; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19665 = 7'h30 == index ? record_olddata_48 : _GEN_19664; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19666 = 7'h31 == index ? record_olddata_49 : _GEN_19665; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19667 = 7'h32 == index ? record_olddata_50 : _GEN_19666; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19668 = 7'h33 == index ? record_olddata_51 : _GEN_19667; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19669 = 7'h34 == index ? record_olddata_52 : _GEN_19668; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19670 = 7'h35 == index ? record_olddata_53 : _GEN_19669; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19671 = 7'h36 == index ? record_olddata_54 : _GEN_19670; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19672 = 7'h37 == index ? record_olddata_55 : _GEN_19671; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19673 = 7'h38 == index ? record_olddata_56 : _GEN_19672; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19674 = 7'h39 == index ? record_olddata_57 : _GEN_19673; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19675 = 7'h3a == index ? record_olddata_58 : _GEN_19674; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19676 = 7'h3b == index ? record_olddata_59 : _GEN_19675; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19677 = 7'h3c == index ? record_olddata_60 : _GEN_19676; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19678 = 7'h3d == index ? record_olddata_61 : _GEN_19677; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19679 = 7'h3e == index ? record_olddata_62 : _GEN_19678; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19680 = 7'h3f == index ? record_olddata_63 : _GEN_19679; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19681 = 7'h40 == index ? record_olddata_64 : _GEN_19680; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19682 = 7'h41 == index ? record_olddata_65 : _GEN_19681; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19683 = 7'h42 == index ? record_olddata_66 : _GEN_19682; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19684 = 7'h43 == index ? record_olddata_67 : _GEN_19683; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19685 = 7'h44 == index ? record_olddata_68 : _GEN_19684; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19686 = 7'h45 == index ? record_olddata_69 : _GEN_19685; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19687 = 7'h46 == index ? record_olddata_70 : _GEN_19686; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19688 = 7'h47 == index ? record_olddata_71 : _GEN_19687; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19689 = 7'h48 == index ? record_olddata_72 : _GEN_19688; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19690 = 7'h49 == index ? record_olddata_73 : _GEN_19689; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19691 = 7'h4a == index ? record_olddata_74 : _GEN_19690; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19692 = 7'h4b == index ? record_olddata_75 : _GEN_19691; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19693 = 7'h4c == index ? record_olddata_76 : _GEN_19692; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19694 = 7'h4d == index ? record_olddata_77 : _GEN_19693; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19695 = 7'h4e == index ? record_olddata_78 : _GEN_19694; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19696 = 7'h4f == index ? record_olddata_79 : _GEN_19695; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19697 = 7'h50 == index ? record_olddata_80 : _GEN_19696; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19698 = 7'h51 == index ? record_olddata_81 : _GEN_19697; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19699 = 7'h52 == index ? record_olddata_82 : _GEN_19698; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19700 = 7'h53 == index ? record_olddata_83 : _GEN_19699; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19701 = 7'h54 == index ? record_olddata_84 : _GEN_19700; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19702 = 7'h55 == index ? record_olddata_85 : _GEN_19701; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19703 = 7'h56 == index ? record_olddata_86 : _GEN_19702; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19704 = 7'h57 == index ? record_olddata_87 : _GEN_19703; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19705 = 7'h58 == index ? record_olddata_88 : _GEN_19704; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19706 = 7'h59 == index ? record_olddata_89 : _GEN_19705; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19707 = 7'h5a == index ? record_olddata_90 : _GEN_19706; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19708 = 7'h5b == index ? record_olddata_91 : _GEN_19707; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19709 = 7'h5c == index ? record_olddata_92 : _GEN_19708; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19710 = 7'h5d == index ? record_olddata_93 : _GEN_19709; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19711 = 7'h5e == index ? record_olddata_94 : _GEN_19710; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19712 = 7'h5f == index ? record_olddata_95 : _GEN_19711; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19713 = 7'h60 == index ? record_olddata_96 : _GEN_19712; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19714 = 7'h61 == index ? record_olddata_97 : _GEN_19713; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19715 = 7'h62 == index ? record_olddata_98 : _GEN_19714; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19716 = 7'h63 == index ? record_olddata_99 : _GEN_19715; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19717 = 7'h64 == index ? record_olddata_100 : _GEN_19716; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19718 = 7'h65 == index ? record_olddata_101 : _GEN_19717; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19719 = 7'h66 == index ? record_olddata_102 : _GEN_19718; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19720 = 7'h67 == index ? record_olddata_103 : _GEN_19719; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19721 = 7'h68 == index ? record_olddata_104 : _GEN_19720; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19722 = 7'h69 == index ? record_olddata_105 : _GEN_19721; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19723 = 7'h6a == index ? record_olddata_106 : _GEN_19722; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19724 = 7'h6b == index ? record_olddata_107 : _GEN_19723; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19725 = 7'h6c == index ? record_olddata_108 : _GEN_19724; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19726 = 7'h6d == index ? record_olddata_109 : _GEN_19725; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19727 = 7'h6e == index ? record_olddata_110 : _GEN_19726; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19728 = 7'h6f == index ? record_olddata_111 : _GEN_19727; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19729 = 7'h70 == index ? record_olddata_112 : _GEN_19728; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19730 = 7'h71 == index ? record_olddata_113 : _GEN_19729; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19731 = 7'h72 == index ? record_olddata_114 : _GEN_19730; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19732 = 7'h73 == index ? record_olddata_115 : _GEN_19731; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19733 = 7'h74 == index ? record_olddata_116 : _GEN_19732; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19734 = 7'h75 == index ? record_olddata_117 : _GEN_19733; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19735 = 7'h76 == index ? record_olddata_118 : _GEN_19734; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19736 = 7'h77 == index ? record_olddata_119 : _GEN_19735; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19737 = 7'h78 == index ? record_olddata_120 : _GEN_19736; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19738 = 7'h79 == index ? record_olddata_121 : _GEN_19737; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19739 = 7'h7a == index ? record_olddata_122 : _GEN_19738; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19740 = 7'h7b == index ? record_olddata_123 : _GEN_19739; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19741 = 7'h7c == index ? record_olddata_124 : _GEN_19740; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19742 = 7'h7d == index ? record_olddata_125 : _GEN_19741; // @[d_cache.scala 374:{11,11}]
  wire [63:0] _GEN_19743 = 7'h7e == index ? record_olddata_126 : _GEN_19742; // @[d_cache.scala 374:{11,11}]
  wire [41:0] _GEN_20774 = reset ? 42'h0 : _GEN_19008; // @[d_cache.scala 38:{34,34}]
  wire  _GEN_20776 = ~_T_14 & _T_15; // @[d_cache.scala 99:27]
  assign io_to_lsu_arready = state == 3'h0 ? io_from_axi_arready : _GEN_19085; // @[d_cache.scala 210:23 212:27]
  assign io_to_lsu_rdata = state == 3'h0 ? 64'h0 : _GEN_19084; // @[d_cache.scala 210:23 211:25]
  assign io_to_lsu_rvalid = state == 3'h0 ? 1'h0 : _GEN_19086; // @[d_cache.scala 210:23 213:26]
  assign io_to_lsu_awready = state == 3'h0 ? io_from_axi_awready : _GEN_19088; // @[d_cache.scala 210:23 216:27]
  assign io_to_lsu_wready = state == 3'h0 ? 1'h0 : _GEN_19087; // @[d_cache.scala 210:23 214:26]
  assign io_to_lsu_bvalid = state == 3'h0 ? 1'h0 : _GEN_19089; // @[d_cache.scala 210:23 215:26]
  assign io_to_axi_araddr = _GEN_19097[31:0];
  assign io_to_axi_arvalid = state == 3'h0 ? 1'h0 : _GEN_19075; // @[d_cache.scala 210:23 217:27]
  assign io_to_axi_rready = state == 3'h0 ? io_from_lsu_rready : _GEN_19077; // @[d_cache.scala 210:23 219:26]
  assign io_to_axi_awaddr = state == 3'h0 ? 32'h0 : _GEN_19078; // @[d_cache.scala 210:23 220:26]
  assign io_to_axi_awvalid = state == 3'h0 ? 1'h0 : _GEN_19079; // @[d_cache.scala 210:23 221:27]
  assign io_to_axi_wdata = state == 3'h0 ? 64'h0 : _GEN_19080; // @[d_cache.scala 210:23 222:25]
  assign io_to_axi_wstrb = state == 3'h0 ? 8'h0 : _GEN_19081; // @[d_cache.scala 210:23 223:25]
  assign io_to_axi_wvalid = state == 3'h0 ? 1'h0 : _GEN_19082; // @[d_cache.scala 210:23 224:26]
  assign io_to_axi_bready = state == 3'h0 ? io_from_lsu_bready : _GEN_19083; // @[d_cache.scala 210:23 225:26]
  always @(posedge clock) begin
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_0 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_0 <= _GEN_3083;
        end else begin
          ram_0_0 <= _GEN_12975;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_1 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_1 <= _GEN_3084;
        end else begin
          ram_0_1 <= _GEN_12976;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_2 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_2 <= _GEN_3085;
        end else begin
          ram_0_2 <= _GEN_12977;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_3 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_3 <= _GEN_3086;
        end else begin
          ram_0_3 <= _GEN_12978;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_4 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_4 <= _GEN_3087;
        end else begin
          ram_0_4 <= _GEN_12979;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_5 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_5 <= _GEN_3088;
        end else begin
          ram_0_5 <= _GEN_12980;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_6 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_6 <= _GEN_3089;
        end else begin
          ram_0_6 <= _GEN_12981;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_7 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_7 <= _GEN_3090;
        end else begin
          ram_0_7 <= _GEN_12982;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_8 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_8 <= _GEN_3091;
        end else begin
          ram_0_8 <= _GEN_12983;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_9 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_9 <= _GEN_3092;
        end else begin
          ram_0_9 <= _GEN_12984;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_10 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_10 <= _GEN_3093;
        end else begin
          ram_0_10 <= _GEN_12985;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_11 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_11 <= _GEN_3094;
        end else begin
          ram_0_11 <= _GEN_12986;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_12 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_12 <= _GEN_3095;
        end else begin
          ram_0_12 <= _GEN_12987;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_13 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_13 <= _GEN_3096;
        end else begin
          ram_0_13 <= _GEN_12988;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_14 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_14 <= _GEN_3097;
        end else begin
          ram_0_14 <= _GEN_12989;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_15 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_15 <= _GEN_3098;
        end else begin
          ram_0_15 <= _GEN_12990;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_16 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_16 <= _GEN_3099;
        end else begin
          ram_0_16 <= _GEN_12991;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_17 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_17 <= _GEN_3100;
        end else begin
          ram_0_17 <= _GEN_12992;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_18 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_18 <= _GEN_3101;
        end else begin
          ram_0_18 <= _GEN_12993;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_19 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_19 <= _GEN_3102;
        end else begin
          ram_0_19 <= _GEN_12994;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_20 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_20 <= _GEN_3103;
        end else begin
          ram_0_20 <= _GEN_12995;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_21 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_21 <= _GEN_3104;
        end else begin
          ram_0_21 <= _GEN_12996;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_22 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_22 <= _GEN_3105;
        end else begin
          ram_0_22 <= _GEN_12997;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_23 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_23 <= _GEN_3106;
        end else begin
          ram_0_23 <= _GEN_12998;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_24 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_24 <= _GEN_3107;
        end else begin
          ram_0_24 <= _GEN_12999;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_25 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_25 <= _GEN_3108;
        end else begin
          ram_0_25 <= _GEN_13000;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_26 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_26 <= _GEN_3109;
        end else begin
          ram_0_26 <= _GEN_13001;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_27 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_27 <= _GEN_3110;
        end else begin
          ram_0_27 <= _GEN_13002;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_28 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_28 <= _GEN_3111;
        end else begin
          ram_0_28 <= _GEN_13003;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_29 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_29 <= _GEN_3112;
        end else begin
          ram_0_29 <= _GEN_13004;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_30 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_30 <= _GEN_3113;
        end else begin
          ram_0_30 <= _GEN_13005;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_31 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_31 <= _GEN_3114;
        end else begin
          ram_0_31 <= _GEN_13006;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_32 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_32 <= _GEN_3115;
        end else begin
          ram_0_32 <= _GEN_13007;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_33 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_33 <= _GEN_3116;
        end else begin
          ram_0_33 <= _GEN_13008;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_34 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_34 <= _GEN_3117;
        end else begin
          ram_0_34 <= _GEN_13009;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_35 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_35 <= _GEN_3118;
        end else begin
          ram_0_35 <= _GEN_13010;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_36 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_36 <= _GEN_3119;
        end else begin
          ram_0_36 <= _GEN_13011;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_37 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_37 <= _GEN_3120;
        end else begin
          ram_0_37 <= _GEN_13012;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_38 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_38 <= _GEN_3121;
        end else begin
          ram_0_38 <= _GEN_13013;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_39 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_39 <= _GEN_3122;
        end else begin
          ram_0_39 <= _GEN_13014;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_40 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_40 <= _GEN_3123;
        end else begin
          ram_0_40 <= _GEN_13015;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_41 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_41 <= _GEN_3124;
        end else begin
          ram_0_41 <= _GEN_13016;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_42 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_42 <= _GEN_3125;
        end else begin
          ram_0_42 <= _GEN_13017;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_43 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_43 <= _GEN_3126;
        end else begin
          ram_0_43 <= _GEN_13018;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_44 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_44 <= _GEN_3127;
        end else begin
          ram_0_44 <= _GEN_13019;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_45 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_45 <= _GEN_3128;
        end else begin
          ram_0_45 <= _GEN_13020;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_46 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_46 <= _GEN_3129;
        end else begin
          ram_0_46 <= _GEN_13021;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_47 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_47 <= _GEN_3130;
        end else begin
          ram_0_47 <= _GEN_13022;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_48 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_48 <= _GEN_3131;
        end else begin
          ram_0_48 <= _GEN_13023;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_49 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_49 <= _GEN_3132;
        end else begin
          ram_0_49 <= _GEN_13024;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_50 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_50 <= _GEN_3133;
        end else begin
          ram_0_50 <= _GEN_13025;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_51 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_51 <= _GEN_3134;
        end else begin
          ram_0_51 <= _GEN_13026;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_52 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_52 <= _GEN_3135;
        end else begin
          ram_0_52 <= _GEN_13027;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_53 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_53 <= _GEN_3136;
        end else begin
          ram_0_53 <= _GEN_13028;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_54 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_54 <= _GEN_3137;
        end else begin
          ram_0_54 <= _GEN_13029;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_55 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_55 <= _GEN_3138;
        end else begin
          ram_0_55 <= _GEN_13030;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_56 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_56 <= _GEN_3139;
        end else begin
          ram_0_56 <= _GEN_13031;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_57 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_57 <= _GEN_3140;
        end else begin
          ram_0_57 <= _GEN_13032;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_58 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_58 <= _GEN_3141;
        end else begin
          ram_0_58 <= _GEN_13033;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_59 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_59 <= _GEN_3142;
        end else begin
          ram_0_59 <= _GEN_13034;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_60 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_60 <= _GEN_3143;
        end else begin
          ram_0_60 <= _GEN_13035;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_61 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_61 <= _GEN_3144;
        end else begin
          ram_0_61 <= _GEN_13036;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_62 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_62 <= _GEN_3145;
        end else begin
          ram_0_62 <= _GEN_13037;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_63 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_63 <= _GEN_3146;
        end else begin
          ram_0_63 <= _GEN_13038;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_64 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_64 <= _GEN_3147;
        end else begin
          ram_0_64 <= _GEN_13039;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_65 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_65 <= _GEN_3148;
        end else begin
          ram_0_65 <= _GEN_13040;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_66 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_66 <= _GEN_3149;
        end else begin
          ram_0_66 <= _GEN_13041;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_67 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_67 <= _GEN_3150;
        end else begin
          ram_0_67 <= _GEN_13042;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_68 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_68 <= _GEN_3151;
        end else begin
          ram_0_68 <= _GEN_13043;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_69 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_69 <= _GEN_3152;
        end else begin
          ram_0_69 <= _GEN_13044;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_70 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_70 <= _GEN_3153;
        end else begin
          ram_0_70 <= _GEN_13045;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_71 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_71 <= _GEN_3154;
        end else begin
          ram_0_71 <= _GEN_13046;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_72 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_72 <= _GEN_3155;
        end else begin
          ram_0_72 <= _GEN_13047;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_73 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_73 <= _GEN_3156;
        end else begin
          ram_0_73 <= _GEN_13048;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_74 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_74 <= _GEN_3157;
        end else begin
          ram_0_74 <= _GEN_13049;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_75 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_75 <= _GEN_3158;
        end else begin
          ram_0_75 <= _GEN_13050;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_76 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_76 <= _GEN_3159;
        end else begin
          ram_0_76 <= _GEN_13051;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_77 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_77 <= _GEN_3160;
        end else begin
          ram_0_77 <= _GEN_13052;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_78 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_78 <= _GEN_3161;
        end else begin
          ram_0_78 <= _GEN_13053;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_79 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_79 <= _GEN_3162;
        end else begin
          ram_0_79 <= _GEN_13054;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_80 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_80 <= _GEN_3163;
        end else begin
          ram_0_80 <= _GEN_13055;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_81 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_81 <= _GEN_3164;
        end else begin
          ram_0_81 <= _GEN_13056;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_82 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_82 <= _GEN_3165;
        end else begin
          ram_0_82 <= _GEN_13057;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_83 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_83 <= _GEN_3166;
        end else begin
          ram_0_83 <= _GEN_13058;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_84 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_84 <= _GEN_3167;
        end else begin
          ram_0_84 <= _GEN_13059;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_85 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_85 <= _GEN_3168;
        end else begin
          ram_0_85 <= _GEN_13060;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_86 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_86 <= _GEN_3169;
        end else begin
          ram_0_86 <= _GEN_13061;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_87 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_87 <= _GEN_3170;
        end else begin
          ram_0_87 <= _GEN_13062;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_88 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_88 <= _GEN_3171;
        end else begin
          ram_0_88 <= _GEN_13063;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_89 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_89 <= _GEN_3172;
        end else begin
          ram_0_89 <= _GEN_13064;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_90 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_90 <= _GEN_3173;
        end else begin
          ram_0_90 <= _GEN_13065;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_91 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_91 <= _GEN_3174;
        end else begin
          ram_0_91 <= _GEN_13066;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_92 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_92 <= _GEN_3175;
        end else begin
          ram_0_92 <= _GEN_13067;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_93 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_93 <= _GEN_3176;
        end else begin
          ram_0_93 <= _GEN_13068;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_94 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_94 <= _GEN_3177;
        end else begin
          ram_0_94 <= _GEN_13069;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_95 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_95 <= _GEN_3178;
        end else begin
          ram_0_95 <= _GEN_13070;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_96 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_96 <= _GEN_3179;
        end else begin
          ram_0_96 <= _GEN_13071;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_97 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_97 <= _GEN_3180;
        end else begin
          ram_0_97 <= _GEN_13072;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_98 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_98 <= _GEN_3181;
        end else begin
          ram_0_98 <= _GEN_13073;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_99 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_99 <= _GEN_3182;
        end else begin
          ram_0_99 <= _GEN_13074;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_100 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_100 <= _GEN_3183;
        end else begin
          ram_0_100 <= _GEN_13075;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_101 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_101 <= _GEN_3184;
        end else begin
          ram_0_101 <= _GEN_13076;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_102 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_102 <= _GEN_3185;
        end else begin
          ram_0_102 <= _GEN_13077;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_103 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_103 <= _GEN_3186;
        end else begin
          ram_0_103 <= _GEN_13078;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_104 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_104 <= _GEN_3187;
        end else begin
          ram_0_104 <= _GEN_13079;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_105 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_105 <= _GEN_3188;
        end else begin
          ram_0_105 <= _GEN_13080;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_106 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_106 <= _GEN_3189;
        end else begin
          ram_0_106 <= _GEN_13081;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_107 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_107 <= _GEN_3190;
        end else begin
          ram_0_107 <= _GEN_13082;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_108 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_108 <= _GEN_3191;
        end else begin
          ram_0_108 <= _GEN_13083;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_109 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_109 <= _GEN_3192;
        end else begin
          ram_0_109 <= _GEN_13084;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_110 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_110 <= _GEN_3193;
        end else begin
          ram_0_110 <= _GEN_13085;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_111 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_111 <= _GEN_3194;
        end else begin
          ram_0_111 <= _GEN_13086;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_112 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_112 <= _GEN_3195;
        end else begin
          ram_0_112 <= _GEN_13087;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_113 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_113 <= _GEN_3196;
        end else begin
          ram_0_113 <= _GEN_13088;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_114 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_114 <= _GEN_3197;
        end else begin
          ram_0_114 <= _GEN_13089;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_115 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_115 <= _GEN_3198;
        end else begin
          ram_0_115 <= _GEN_13090;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_116 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_116 <= _GEN_3199;
        end else begin
          ram_0_116 <= _GEN_13091;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_117 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_117 <= _GEN_3200;
        end else begin
          ram_0_117 <= _GEN_13092;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_118 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_118 <= _GEN_3201;
        end else begin
          ram_0_118 <= _GEN_13093;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_119 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_119 <= _GEN_3202;
        end else begin
          ram_0_119 <= _GEN_13094;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_120 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_120 <= _GEN_3203;
        end else begin
          ram_0_120 <= _GEN_13095;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_121 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_121 <= _GEN_3204;
        end else begin
          ram_0_121 <= _GEN_13096;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_122 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_122 <= _GEN_3205;
        end else begin
          ram_0_122 <= _GEN_13097;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_123 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_123 <= _GEN_3206;
        end else begin
          ram_0_123 <= _GEN_13098;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_124 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_124 <= _GEN_3207;
        end else begin
          ram_0_124 <= _GEN_13099;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_125 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_125 <= _GEN_3208;
        end else begin
          ram_0_125 <= _GEN_13100;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_126 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_126 <= _GEN_3209;
        end else begin
          ram_0_126 <= _GEN_13101;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_127 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_127 <= _GEN_3210;
        end else begin
          ram_0_127 <= _GEN_13102;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_0 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_0 <= _GEN_3467;
        end else begin
          ram_1_0 <= _GEN_13360;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_1 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_1 <= _GEN_3468;
        end else begin
          ram_1_1 <= _GEN_13361;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_2 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_2 <= _GEN_3469;
        end else begin
          ram_1_2 <= _GEN_13362;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_3 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_3 <= _GEN_3470;
        end else begin
          ram_1_3 <= _GEN_13363;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_4 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_4 <= _GEN_3471;
        end else begin
          ram_1_4 <= _GEN_13364;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_5 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_5 <= _GEN_3472;
        end else begin
          ram_1_5 <= _GEN_13365;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_6 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_6 <= _GEN_3473;
        end else begin
          ram_1_6 <= _GEN_13366;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_7 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_7 <= _GEN_3474;
        end else begin
          ram_1_7 <= _GEN_13367;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_8 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_8 <= _GEN_3475;
        end else begin
          ram_1_8 <= _GEN_13368;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_9 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_9 <= _GEN_3476;
        end else begin
          ram_1_9 <= _GEN_13369;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_10 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_10 <= _GEN_3477;
        end else begin
          ram_1_10 <= _GEN_13370;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_11 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_11 <= _GEN_3478;
        end else begin
          ram_1_11 <= _GEN_13371;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_12 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_12 <= _GEN_3479;
        end else begin
          ram_1_12 <= _GEN_13372;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_13 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_13 <= _GEN_3480;
        end else begin
          ram_1_13 <= _GEN_13373;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_14 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_14 <= _GEN_3481;
        end else begin
          ram_1_14 <= _GEN_13374;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_15 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_15 <= _GEN_3482;
        end else begin
          ram_1_15 <= _GEN_13375;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_16 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_16 <= _GEN_3483;
        end else begin
          ram_1_16 <= _GEN_13376;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_17 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_17 <= _GEN_3484;
        end else begin
          ram_1_17 <= _GEN_13377;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_18 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_18 <= _GEN_3485;
        end else begin
          ram_1_18 <= _GEN_13378;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_19 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_19 <= _GEN_3486;
        end else begin
          ram_1_19 <= _GEN_13379;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_20 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_20 <= _GEN_3487;
        end else begin
          ram_1_20 <= _GEN_13380;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_21 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_21 <= _GEN_3488;
        end else begin
          ram_1_21 <= _GEN_13381;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_22 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_22 <= _GEN_3489;
        end else begin
          ram_1_22 <= _GEN_13382;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_23 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_23 <= _GEN_3490;
        end else begin
          ram_1_23 <= _GEN_13383;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_24 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_24 <= _GEN_3491;
        end else begin
          ram_1_24 <= _GEN_13384;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_25 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_25 <= _GEN_3492;
        end else begin
          ram_1_25 <= _GEN_13385;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_26 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_26 <= _GEN_3493;
        end else begin
          ram_1_26 <= _GEN_13386;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_27 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_27 <= _GEN_3494;
        end else begin
          ram_1_27 <= _GEN_13387;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_28 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_28 <= _GEN_3495;
        end else begin
          ram_1_28 <= _GEN_13388;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_29 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_29 <= _GEN_3496;
        end else begin
          ram_1_29 <= _GEN_13389;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_30 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_30 <= _GEN_3497;
        end else begin
          ram_1_30 <= _GEN_13390;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_31 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_31 <= _GEN_3498;
        end else begin
          ram_1_31 <= _GEN_13391;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_32 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_32 <= _GEN_3499;
        end else begin
          ram_1_32 <= _GEN_13392;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_33 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_33 <= _GEN_3500;
        end else begin
          ram_1_33 <= _GEN_13393;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_34 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_34 <= _GEN_3501;
        end else begin
          ram_1_34 <= _GEN_13394;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_35 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_35 <= _GEN_3502;
        end else begin
          ram_1_35 <= _GEN_13395;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_36 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_36 <= _GEN_3503;
        end else begin
          ram_1_36 <= _GEN_13396;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_37 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_37 <= _GEN_3504;
        end else begin
          ram_1_37 <= _GEN_13397;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_38 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_38 <= _GEN_3505;
        end else begin
          ram_1_38 <= _GEN_13398;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_39 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_39 <= _GEN_3506;
        end else begin
          ram_1_39 <= _GEN_13399;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_40 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_40 <= _GEN_3507;
        end else begin
          ram_1_40 <= _GEN_13400;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_41 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_41 <= _GEN_3508;
        end else begin
          ram_1_41 <= _GEN_13401;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_42 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_42 <= _GEN_3509;
        end else begin
          ram_1_42 <= _GEN_13402;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_43 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_43 <= _GEN_3510;
        end else begin
          ram_1_43 <= _GEN_13403;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_44 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_44 <= _GEN_3511;
        end else begin
          ram_1_44 <= _GEN_13404;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_45 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_45 <= _GEN_3512;
        end else begin
          ram_1_45 <= _GEN_13405;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_46 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_46 <= _GEN_3513;
        end else begin
          ram_1_46 <= _GEN_13406;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_47 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_47 <= _GEN_3514;
        end else begin
          ram_1_47 <= _GEN_13407;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_48 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_48 <= _GEN_3515;
        end else begin
          ram_1_48 <= _GEN_13408;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_49 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_49 <= _GEN_3516;
        end else begin
          ram_1_49 <= _GEN_13409;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_50 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_50 <= _GEN_3517;
        end else begin
          ram_1_50 <= _GEN_13410;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_51 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_51 <= _GEN_3518;
        end else begin
          ram_1_51 <= _GEN_13411;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_52 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_52 <= _GEN_3519;
        end else begin
          ram_1_52 <= _GEN_13412;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_53 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_53 <= _GEN_3520;
        end else begin
          ram_1_53 <= _GEN_13413;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_54 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_54 <= _GEN_3521;
        end else begin
          ram_1_54 <= _GEN_13414;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_55 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_55 <= _GEN_3522;
        end else begin
          ram_1_55 <= _GEN_13415;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_56 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_56 <= _GEN_3523;
        end else begin
          ram_1_56 <= _GEN_13416;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_57 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_57 <= _GEN_3524;
        end else begin
          ram_1_57 <= _GEN_13417;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_58 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_58 <= _GEN_3525;
        end else begin
          ram_1_58 <= _GEN_13418;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_59 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_59 <= _GEN_3526;
        end else begin
          ram_1_59 <= _GEN_13419;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_60 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_60 <= _GEN_3527;
        end else begin
          ram_1_60 <= _GEN_13420;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_61 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_61 <= _GEN_3528;
        end else begin
          ram_1_61 <= _GEN_13421;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_62 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_62 <= _GEN_3529;
        end else begin
          ram_1_62 <= _GEN_13422;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_63 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_63 <= _GEN_3530;
        end else begin
          ram_1_63 <= _GEN_13423;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_64 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_64 <= _GEN_3531;
        end else begin
          ram_1_64 <= _GEN_13424;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_65 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_65 <= _GEN_3532;
        end else begin
          ram_1_65 <= _GEN_13425;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_66 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_66 <= _GEN_3533;
        end else begin
          ram_1_66 <= _GEN_13426;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_67 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_67 <= _GEN_3534;
        end else begin
          ram_1_67 <= _GEN_13427;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_68 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_68 <= _GEN_3535;
        end else begin
          ram_1_68 <= _GEN_13428;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_69 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_69 <= _GEN_3536;
        end else begin
          ram_1_69 <= _GEN_13429;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_70 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_70 <= _GEN_3537;
        end else begin
          ram_1_70 <= _GEN_13430;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_71 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_71 <= _GEN_3538;
        end else begin
          ram_1_71 <= _GEN_13431;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_72 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_72 <= _GEN_3539;
        end else begin
          ram_1_72 <= _GEN_13432;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_73 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_73 <= _GEN_3540;
        end else begin
          ram_1_73 <= _GEN_13433;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_74 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_74 <= _GEN_3541;
        end else begin
          ram_1_74 <= _GEN_13434;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_75 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_75 <= _GEN_3542;
        end else begin
          ram_1_75 <= _GEN_13435;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_76 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_76 <= _GEN_3543;
        end else begin
          ram_1_76 <= _GEN_13436;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_77 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_77 <= _GEN_3544;
        end else begin
          ram_1_77 <= _GEN_13437;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_78 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_78 <= _GEN_3545;
        end else begin
          ram_1_78 <= _GEN_13438;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_79 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_79 <= _GEN_3546;
        end else begin
          ram_1_79 <= _GEN_13439;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_80 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_80 <= _GEN_3547;
        end else begin
          ram_1_80 <= _GEN_13440;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_81 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_81 <= _GEN_3548;
        end else begin
          ram_1_81 <= _GEN_13441;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_82 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_82 <= _GEN_3549;
        end else begin
          ram_1_82 <= _GEN_13442;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_83 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_83 <= _GEN_3550;
        end else begin
          ram_1_83 <= _GEN_13443;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_84 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_84 <= _GEN_3551;
        end else begin
          ram_1_84 <= _GEN_13444;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_85 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_85 <= _GEN_3552;
        end else begin
          ram_1_85 <= _GEN_13445;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_86 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_86 <= _GEN_3553;
        end else begin
          ram_1_86 <= _GEN_13446;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_87 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_87 <= _GEN_3554;
        end else begin
          ram_1_87 <= _GEN_13447;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_88 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_88 <= _GEN_3555;
        end else begin
          ram_1_88 <= _GEN_13448;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_89 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_89 <= _GEN_3556;
        end else begin
          ram_1_89 <= _GEN_13449;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_90 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_90 <= _GEN_3557;
        end else begin
          ram_1_90 <= _GEN_13450;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_91 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_91 <= _GEN_3558;
        end else begin
          ram_1_91 <= _GEN_13451;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_92 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_92 <= _GEN_3559;
        end else begin
          ram_1_92 <= _GEN_13452;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_93 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_93 <= _GEN_3560;
        end else begin
          ram_1_93 <= _GEN_13453;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_94 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_94 <= _GEN_3561;
        end else begin
          ram_1_94 <= _GEN_13454;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_95 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_95 <= _GEN_3562;
        end else begin
          ram_1_95 <= _GEN_13455;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_96 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_96 <= _GEN_3563;
        end else begin
          ram_1_96 <= _GEN_13456;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_97 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_97 <= _GEN_3564;
        end else begin
          ram_1_97 <= _GEN_13457;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_98 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_98 <= _GEN_3565;
        end else begin
          ram_1_98 <= _GEN_13458;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_99 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_99 <= _GEN_3566;
        end else begin
          ram_1_99 <= _GEN_13459;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_100 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_100 <= _GEN_3567;
        end else begin
          ram_1_100 <= _GEN_13460;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_101 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_101 <= _GEN_3568;
        end else begin
          ram_1_101 <= _GEN_13461;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_102 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_102 <= _GEN_3569;
        end else begin
          ram_1_102 <= _GEN_13462;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_103 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_103 <= _GEN_3570;
        end else begin
          ram_1_103 <= _GEN_13463;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_104 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_104 <= _GEN_3571;
        end else begin
          ram_1_104 <= _GEN_13464;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_105 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_105 <= _GEN_3572;
        end else begin
          ram_1_105 <= _GEN_13465;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_106 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_106 <= _GEN_3573;
        end else begin
          ram_1_106 <= _GEN_13466;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_107 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_107 <= _GEN_3574;
        end else begin
          ram_1_107 <= _GEN_13467;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_108 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_108 <= _GEN_3575;
        end else begin
          ram_1_108 <= _GEN_13468;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_109 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_109 <= _GEN_3576;
        end else begin
          ram_1_109 <= _GEN_13469;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_110 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_110 <= _GEN_3577;
        end else begin
          ram_1_110 <= _GEN_13470;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_111 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_111 <= _GEN_3578;
        end else begin
          ram_1_111 <= _GEN_13471;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_112 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_112 <= _GEN_3579;
        end else begin
          ram_1_112 <= _GEN_13472;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_113 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_113 <= _GEN_3580;
        end else begin
          ram_1_113 <= _GEN_13473;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_114 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_114 <= _GEN_3581;
        end else begin
          ram_1_114 <= _GEN_13474;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_115 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_115 <= _GEN_3582;
        end else begin
          ram_1_115 <= _GEN_13475;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_116 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_116 <= _GEN_3583;
        end else begin
          ram_1_116 <= _GEN_13476;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_117 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_117 <= _GEN_3584;
        end else begin
          ram_1_117 <= _GEN_13477;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_118 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_118 <= _GEN_3585;
        end else begin
          ram_1_118 <= _GEN_13478;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_119 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_119 <= _GEN_3586;
        end else begin
          ram_1_119 <= _GEN_13479;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_120 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_120 <= _GEN_3587;
        end else begin
          ram_1_120 <= _GEN_13480;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_121 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_121 <= _GEN_3588;
        end else begin
          ram_1_121 <= _GEN_13481;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_122 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_122 <= _GEN_3589;
        end else begin
          ram_1_122 <= _GEN_13482;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_123 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_123 <= _GEN_3590;
        end else begin
          ram_1_123 <= _GEN_13483;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_124 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_124 <= _GEN_3591;
        end else begin
          ram_1_124 <= _GEN_13484;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_125 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_125 <= _GEN_3592;
        end else begin
          ram_1_125 <= _GEN_13485;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_126 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_126 <= _GEN_3593;
        end else begin
          ram_1_126 <= _GEN_13486;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_127 <= 64'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_127 <= _GEN_3594;
        end else begin
          ram_1_127 <= _GEN_13487;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_0 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_0 <= _GEN_3595;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_1 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_1 <= _GEN_3596;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_2 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_2 <= _GEN_3597;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_3 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_3 <= _GEN_3598;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_4 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_4 <= _GEN_3599;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_5 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_5 <= _GEN_3600;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_6 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_6 <= _GEN_3601;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_7 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_7 <= _GEN_3602;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_8 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_8 <= _GEN_3603;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_9 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_9 <= _GEN_3604;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_10 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_10 <= _GEN_3605;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_11 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_11 <= _GEN_3606;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_12 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_12 <= _GEN_3607;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_13 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_13 <= _GEN_3608;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_14 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_14 <= _GEN_3609;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_15 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_15 <= _GEN_3610;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_16 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_16 <= _GEN_3611;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_17 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_17 <= _GEN_3612;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_18 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_18 <= _GEN_3613;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_19 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_19 <= _GEN_3614;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_20 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_20 <= _GEN_3615;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_21 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_21 <= _GEN_3616;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_22 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_22 <= _GEN_3617;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_23 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_23 <= _GEN_3618;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_24 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_24 <= _GEN_3619;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_25 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_25 <= _GEN_3620;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_26 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_26 <= _GEN_3621;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_27 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_27 <= _GEN_3622;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_28 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_28 <= _GEN_3623;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_29 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_29 <= _GEN_3624;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_30 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_30 <= _GEN_3625;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_31 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_31 <= _GEN_3626;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_32 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_32 <= _GEN_3627;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_33 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_33 <= _GEN_3628;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_34 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_34 <= _GEN_3629;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_35 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_35 <= _GEN_3630;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_36 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_36 <= _GEN_3631;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_37 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_37 <= _GEN_3632;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_38 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_38 <= _GEN_3633;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_39 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_39 <= _GEN_3634;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_40 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_40 <= _GEN_3635;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_41 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_41 <= _GEN_3636;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_42 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_42 <= _GEN_3637;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_43 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_43 <= _GEN_3638;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_44 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_44 <= _GEN_3639;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_45 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_45 <= _GEN_3640;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_46 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_46 <= _GEN_3641;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_47 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_47 <= _GEN_3642;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_48 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_48 <= _GEN_3643;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_49 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_49 <= _GEN_3644;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_50 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_50 <= _GEN_3645;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_51 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_51 <= _GEN_3646;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_52 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_52 <= _GEN_3647;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_53 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_53 <= _GEN_3648;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_54 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_54 <= _GEN_3649;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_55 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_55 <= _GEN_3650;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_56 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_56 <= _GEN_3651;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_57 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_57 <= _GEN_3652;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_58 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_58 <= _GEN_3653;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_59 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_59 <= _GEN_3654;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_60 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_60 <= _GEN_3655;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_61 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_61 <= _GEN_3656;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_62 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_62 <= _GEN_3657;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_63 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_63 <= _GEN_3658;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_64 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_64 <= _GEN_3659;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_65 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_65 <= _GEN_3660;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_66 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_66 <= _GEN_3661;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_67 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_67 <= _GEN_3662;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_68 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_68 <= _GEN_3663;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_69 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_69 <= _GEN_3664;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_70 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_70 <= _GEN_3665;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_71 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_71 <= _GEN_3666;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_72 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_72 <= _GEN_3667;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_73 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_73 <= _GEN_3668;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_74 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_74 <= _GEN_3669;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_75 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_75 <= _GEN_3670;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_76 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_76 <= _GEN_3671;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_77 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_77 <= _GEN_3672;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_78 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_78 <= _GEN_3673;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_79 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_79 <= _GEN_3674;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_80 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_80 <= _GEN_3675;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_81 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_81 <= _GEN_3676;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_82 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_82 <= _GEN_3677;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_83 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_83 <= _GEN_3678;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_84 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_84 <= _GEN_3679;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_85 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_85 <= _GEN_3680;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_86 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_86 <= _GEN_3681;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_87 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_87 <= _GEN_3682;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_88 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_88 <= _GEN_3683;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_89 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_89 <= _GEN_3684;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_90 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_90 <= _GEN_3685;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_91 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_91 <= _GEN_3686;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_92 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_92 <= _GEN_3687;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_93 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_93 <= _GEN_3688;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_94 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_94 <= _GEN_3689;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_95 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_95 <= _GEN_3690;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_96 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_96 <= _GEN_3691;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_97 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_97 <= _GEN_3692;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_98 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_98 <= _GEN_3693;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_99 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_99 <= _GEN_3694;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_100 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_100 <= _GEN_3695;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_101 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_101 <= _GEN_3696;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_102 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_102 <= _GEN_3697;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_103 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_103 <= _GEN_3698;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_104 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_104 <= _GEN_3699;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_105 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_105 <= _GEN_3700;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_106 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_106 <= _GEN_3701;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_107 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_107 <= _GEN_3702;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_108 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_108 <= _GEN_3703;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_109 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_109 <= _GEN_3704;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_110 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_110 <= _GEN_3705;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_111 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_111 <= _GEN_3706;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_112 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_112 <= _GEN_3707;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_113 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_113 <= _GEN_3708;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_114 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_114 <= _GEN_3709;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_115 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_115 <= _GEN_3710;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_116 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_116 <= _GEN_3711;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_117 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_117 <= _GEN_3712;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_118 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_118 <= _GEN_3713;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_119 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_119 <= _GEN_3714;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_120 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_120 <= _GEN_3715;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_121 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_121 <= _GEN_3716;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_122 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_122 <= _GEN_3717;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_123 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_123 <= _GEN_3718;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_124 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_124 <= _GEN_3719;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_125 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_125 <= _GEN_3720;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_126 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_126 <= _GEN_3721;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:32]
      record_wdata1_127 <= 64'h0; // @[d_cache.scala 21:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wdata1_127 <= _GEN_3722;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_0 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_0 <= _GEN_3723;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_1 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_1 <= _GEN_3724;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_2 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_2 <= _GEN_3725;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_3 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_3 <= _GEN_3726;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_4 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_4 <= _GEN_3727;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_5 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_5 <= _GEN_3728;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_6 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_6 <= _GEN_3729;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_7 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_7 <= _GEN_3730;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_8 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_8 <= _GEN_3731;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_9 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_9 <= _GEN_3732;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_10 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_10 <= _GEN_3733;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_11 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_11 <= _GEN_3734;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_12 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_12 <= _GEN_3735;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_13 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_13 <= _GEN_3736;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_14 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_14 <= _GEN_3737;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_15 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_15 <= _GEN_3738;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_16 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_16 <= _GEN_3739;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_17 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_17 <= _GEN_3740;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_18 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_18 <= _GEN_3741;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_19 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_19 <= _GEN_3742;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_20 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_20 <= _GEN_3743;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_21 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_21 <= _GEN_3744;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_22 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_22 <= _GEN_3745;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_23 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_23 <= _GEN_3746;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_24 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_24 <= _GEN_3747;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_25 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_25 <= _GEN_3748;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_26 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_26 <= _GEN_3749;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_27 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_27 <= _GEN_3750;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_28 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_28 <= _GEN_3751;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_29 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_29 <= _GEN_3752;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_30 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_30 <= _GEN_3753;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_31 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_31 <= _GEN_3754;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_32 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_32 <= _GEN_3755;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_33 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_33 <= _GEN_3756;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_34 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_34 <= _GEN_3757;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_35 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_35 <= _GEN_3758;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_36 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_36 <= _GEN_3759;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_37 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_37 <= _GEN_3760;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_38 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_38 <= _GEN_3761;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_39 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_39 <= _GEN_3762;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_40 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_40 <= _GEN_3763;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_41 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_41 <= _GEN_3764;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_42 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_42 <= _GEN_3765;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_43 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_43 <= _GEN_3766;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_44 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_44 <= _GEN_3767;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_45 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_45 <= _GEN_3768;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_46 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_46 <= _GEN_3769;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_47 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_47 <= _GEN_3770;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_48 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_48 <= _GEN_3771;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_49 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_49 <= _GEN_3772;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_50 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_50 <= _GEN_3773;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_51 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_51 <= _GEN_3774;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_52 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_52 <= _GEN_3775;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_53 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_53 <= _GEN_3776;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_54 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_54 <= _GEN_3777;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_55 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_55 <= _GEN_3778;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_56 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_56 <= _GEN_3779;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_57 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_57 <= _GEN_3780;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_58 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_58 <= _GEN_3781;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_59 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_59 <= _GEN_3782;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_60 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_60 <= _GEN_3783;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_61 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_61 <= _GEN_3784;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_62 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_62 <= _GEN_3785;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_63 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_63 <= _GEN_3786;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_64 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_64 <= _GEN_3787;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_65 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_65 <= _GEN_3788;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_66 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_66 <= _GEN_3789;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_67 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_67 <= _GEN_3790;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_68 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_68 <= _GEN_3791;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_69 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_69 <= _GEN_3792;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_70 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_70 <= _GEN_3793;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_71 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_71 <= _GEN_3794;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_72 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_72 <= _GEN_3795;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_73 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_73 <= _GEN_3796;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_74 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_74 <= _GEN_3797;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_75 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_75 <= _GEN_3798;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_76 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_76 <= _GEN_3799;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_77 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_77 <= _GEN_3800;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_78 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_78 <= _GEN_3801;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_79 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_79 <= _GEN_3802;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_80 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_80 <= _GEN_3803;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_81 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_81 <= _GEN_3804;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_82 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_82 <= _GEN_3805;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_83 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_83 <= _GEN_3806;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_84 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_84 <= _GEN_3807;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_85 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_85 <= _GEN_3808;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_86 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_86 <= _GEN_3809;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_87 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_87 <= _GEN_3810;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_88 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_88 <= _GEN_3811;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_89 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_89 <= _GEN_3812;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_90 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_90 <= _GEN_3813;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_91 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_91 <= _GEN_3814;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_92 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_92 <= _GEN_3815;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_93 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_93 <= _GEN_3816;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_94 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_94 <= _GEN_3817;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_95 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_95 <= _GEN_3818;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_96 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_96 <= _GEN_3819;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_97 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_97 <= _GEN_3820;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_98 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_98 <= _GEN_3821;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_99 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_99 <= _GEN_3822;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_100 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_100 <= _GEN_3823;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_101 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_101 <= _GEN_3824;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_102 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_102 <= _GEN_3825;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_103 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_103 <= _GEN_3826;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_104 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_104 <= _GEN_3827;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_105 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_105 <= _GEN_3828;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_106 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_106 <= _GEN_3829;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_107 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_107 <= _GEN_3830;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_108 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_108 <= _GEN_3831;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_109 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_109 <= _GEN_3832;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_110 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_110 <= _GEN_3833;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_111 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_111 <= _GEN_3834;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_112 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_112 <= _GEN_3835;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_113 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_113 <= _GEN_3836;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_114 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_114 <= _GEN_3837;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_115 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_115 <= _GEN_3838;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_116 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_116 <= _GEN_3839;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_117 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_117 <= _GEN_3840;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_118 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_118 <= _GEN_3841;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_119 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_119 <= _GEN_3842;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_120 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_120 <= _GEN_3843;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_121 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_121 <= _GEN_3844;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_122 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_122 <= _GEN_3845;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_123 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_123 <= _GEN_3846;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_124 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_124 <= _GEN_3847;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_125 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_125 <= _GEN_3848;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_126 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_126 <= _GEN_3849;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:32]
      record_wstrb1_127 <= 8'h0; // @[d_cache.scala 22:32]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_wstrb1_127 <= _GEN_3850;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_0 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_0 <= _GEN_3851;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_1 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_1 <= _GEN_3852;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_2 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_2 <= _GEN_3853;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_3 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_3 <= _GEN_3854;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_4 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_4 <= _GEN_3855;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_5 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_5 <= _GEN_3856;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_6 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_6 <= _GEN_3857;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_7 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_7 <= _GEN_3858;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_8 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_8 <= _GEN_3859;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_9 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_9 <= _GEN_3860;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_10 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_10 <= _GEN_3861;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_11 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_11 <= _GEN_3862;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_12 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_12 <= _GEN_3863;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_13 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_13 <= _GEN_3864;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_14 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_14 <= _GEN_3865;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_15 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_15 <= _GEN_3866;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_16 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_16 <= _GEN_3867;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_17 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_17 <= _GEN_3868;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_18 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_18 <= _GEN_3869;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_19 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_19 <= _GEN_3870;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_20 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_20 <= _GEN_3871;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_21 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_21 <= _GEN_3872;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_22 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_22 <= _GEN_3873;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_23 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_23 <= _GEN_3874;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_24 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_24 <= _GEN_3875;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_25 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_25 <= _GEN_3876;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_26 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_26 <= _GEN_3877;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_27 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_27 <= _GEN_3878;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_28 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_28 <= _GEN_3879;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_29 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_29 <= _GEN_3880;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_30 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_30 <= _GEN_3881;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_31 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_31 <= _GEN_3882;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_32 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_32 <= _GEN_3883;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_33 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_33 <= _GEN_3884;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_34 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_34 <= _GEN_3885;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_35 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_35 <= _GEN_3886;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_36 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_36 <= _GEN_3887;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_37 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_37 <= _GEN_3888;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_38 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_38 <= _GEN_3889;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_39 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_39 <= _GEN_3890;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_40 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_40 <= _GEN_3891;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_41 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_41 <= _GEN_3892;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_42 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_42 <= _GEN_3893;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_43 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_43 <= _GEN_3894;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_44 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_44 <= _GEN_3895;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_45 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_45 <= _GEN_3896;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_46 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_46 <= _GEN_3897;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_47 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_47 <= _GEN_3898;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_48 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_48 <= _GEN_3899;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_49 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_49 <= _GEN_3900;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_50 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_50 <= _GEN_3901;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_51 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_51 <= _GEN_3902;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_52 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_52 <= _GEN_3903;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_53 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_53 <= _GEN_3904;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_54 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_54 <= _GEN_3905;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_55 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_55 <= _GEN_3906;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_56 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_56 <= _GEN_3907;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_57 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_57 <= _GEN_3908;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_58 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_58 <= _GEN_3909;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_59 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_59 <= _GEN_3910;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_60 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_60 <= _GEN_3911;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_61 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_61 <= _GEN_3912;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_62 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_62 <= _GEN_3913;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_63 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_63 <= _GEN_3914;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_64 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_64 <= _GEN_3915;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_65 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_65 <= _GEN_3916;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_66 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_66 <= _GEN_3917;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_67 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_67 <= _GEN_3918;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_68 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_68 <= _GEN_3919;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_69 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_69 <= _GEN_3920;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_70 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_70 <= _GEN_3921;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_71 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_71 <= _GEN_3922;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_72 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_72 <= _GEN_3923;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_73 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_73 <= _GEN_3924;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_74 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_74 <= _GEN_3925;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_75 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_75 <= _GEN_3926;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_76 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_76 <= _GEN_3927;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_77 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_77 <= _GEN_3928;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_78 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_78 <= _GEN_3929;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_79 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_79 <= _GEN_3930;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_80 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_80 <= _GEN_3931;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_81 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_81 <= _GEN_3932;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_82 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_82 <= _GEN_3933;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_83 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_83 <= _GEN_3934;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_84 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_84 <= _GEN_3935;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_85 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_85 <= _GEN_3936;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_86 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_86 <= _GEN_3937;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_87 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_87 <= _GEN_3938;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_88 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_88 <= _GEN_3939;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_89 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_89 <= _GEN_3940;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_90 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_90 <= _GEN_3941;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_91 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_91 <= _GEN_3942;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_92 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_92 <= _GEN_3943;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_93 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_93 <= _GEN_3944;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_94 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_94 <= _GEN_3945;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_95 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_95 <= _GEN_3946;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_96 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_96 <= _GEN_3947;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_97 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_97 <= _GEN_3948;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_98 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_98 <= _GEN_3949;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_99 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_99 <= _GEN_3950;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_100 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_100 <= _GEN_3951;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_101 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_101 <= _GEN_3952;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_102 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_102 <= _GEN_3953;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_103 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_103 <= _GEN_3954;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_104 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_104 <= _GEN_3955;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_105 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_105 <= _GEN_3956;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_106 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_106 <= _GEN_3957;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_107 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_107 <= _GEN_3958;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_108 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_108 <= _GEN_3959;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_109 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_109 <= _GEN_3960;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_110 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_110 <= _GEN_3961;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_111 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_111 <= _GEN_3962;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_112 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_112 <= _GEN_3963;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_113 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_113 <= _GEN_3964;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_114 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_114 <= _GEN_3965;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_115 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_115 <= _GEN_3966;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_116 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_116 <= _GEN_3967;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_117 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_117 <= _GEN_3968;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_118 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_118 <= _GEN_3969;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_119 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_119 <= _GEN_3970;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_120 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_120 <= _GEN_3971;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_121 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_121 <= _GEN_3972;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_122 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_122 <= _GEN_3973;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_123 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_123 <= _GEN_3974;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_124 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_124 <= _GEN_3975;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_125 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_125 <= _GEN_3976;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_126 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_126 <= _GEN_3977;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:28]
      record_pc_127 <= 64'h0; // @[d_cache.scala 23:28]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_pc_127 <= _GEN_3978;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_0 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_0 <= _GEN_3979;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_1 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_1 <= _GEN_3980;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_2 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_2 <= _GEN_3981;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_3 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_3 <= _GEN_3982;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_4 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_4 <= _GEN_3983;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_5 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_5 <= _GEN_3984;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_6 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_6 <= _GEN_3985;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_7 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_7 <= _GEN_3986;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_8 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_8 <= _GEN_3987;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_9 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_9 <= _GEN_3988;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_10 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_10 <= _GEN_3989;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_11 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_11 <= _GEN_3990;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_12 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_12 <= _GEN_3991;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_13 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_13 <= _GEN_3992;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_14 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_14 <= _GEN_3993;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_15 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_15 <= _GEN_3994;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_16 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_16 <= _GEN_3995;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_17 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_17 <= _GEN_3996;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_18 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_18 <= _GEN_3997;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_19 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_19 <= _GEN_3998;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_20 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_20 <= _GEN_3999;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_21 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_21 <= _GEN_4000;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_22 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_22 <= _GEN_4001;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_23 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_23 <= _GEN_4002;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_24 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_24 <= _GEN_4003;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_25 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_25 <= _GEN_4004;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_26 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_26 <= _GEN_4005;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_27 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_27 <= _GEN_4006;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_28 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_28 <= _GEN_4007;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_29 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_29 <= _GEN_4008;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_30 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_30 <= _GEN_4009;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_31 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_31 <= _GEN_4010;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_32 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_32 <= _GEN_4011;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_33 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_33 <= _GEN_4012;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_34 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_34 <= _GEN_4013;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_35 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_35 <= _GEN_4014;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_36 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_36 <= _GEN_4015;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_37 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_37 <= _GEN_4016;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_38 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_38 <= _GEN_4017;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_39 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_39 <= _GEN_4018;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_40 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_40 <= _GEN_4019;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_41 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_41 <= _GEN_4020;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_42 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_42 <= _GEN_4021;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_43 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_43 <= _GEN_4022;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_44 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_44 <= _GEN_4023;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_45 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_45 <= _GEN_4024;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_46 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_46 <= _GEN_4025;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_47 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_47 <= _GEN_4026;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_48 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_48 <= _GEN_4027;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_49 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_49 <= _GEN_4028;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_50 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_50 <= _GEN_4029;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_51 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_51 <= _GEN_4030;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_52 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_52 <= _GEN_4031;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_53 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_53 <= _GEN_4032;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_54 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_54 <= _GEN_4033;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_55 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_55 <= _GEN_4034;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_56 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_56 <= _GEN_4035;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_57 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_57 <= _GEN_4036;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_58 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_58 <= _GEN_4037;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_59 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_59 <= _GEN_4038;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_60 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_60 <= _GEN_4039;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_61 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_61 <= _GEN_4040;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_62 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_62 <= _GEN_4041;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_63 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_63 <= _GEN_4042;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_64 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_64 <= _GEN_4043;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_65 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_65 <= _GEN_4044;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_66 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_66 <= _GEN_4045;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_67 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_67 <= _GEN_4046;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_68 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_68 <= _GEN_4047;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_69 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_69 <= _GEN_4048;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_70 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_70 <= _GEN_4049;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_71 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_71 <= _GEN_4050;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_72 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_72 <= _GEN_4051;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_73 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_73 <= _GEN_4052;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_74 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_74 <= _GEN_4053;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_75 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_75 <= _GEN_4054;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_76 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_76 <= _GEN_4055;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_77 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_77 <= _GEN_4056;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_78 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_78 <= _GEN_4057;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_79 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_79 <= _GEN_4058;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_80 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_80 <= _GEN_4059;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_81 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_81 <= _GEN_4060;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_82 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_82 <= _GEN_4061;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_83 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_83 <= _GEN_4062;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_84 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_84 <= _GEN_4063;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_85 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_85 <= _GEN_4064;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_86 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_86 <= _GEN_4065;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_87 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_87 <= _GEN_4066;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_88 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_88 <= _GEN_4067;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_89 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_89 <= _GEN_4068;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_90 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_90 <= _GEN_4069;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_91 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_91 <= _GEN_4070;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_92 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_92 <= _GEN_4071;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_93 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_93 <= _GEN_4072;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_94 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_94 <= _GEN_4073;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_95 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_95 <= _GEN_4074;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_96 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_96 <= _GEN_4075;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_97 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_97 <= _GEN_4076;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_98 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_98 <= _GEN_4077;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_99 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_99 <= _GEN_4078;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_100 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_100 <= _GEN_4079;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_101 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_101 <= _GEN_4080;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_102 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_102 <= _GEN_4081;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_103 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_103 <= _GEN_4082;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_104 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_104 <= _GEN_4083;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_105 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_105 <= _GEN_4084;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_106 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_106 <= _GEN_4085;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_107 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_107 <= _GEN_4086;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_108 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_108 <= _GEN_4087;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_109 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_109 <= _GEN_4088;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_110 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_110 <= _GEN_4089;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_111 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_111 <= _GEN_4090;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_112 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_112 <= _GEN_4091;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_113 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_113 <= _GEN_4092;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_114 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_114 <= _GEN_4093;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_115 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_115 <= _GEN_4094;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_116 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_116 <= _GEN_4095;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_117 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_117 <= _GEN_4096;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_118 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_118 <= _GEN_4097;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_119 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_119 <= _GEN_4098;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_120 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_120 <= _GEN_4099;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_121 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_121 <= _GEN_4100;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_122 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_122 <= _GEN_4101;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_123 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_123 <= _GEN_4102;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_124 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_124 <= _GEN_4103;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_125 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_125 <= _GEN_4104;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_126 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_126 <= _GEN_4105;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:30]
      record_addr_127 <= 32'h0; // @[d_cache.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_addr_127 <= _GEN_4106;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_0 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_0 <= _GEN_3339;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_1 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_1 <= _GEN_3340;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_2 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_2 <= _GEN_3341;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_3 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_3 <= _GEN_3342;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_4 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_4 <= _GEN_3343;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_5 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_5 <= _GEN_3344;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_6 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_6 <= _GEN_3345;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_7 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_7 <= _GEN_3346;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_8 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_8 <= _GEN_3347;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_9 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_9 <= _GEN_3348;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_10 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_10 <= _GEN_3349;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_11 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_11 <= _GEN_3350;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_12 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_12 <= _GEN_3351;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_13 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_13 <= _GEN_3352;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_14 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_14 <= _GEN_3353;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_15 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_15 <= _GEN_3354;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_16 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_16 <= _GEN_3355;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_17 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_17 <= _GEN_3356;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_18 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_18 <= _GEN_3357;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_19 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_19 <= _GEN_3358;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_20 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_20 <= _GEN_3359;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_21 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_21 <= _GEN_3360;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_22 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_22 <= _GEN_3361;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_23 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_23 <= _GEN_3362;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_24 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_24 <= _GEN_3363;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_25 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_25 <= _GEN_3364;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_26 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_26 <= _GEN_3365;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_27 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_27 <= _GEN_3366;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_28 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_28 <= _GEN_3367;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_29 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_29 <= _GEN_3368;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_30 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_30 <= _GEN_3369;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_31 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_31 <= _GEN_3370;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_32 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_32 <= _GEN_3371;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_33 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_33 <= _GEN_3372;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_34 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_34 <= _GEN_3373;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_35 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_35 <= _GEN_3374;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_36 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_36 <= _GEN_3375;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_37 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_37 <= _GEN_3376;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_38 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_38 <= _GEN_3377;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_39 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_39 <= _GEN_3378;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_40 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_40 <= _GEN_3379;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_41 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_41 <= _GEN_3380;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_42 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_42 <= _GEN_3381;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_43 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_43 <= _GEN_3382;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_44 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_44 <= _GEN_3383;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_45 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_45 <= _GEN_3384;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_46 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_46 <= _GEN_3385;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_47 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_47 <= _GEN_3386;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_48 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_48 <= _GEN_3387;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_49 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_49 <= _GEN_3388;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_50 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_50 <= _GEN_3389;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_51 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_51 <= _GEN_3390;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_52 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_52 <= _GEN_3391;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_53 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_53 <= _GEN_3392;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_54 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_54 <= _GEN_3393;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_55 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_55 <= _GEN_3394;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_56 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_56 <= _GEN_3395;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_57 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_57 <= _GEN_3396;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_58 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_58 <= _GEN_3397;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_59 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_59 <= _GEN_3398;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_60 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_60 <= _GEN_3399;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_61 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_61 <= _GEN_3400;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_62 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_62 <= _GEN_3401;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_63 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_63 <= _GEN_3402;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_64 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_64 <= _GEN_3403;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_65 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_65 <= _GEN_3404;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_66 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_66 <= _GEN_3405;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_67 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_67 <= _GEN_3406;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_68 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_68 <= _GEN_3407;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_69 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_69 <= _GEN_3408;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_70 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_70 <= _GEN_3409;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_71 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_71 <= _GEN_3410;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_72 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_72 <= _GEN_3411;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_73 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_73 <= _GEN_3412;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_74 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_74 <= _GEN_3413;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_75 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_75 <= _GEN_3414;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_76 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_76 <= _GEN_3415;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_77 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_77 <= _GEN_3416;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_78 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_78 <= _GEN_3417;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_79 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_79 <= _GEN_3418;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_80 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_80 <= _GEN_3419;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_81 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_81 <= _GEN_3420;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_82 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_82 <= _GEN_3421;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_83 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_83 <= _GEN_3422;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_84 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_84 <= _GEN_3423;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_85 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_85 <= _GEN_3424;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_86 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_86 <= _GEN_3425;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_87 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_87 <= _GEN_3426;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_88 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_88 <= _GEN_3427;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_89 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_89 <= _GEN_3428;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_90 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_90 <= _GEN_3429;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_91 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_91 <= _GEN_3430;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_92 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_92 <= _GEN_3431;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_93 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_93 <= _GEN_3432;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_94 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_94 <= _GEN_3433;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_95 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_95 <= _GEN_3434;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_96 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_96 <= _GEN_3435;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_97 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_97 <= _GEN_3436;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_98 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_98 <= _GEN_3437;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_99 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_99 <= _GEN_3438;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_100 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_100 <= _GEN_3439;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_101 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_101 <= _GEN_3440;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_102 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_102 <= _GEN_3441;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_103 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_103 <= _GEN_3442;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_104 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_104 <= _GEN_3443;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_105 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_105 <= _GEN_3444;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_106 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_106 <= _GEN_3445;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_107 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_107 <= _GEN_3446;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_108 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_108 <= _GEN_3447;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_109 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_109 <= _GEN_3448;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_110 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_110 <= _GEN_3449;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_111 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_111 <= _GEN_3450;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_112 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_112 <= _GEN_3451;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_113 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_113 <= _GEN_3452;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_114 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_114 <= _GEN_3453;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_115 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_115 <= _GEN_3454;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_116 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_116 <= _GEN_3455;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_117 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_117 <= _GEN_3456;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_118 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_118 <= _GEN_3457;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_119 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_119 <= _GEN_3458;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_120 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_120 <= _GEN_3459;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_121 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_121 <= _GEN_3460;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_122 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_122 <= _GEN_3461;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_123 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_123 <= _GEN_3462;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_124 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_124 <= _GEN_3463;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_125 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_125 <= _GEN_3464;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_126 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_126 <= _GEN_3465;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:33]
      record_olddata_127 <= 64'h0; // @[d_cache.scala 25:33]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          record_olddata_127 <= _GEN_3466;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_0 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_0 <= _GEN_13103;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_1 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_1 <= _GEN_13104;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_2 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_2 <= _GEN_13105;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_3 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_3 <= _GEN_13106;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_4 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_4 <= _GEN_13107;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_5 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_5 <= _GEN_13108;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_6 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_6 <= _GEN_13109;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_7 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_7 <= _GEN_13110;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_8 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_8 <= _GEN_13111;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_9 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_9 <= _GEN_13112;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_10 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_10 <= _GEN_13113;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_11 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_11 <= _GEN_13114;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_12 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_12 <= _GEN_13115;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_13 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_13 <= _GEN_13116;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_14 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_14 <= _GEN_13117;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_15 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_15 <= _GEN_13118;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_16 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_16 <= _GEN_13119;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_17 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_17 <= _GEN_13120;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_18 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_18 <= _GEN_13121;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_19 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_19 <= _GEN_13122;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_20 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_20 <= _GEN_13123;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_21 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_21 <= _GEN_13124;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_22 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_22 <= _GEN_13125;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_23 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_23 <= _GEN_13126;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_24 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_24 <= _GEN_13127;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_25 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_25 <= _GEN_13128;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_26 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_26 <= _GEN_13129;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_27 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_27 <= _GEN_13130;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_28 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_28 <= _GEN_13131;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_29 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_29 <= _GEN_13132;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_30 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_30 <= _GEN_13133;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_31 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_31 <= _GEN_13134;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_32 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_32 <= _GEN_13135;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_33 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_33 <= _GEN_13136;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_34 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_34 <= _GEN_13137;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_35 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_35 <= _GEN_13138;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_36 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_36 <= _GEN_13139;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_37 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_37 <= _GEN_13140;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_38 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_38 <= _GEN_13141;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_39 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_39 <= _GEN_13142;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_40 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_40 <= _GEN_13143;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_41 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_41 <= _GEN_13144;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_42 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_42 <= _GEN_13145;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_43 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_43 <= _GEN_13146;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_44 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_44 <= _GEN_13147;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_45 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_45 <= _GEN_13148;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_46 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_46 <= _GEN_13149;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_47 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_47 <= _GEN_13150;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_48 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_48 <= _GEN_13151;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_49 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_49 <= _GEN_13152;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_50 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_50 <= _GEN_13153;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_51 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_51 <= _GEN_13154;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_52 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_52 <= _GEN_13155;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_53 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_53 <= _GEN_13156;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_54 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_54 <= _GEN_13157;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_55 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_55 <= _GEN_13158;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_56 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_56 <= _GEN_13159;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_57 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_57 <= _GEN_13160;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_58 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_58 <= _GEN_13161;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_59 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_59 <= _GEN_13162;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_60 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_60 <= _GEN_13163;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_61 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_61 <= _GEN_13164;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_62 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_62 <= _GEN_13165;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_63 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_63 <= _GEN_13166;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_64 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_64 <= _GEN_13167;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_65 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_65 <= _GEN_13168;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_66 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_66 <= _GEN_13169;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_67 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_67 <= _GEN_13170;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_68 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_68 <= _GEN_13171;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_69 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_69 <= _GEN_13172;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_70 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_70 <= _GEN_13173;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_71 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_71 <= _GEN_13174;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_72 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_72 <= _GEN_13175;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_73 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_73 <= _GEN_13176;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_74 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_74 <= _GEN_13177;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_75 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_75 <= _GEN_13178;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_76 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_76 <= _GEN_13179;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_77 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_77 <= _GEN_13180;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_78 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_78 <= _GEN_13181;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_79 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_79 <= _GEN_13182;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_80 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_80 <= _GEN_13183;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_81 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_81 <= _GEN_13184;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_82 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_82 <= _GEN_13185;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_83 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_83 <= _GEN_13186;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_84 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_84 <= _GEN_13187;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_85 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_85 <= _GEN_13188;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_86 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_86 <= _GEN_13189;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_87 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_87 <= _GEN_13190;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_88 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_88 <= _GEN_13191;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_89 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_89 <= _GEN_13192;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_90 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_90 <= _GEN_13193;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_91 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_91 <= _GEN_13194;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_92 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_92 <= _GEN_13195;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_93 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_93 <= _GEN_13196;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_94 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_94 <= _GEN_13197;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_95 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_95 <= _GEN_13198;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_96 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_96 <= _GEN_13199;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_97 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_97 <= _GEN_13200;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_98 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_98 <= _GEN_13201;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_99 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_99 <= _GEN_13202;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_100 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_100 <= _GEN_13203;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_101 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_101 <= _GEN_13204;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_102 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_102 <= _GEN_13205;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_103 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_103 <= _GEN_13206;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_104 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_104 <= _GEN_13207;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_105 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_105 <= _GEN_13208;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_106 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_106 <= _GEN_13209;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_107 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_107 <= _GEN_13210;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_108 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_108 <= _GEN_13211;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_109 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_109 <= _GEN_13212;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_110 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_110 <= _GEN_13213;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_111 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_111 <= _GEN_13214;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_112 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_112 <= _GEN_13215;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_113 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_113 <= _GEN_13216;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_114 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_114 <= _GEN_13217;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_115 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_115 <= _GEN_13218;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_116 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_116 <= _GEN_13219;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_117 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_117 <= _GEN_13220;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_118 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_118 <= _GEN_13221;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_119 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_119 <= _GEN_13222;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_120 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_120 <= _GEN_13223;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_121 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_121 <= _GEN_13224;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_122 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_122 <= _GEN_13225;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_123 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_123 <= _GEN_13226;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_124 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_124 <= _GEN_13227;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_125 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_125 <= _GEN_13228;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_126 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_126 <= _GEN_13229;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:24]
      tag_0_127 <= 32'h0; // @[d_cache.scala 28:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_127 <= _GEN_13230;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_0 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_0 <= _GEN_13488;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_1 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_1 <= _GEN_13489;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_2 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_2 <= _GEN_13490;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_3 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_3 <= _GEN_13491;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_4 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_4 <= _GEN_13492;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_5 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_5 <= _GEN_13493;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_6 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_6 <= _GEN_13494;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_7 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_7 <= _GEN_13495;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_8 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_8 <= _GEN_13496;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_9 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_9 <= _GEN_13497;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_10 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_10 <= _GEN_13498;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_11 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_11 <= _GEN_13499;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_12 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_12 <= _GEN_13500;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_13 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_13 <= _GEN_13501;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_14 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_14 <= _GEN_13502;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_15 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_15 <= _GEN_13503;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_16 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_16 <= _GEN_13504;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_17 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_17 <= _GEN_13505;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_18 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_18 <= _GEN_13506;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_19 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_19 <= _GEN_13507;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_20 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_20 <= _GEN_13508;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_21 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_21 <= _GEN_13509;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_22 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_22 <= _GEN_13510;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_23 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_23 <= _GEN_13511;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_24 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_24 <= _GEN_13512;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_25 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_25 <= _GEN_13513;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_26 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_26 <= _GEN_13514;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_27 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_27 <= _GEN_13515;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_28 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_28 <= _GEN_13516;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_29 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_29 <= _GEN_13517;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_30 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_30 <= _GEN_13518;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_31 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_31 <= _GEN_13519;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_32 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_32 <= _GEN_13520;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_33 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_33 <= _GEN_13521;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_34 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_34 <= _GEN_13522;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_35 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_35 <= _GEN_13523;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_36 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_36 <= _GEN_13524;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_37 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_37 <= _GEN_13525;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_38 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_38 <= _GEN_13526;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_39 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_39 <= _GEN_13527;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_40 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_40 <= _GEN_13528;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_41 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_41 <= _GEN_13529;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_42 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_42 <= _GEN_13530;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_43 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_43 <= _GEN_13531;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_44 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_44 <= _GEN_13532;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_45 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_45 <= _GEN_13533;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_46 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_46 <= _GEN_13534;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_47 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_47 <= _GEN_13535;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_48 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_48 <= _GEN_13536;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_49 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_49 <= _GEN_13537;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_50 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_50 <= _GEN_13538;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_51 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_51 <= _GEN_13539;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_52 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_52 <= _GEN_13540;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_53 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_53 <= _GEN_13541;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_54 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_54 <= _GEN_13542;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_55 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_55 <= _GEN_13543;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_56 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_56 <= _GEN_13544;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_57 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_57 <= _GEN_13545;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_58 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_58 <= _GEN_13546;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_59 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_59 <= _GEN_13547;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_60 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_60 <= _GEN_13548;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_61 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_61 <= _GEN_13549;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_62 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_62 <= _GEN_13550;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_63 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_63 <= _GEN_13551;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_64 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_64 <= _GEN_13552;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_65 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_65 <= _GEN_13553;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_66 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_66 <= _GEN_13554;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_67 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_67 <= _GEN_13555;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_68 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_68 <= _GEN_13556;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_69 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_69 <= _GEN_13557;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_70 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_70 <= _GEN_13558;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_71 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_71 <= _GEN_13559;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_72 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_72 <= _GEN_13560;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_73 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_73 <= _GEN_13561;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_74 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_74 <= _GEN_13562;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_75 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_75 <= _GEN_13563;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_76 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_76 <= _GEN_13564;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_77 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_77 <= _GEN_13565;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_78 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_78 <= _GEN_13566;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_79 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_79 <= _GEN_13567;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_80 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_80 <= _GEN_13568;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_81 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_81 <= _GEN_13569;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_82 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_82 <= _GEN_13570;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_83 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_83 <= _GEN_13571;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_84 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_84 <= _GEN_13572;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_85 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_85 <= _GEN_13573;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_86 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_86 <= _GEN_13574;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_87 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_87 <= _GEN_13575;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_88 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_88 <= _GEN_13576;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_89 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_89 <= _GEN_13577;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_90 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_90 <= _GEN_13578;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_91 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_91 <= _GEN_13579;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_92 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_92 <= _GEN_13580;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_93 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_93 <= _GEN_13581;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_94 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_94 <= _GEN_13582;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_95 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_95 <= _GEN_13583;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_96 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_96 <= _GEN_13584;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_97 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_97 <= _GEN_13585;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_98 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_98 <= _GEN_13586;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_99 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_99 <= _GEN_13587;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_100 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_100 <= _GEN_13588;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_101 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_101 <= _GEN_13589;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_102 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_102 <= _GEN_13590;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_103 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_103 <= _GEN_13591;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_104 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_104 <= _GEN_13592;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_105 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_105 <= _GEN_13593;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_106 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_106 <= _GEN_13594;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_107 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_107 <= _GEN_13595;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_108 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_108 <= _GEN_13596;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_109 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_109 <= _GEN_13597;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_110 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_110 <= _GEN_13598;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_111 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_111 <= _GEN_13599;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_112 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_112 <= _GEN_13600;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_113 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_113 <= _GEN_13601;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_114 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_114 <= _GEN_13602;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_115 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_115 <= _GEN_13603;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_116 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_116 <= _GEN_13604;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_117 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_117 <= _GEN_13605;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_118 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_118 <= _GEN_13606;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_119 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_119 <= _GEN_13607;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_120 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_120 <= _GEN_13608;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_121 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_121 <= _GEN_13609;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_122 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_122 <= _GEN_13610;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_123 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_123 <= _GEN_13611;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_124 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_124 <= _GEN_13612;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_125 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_125 <= _GEN_13613;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_126 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_126 <= _GEN_13614;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:24]
      tag_1_127 <= 32'h0; // @[d_cache.scala 29:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_127 <= _GEN_13615;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_0 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_0 <= _GEN_13231;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_1 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_1 <= _GEN_13232;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_2 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_2 <= _GEN_13233;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_3 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_3 <= _GEN_13234;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_4 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_4 <= _GEN_13235;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_5 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_5 <= _GEN_13236;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_6 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_6 <= _GEN_13237;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_7 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_7 <= _GEN_13238;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_8 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_8 <= _GEN_13239;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_9 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_9 <= _GEN_13240;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_10 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_10 <= _GEN_13241;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_11 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_11 <= _GEN_13242;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_12 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_12 <= _GEN_13243;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_13 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_13 <= _GEN_13244;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_14 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_14 <= _GEN_13245;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_15 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_15 <= _GEN_13246;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_16 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_16 <= _GEN_13247;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_17 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_17 <= _GEN_13248;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_18 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_18 <= _GEN_13249;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_19 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_19 <= _GEN_13250;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_20 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_20 <= _GEN_13251;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_21 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_21 <= _GEN_13252;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_22 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_22 <= _GEN_13253;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_23 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_23 <= _GEN_13254;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_24 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_24 <= _GEN_13255;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_25 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_25 <= _GEN_13256;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_26 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_26 <= _GEN_13257;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_27 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_27 <= _GEN_13258;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_28 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_28 <= _GEN_13259;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_29 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_29 <= _GEN_13260;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_30 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_30 <= _GEN_13261;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_31 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_31 <= _GEN_13262;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_32 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_32 <= _GEN_13263;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_33 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_33 <= _GEN_13264;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_34 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_34 <= _GEN_13265;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_35 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_35 <= _GEN_13266;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_36 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_36 <= _GEN_13267;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_37 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_37 <= _GEN_13268;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_38 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_38 <= _GEN_13269;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_39 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_39 <= _GEN_13270;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_40 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_40 <= _GEN_13271;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_41 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_41 <= _GEN_13272;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_42 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_42 <= _GEN_13273;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_43 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_43 <= _GEN_13274;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_44 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_44 <= _GEN_13275;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_45 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_45 <= _GEN_13276;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_46 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_46 <= _GEN_13277;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_47 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_47 <= _GEN_13278;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_48 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_48 <= _GEN_13279;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_49 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_49 <= _GEN_13280;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_50 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_50 <= _GEN_13281;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_51 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_51 <= _GEN_13282;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_52 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_52 <= _GEN_13283;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_53 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_53 <= _GEN_13284;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_54 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_54 <= _GEN_13285;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_55 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_55 <= _GEN_13286;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_56 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_56 <= _GEN_13287;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_57 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_57 <= _GEN_13288;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_58 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_58 <= _GEN_13289;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_59 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_59 <= _GEN_13290;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_60 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_60 <= _GEN_13291;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_61 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_61 <= _GEN_13292;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_62 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_62 <= _GEN_13293;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_63 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_63 <= _GEN_13294;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_64 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_64 <= _GEN_13295;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_65 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_65 <= _GEN_13296;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_66 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_66 <= _GEN_13297;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_67 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_67 <= _GEN_13298;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_68 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_68 <= _GEN_13299;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_69 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_69 <= _GEN_13300;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_70 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_70 <= _GEN_13301;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_71 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_71 <= _GEN_13302;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_72 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_72 <= _GEN_13303;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_73 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_73 <= _GEN_13304;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_74 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_74 <= _GEN_13305;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_75 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_75 <= _GEN_13306;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_76 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_76 <= _GEN_13307;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_77 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_77 <= _GEN_13308;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_78 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_78 <= _GEN_13309;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_79 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_79 <= _GEN_13310;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_80 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_80 <= _GEN_13311;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_81 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_81 <= _GEN_13312;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_82 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_82 <= _GEN_13313;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_83 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_83 <= _GEN_13314;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_84 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_84 <= _GEN_13315;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_85 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_85 <= _GEN_13316;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_86 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_86 <= _GEN_13317;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_87 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_87 <= _GEN_13318;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_88 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_88 <= _GEN_13319;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_89 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_89 <= _GEN_13320;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_90 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_90 <= _GEN_13321;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_91 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_91 <= _GEN_13322;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_92 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_92 <= _GEN_13323;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_93 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_93 <= _GEN_13324;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_94 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_94 <= _GEN_13325;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_95 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_95 <= _GEN_13326;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_96 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_96 <= _GEN_13327;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_97 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_97 <= _GEN_13328;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_98 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_98 <= _GEN_13329;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_99 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_99 <= _GEN_13330;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_100 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_100 <= _GEN_13331;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_101 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_101 <= _GEN_13332;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_102 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_102 <= _GEN_13333;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_103 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_103 <= _GEN_13334;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_104 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_104 <= _GEN_13335;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_105 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_105 <= _GEN_13336;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_106 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_106 <= _GEN_13337;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_107 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_107 <= _GEN_13338;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_108 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_108 <= _GEN_13339;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_109 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_109 <= _GEN_13340;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_110 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_110 <= _GEN_13341;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_111 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_111 <= _GEN_13342;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_112 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_112 <= _GEN_13343;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_113 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_113 <= _GEN_13344;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_114 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_114 <= _GEN_13345;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_115 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_115 <= _GEN_13346;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_116 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_116 <= _GEN_13347;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_117 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_117 <= _GEN_13348;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_118 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_118 <= _GEN_13349;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_119 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_119 <= _GEN_13350;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_120 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_120 <= _GEN_13351;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_121 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_121 <= _GEN_13352;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_122 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_122 <= _GEN_13353;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_123 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_123 <= _GEN_13354;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_124 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_124 <= _GEN_13355;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_125 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_125 <= _GEN_13356;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_126 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_126 <= _GEN_13357;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_0_127 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_127 <= _GEN_13358;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_0 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_0 <= _GEN_13616;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_1 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_1 <= _GEN_13617;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_2 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_2 <= _GEN_13618;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_3 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_3 <= _GEN_13619;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_4 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_4 <= _GEN_13620;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_5 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_5 <= _GEN_13621;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_6 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_6 <= _GEN_13622;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_7 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_7 <= _GEN_13623;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_8 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_8 <= _GEN_13624;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_9 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_9 <= _GEN_13625;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_10 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_10 <= _GEN_13626;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_11 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_11 <= _GEN_13627;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_12 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_12 <= _GEN_13628;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_13 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_13 <= _GEN_13629;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_14 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_14 <= _GEN_13630;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_15 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_15 <= _GEN_13631;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_16 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_16 <= _GEN_13632;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_17 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_17 <= _GEN_13633;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_18 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_18 <= _GEN_13634;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_19 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_19 <= _GEN_13635;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_20 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_20 <= _GEN_13636;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_21 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_21 <= _GEN_13637;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_22 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_22 <= _GEN_13638;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_23 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_23 <= _GEN_13639;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_24 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_24 <= _GEN_13640;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_25 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_25 <= _GEN_13641;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_26 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_26 <= _GEN_13642;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_27 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_27 <= _GEN_13643;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_28 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_28 <= _GEN_13644;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_29 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_29 <= _GEN_13645;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_30 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_30 <= _GEN_13646;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_31 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_31 <= _GEN_13647;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_32 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_32 <= _GEN_13648;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_33 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_33 <= _GEN_13649;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_34 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_34 <= _GEN_13650;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_35 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_35 <= _GEN_13651;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_36 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_36 <= _GEN_13652;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_37 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_37 <= _GEN_13653;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_38 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_38 <= _GEN_13654;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_39 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_39 <= _GEN_13655;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_40 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_40 <= _GEN_13656;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_41 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_41 <= _GEN_13657;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_42 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_42 <= _GEN_13658;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_43 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_43 <= _GEN_13659;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_44 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_44 <= _GEN_13660;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_45 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_45 <= _GEN_13661;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_46 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_46 <= _GEN_13662;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_47 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_47 <= _GEN_13663;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_48 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_48 <= _GEN_13664;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_49 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_49 <= _GEN_13665;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_50 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_50 <= _GEN_13666;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_51 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_51 <= _GEN_13667;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_52 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_52 <= _GEN_13668;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_53 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_53 <= _GEN_13669;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_54 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_54 <= _GEN_13670;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_55 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_55 <= _GEN_13671;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_56 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_56 <= _GEN_13672;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_57 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_57 <= _GEN_13673;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_58 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_58 <= _GEN_13674;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_59 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_59 <= _GEN_13675;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_60 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_60 <= _GEN_13676;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_61 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_61 <= _GEN_13677;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_62 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_62 <= _GEN_13678;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_63 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_63 <= _GEN_13679;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_64 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_64 <= _GEN_13680;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_65 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_65 <= _GEN_13681;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_66 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_66 <= _GEN_13682;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_67 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_67 <= _GEN_13683;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_68 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_68 <= _GEN_13684;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_69 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_69 <= _GEN_13685;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_70 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_70 <= _GEN_13686;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_71 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_71 <= _GEN_13687;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_72 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_72 <= _GEN_13688;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_73 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_73 <= _GEN_13689;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_74 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_74 <= _GEN_13690;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_75 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_75 <= _GEN_13691;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_76 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_76 <= _GEN_13692;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_77 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_77 <= _GEN_13693;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_78 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_78 <= _GEN_13694;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_79 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_79 <= _GEN_13695;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_80 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_80 <= _GEN_13696;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_81 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_81 <= _GEN_13697;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_82 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_82 <= _GEN_13698;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_83 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_83 <= _GEN_13699;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_84 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_84 <= _GEN_13700;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_85 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_85 <= _GEN_13701;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_86 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_86 <= _GEN_13702;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_87 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_87 <= _GEN_13703;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_88 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_88 <= _GEN_13704;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_89 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_89 <= _GEN_13705;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_90 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_90 <= _GEN_13706;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_91 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_91 <= _GEN_13707;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_92 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_92 <= _GEN_13708;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_93 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_93 <= _GEN_13709;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_94 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_94 <= _GEN_13710;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_95 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_95 <= _GEN_13711;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_96 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_96 <= _GEN_13712;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_97 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_97 <= _GEN_13713;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_98 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_98 <= _GEN_13714;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_99 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_99 <= _GEN_13715;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_100 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_100 <= _GEN_13716;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_101 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_101 <= _GEN_13717;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_102 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_102 <= _GEN_13718;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_103 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_103 <= _GEN_13719;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_104 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_104 <= _GEN_13720;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_105 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_105 <= _GEN_13721;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_106 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_106 <= _GEN_13722;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_107 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_107 <= _GEN_13723;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_108 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_108 <= _GEN_13724;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_109 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_109 <= _GEN_13725;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_110 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_110 <= _GEN_13726;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_111 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_111 <= _GEN_13727;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_112 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_112 <= _GEN_13728;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_113 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_113 <= _GEN_13729;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_114 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_114 <= _GEN_13730;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_115 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_115 <= _GEN_13731;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_116 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_116 <= _GEN_13732;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_117 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_117 <= _GEN_13733;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_118 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_118 <= _GEN_13734;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_119 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_119 <= _GEN_13735;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_120 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_120 <= _GEN_13736;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_121 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_121 <= _GEN_13737;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_122 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_122 <= _GEN_13738;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_123 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_123 <= _GEN_13739;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_124 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_124 <= _GEN_13740;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_125 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_125 <= _GEN_13741;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_126 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_126 <= _GEN_13742;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_1_127 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_127 <= _GEN_13743;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_0 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_0 <= _GEN_3211;
        end else begin
          dirty_0_0 <= _GEN_13746;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_1 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_1 <= _GEN_3212;
        end else begin
          dirty_0_1 <= _GEN_13747;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_2 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_2 <= _GEN_3213;
        end else begin
          dirty_0_2 <= _GEN_13748;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_3 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_3 <= _GEN_3214;
        end else begin
          dirty_0_3 <= _GEN_13749;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_4 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_4 <= _GEN_3215;
        end else begin
          dirty_0_4 <= _GEN_13750;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_5 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_5 <= _GEN_3216;
        end else begin
          dirty_0_5 <= _GEN_13751;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_6 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_6 <= _GEN_3217;
        end else begin
          dirty_0_6 <= _GEN_13752;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_7 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_7 <= _GEN_3218;
        end else begin
          dirty_0_7 <= _GEN_13753;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_8 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_8 <= _GEN_3219;
        end else begin
          dirty_0_8 <= _GEN_13754;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_9 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_9 <= _GEN_3220;
        end else begin
          dirty_0_9 <= _GEN_13755;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_10 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_10 <= _GEN_3221;
        end else begin
          dirty_0_10 <= _GEN_13756;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_11 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_11 <= _GEN_3222;
        end else begin
          dirty_0_11 <= _GEN_13757;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_12 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_12 <= _GEN_3223;
        end else begin
          dirty_0_12 <= _GEN_13758;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_13 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_13 <= _GEN_3224;
        end else begin
          dirty_0_13 <= _GEN_13759;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_14 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_14 <= _GEN_3225;
        end else begin
          dirty_0_14 <= _GEN_13760;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_15 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_15 <= _GEN_3226;
        end else begin
          dirty_0_15 <= _GEN_13761;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_16 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_16 <= _GEN_3227;
        end else begin
          dirty_0_16 <= _GEN_13762;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_17 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_17 <= _GEN_3228;
        end else begin
          dirty_0_17 <= _GEN_13763;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_18 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_18 <= _GEN_3229;
        end else begin
          dirty_0_18 <= _GEN_13764;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_19 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_19 <= _GEN_3230;
        end else begin
          dirty_0_19 <= _GEN_13765;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_20 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_20 <= _GEN_3231;
        end else begin
          dirty_0_20 <= _GEN_13766;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_21 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_21 <= _GEN_3232;
        end else begin
          dirty_0_21 <= _GEN_13767;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_22 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_22 <= _GEN_3233;
        end else begin
          dirty_0_22 <= _GEN_13768;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_23 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_23 <= _GEN_3234;
        end else begin
          dirty_0_23 <= _GEN_13769;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_24 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_24 <= _GEN_3235;
        end else begin
          dirty_0_24 <= _GEN_13770;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_25 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_25 <= _GEN_3236;
        end else begin
          dirty_0_25 <= _GEN_13771;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_26 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_26 <= _GEN_3237;
        end else begin
          dirty_0_26 <= _GEN_13772;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_27 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_27 <= _GEN_3238;
        end else begin
          dirty_0_27 <= _GEN_13773;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_28 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_28 <= _GEN_3239;
        end else begin
          dirty_0_28 <= _GEN_13774;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_29 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_29 <= _GEN_3240;
        end else begin
          dirty_0_29 <= _GEN_13775;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_30 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_30 <= _GEN_3241;
        end else begin
          dirty_0_30 <= _GEN_13776;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_31 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_31 <= _GEN_3242;
        end else begin
          dirty_0_31 <= _GEN_13777;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_32 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_32 <= _GEN_3243;
        end else begin
          dirty_0_32 <= _GEN_13778;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_33 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_33 <= _GEN_3244;
        end else begin
          dirty_0_33 <= _GEN_13779;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_34 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_34 <= _GEN_3245;
        end else begin
          dirty_0_34 <= _GEN_13780;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_35 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_35 <= _GEN_3246;
        end else begin
          dirty_0_35 <= _GEN_13781;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_36 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_36 <= _GEN_3247;
        end else begin
          dirty_0_36 <= _GEN_13782;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_37 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_37 <= _GEN_3248;
        end else begin
          dirty_0_37 <= _GEN_13783;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_38 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_38 <= _GEN_3249;
        end else begin
          dirty_0_38 <= _GEN_13784;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_39 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_39 <= _GEN_3250;
        end else begin
          dirty_0_39 <= _GEN_13785;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_40 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_40 <= _GEN_3251;
        end else begin
          dirty_0_40 <= _GEN_13786;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_41 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_41 <= _GEN_3252;
        end else begin
          dirty_0_41 <= _GEN_13787;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_42 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_42 <= _GEN_3253;
        end else begin
          dirty_0_42 <= _GEN_13788;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_43 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_43 <= _GEN_3254;
        end else begin
          dirty_0_43 <= _GEN_13789;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_44 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_44 <= _GEN_3255;
        end else begin
          dirty_0_44 <= _GEN_13790;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_45 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_45 <= _GEN_3256;
        end else begin
          dirty_0_45 <= _GEN_13791;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_46 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_46 <= _GEN_3257;
        end else begin
          dirty_0_46 <= _GEN_13792;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_47 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_47 <= _GEN_3258;
        end else begin
          dirty_0_47 <= _GEN_13793;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_48 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_48 <= _GEN_3259;
        end else begin
          dirty_0_48 <= _GEN_13794;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_49 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_49 <= _GEN_3260;
        end else begin
          dirty_0_49 <= _GEN_13795;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_50 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_50 <= _GEN_3261;
        end else begin
          dirty_0_50 <= _GEN_13796;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_51 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_51 <= _GEN_3262;
        end else begin
          dirty_0_51 <= _GEN_13797;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_52 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_52 <= _GEN_3263;
        end else begin
          dirty_0_52 <= _GEN_13798;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_53 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_53 <= _GEN_3264;
        end else begin
          dirty_0_53 <= _GEN_13799;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_54 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_54 <= _GEN_3265;
        end else begin
          dirty_0_54 <= _GEN_13800;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_55 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_55 <= _GEN_3266;
        end else begin
          dirty_0_55 <= _GEN_13801;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_56 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_56 <= _GEN_3267;
        end else begin
          dirty_0_56 <= _GEN_13802;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_57 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_57 <= _GEN_3268;
        end else begin
          dirty_0_57 <= _GEN_13803;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_58 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_58 <= _GEN_3269;
        end else begin
          dirty_0_58 <= _GEN_13804;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_59 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_59 <= _GEN_3270;
        end else begin
          dirty_0_59 <= _GEN_13805;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_60 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_60 <= _GEN_3271;
        end else begin
          dirty_0_60 <= _GEN_13806;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_61 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_61 <= _GEN_3272;
        end else begin
          dirty_0_61 <= _GEN_13807;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_62 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_62 <= _GEN_3273;
        end else begin
          dirty_0_62 <= _GEN_13808;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_63 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_63 <= _GEN_3274;
        end else begin
          dirty_0_63 <= _GEN_13809;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_64 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_64 <= _GEN_3275;
        end else begin
          dirty_0_64 <= _GEN_13810;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_65 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_65 <= _GEN_3276;
        end else begin
          dirty_0_65 <= _GEN_13811;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_66 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_66 <= _GEN_3277;
        end else begin
          dirty_0_66 <= _GEN_13812;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_67 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_67 <= _GEN_3278;
        end else begin
          dirty_0_67 <= _GEN_13813;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_68 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_68 <= _GEN_3279;
        end else begin
          dirty_0_68 <= _GEN_13814;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_69 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_69 <= _GEN_3280;
        end else begin
          dirty_0_69 <= _GEN_13815;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_70 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_70 <= _GEN_3281;
        end else begin
          dirty_0_70 <= _GEN_13816;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_71 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_71 <= _GEN_3282;
        end else begin
          dirty_0_71 <= _GEN_13817;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_72 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_72 <= _GEN_3283;
        end else begin
          dirty_0_72 <= _GEN_13818;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_73 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_73 <= _GEN_3284;
        end else begin
          dirty_0_73 <= _GEN_13819;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_74 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_74 <= _GEN_3285;
        end else begin
          dirty_0_74 <= _GEN_13820;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_75 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_75 <= _GEN_3286;
        end else begin
          dirty_0_75 <= _GEN_13821;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_76 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_76 <= _GEN_3287;
        end else begin
          dirty_0_76 <= _GEN_13822;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_77 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_77 <= _GEN_3288;
        end else begin
          dirty_0_77 <= _GEN_13823;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_78 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_78 <= _GEN_3289;
        end else begin
          dirty_0_78 <= _GEN_13824;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_79 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_79 <= _GEN_3290;
        end else begin
          dirty_0_79 <= _GEN_13825;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_80 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_80 <= _GEN_3291;
        end else begin
          dirty_0_80 <= _GEN_13826;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_81 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_81 <= _GEN_3292;
        end else begin
          dirty_0_81 <= _GEN_13827;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_82 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_82 <= _GEN_3293;
        end else begin
          dirty_0_82 <= _GEN_13828;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_83 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_83 <= _GEN_3294;
        end else begin
          dirty_0_83 <= _GEN_13829;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_84 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_84 <= _GEN_3295;
        end else begin
          dirty_0_84 <= _GEN_13830;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_85 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_85 <= _GEN_3296;
        end else begin
          dirty_0_85 <= _GEN_13831;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_86 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_86 <= _GEN_3297;
        end else begin
          dirty_0_86 <= _GEN_13832;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_87 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_87 <= _GEN_3298;
        end else begin
          dirty_0_87 <= _GEN_13833;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_88 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_88 <= _GEN_3299;
        end else begin
          dirty_0_88 <= _GEN_13834;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_89 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_89 <= _GEN_3300;
        end else begin
          dirty_0_89 <= _GEN_13835;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_90 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_90 <= _GEN_3301;
        end else begin
          dirty_0_90 <= _GEN_13836;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_91 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_91 <= _GEN_3302;
        end else begin
          dirty_0_91 <= _GEN_13837;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_92 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_92 <= _GEN_3303;
        end else begin
          dirty_0_92 <= _GEN_13838;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_93 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_93 <= _GEN_3304;
        end else begin
          dirty_0_93 <= _GEN_13839;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_94 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_94 <= _GEN_3305;
        end else begin
          dirty_0_94 <= _GEN_13840;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_95 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_95 <= _GEN_3306;
        end else begin
          dirty_0_95 <= _GEN_13841;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_96 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_96 <= _GEN_3307;
        end else begin
          dirty_0_96 <= _GEN_13842;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_97 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_97 <= _GEN_3308;
        end else begin
          dirty_0_97 <= _GEN_13843;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_98 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_98 <= _GEN_3309;
        end else begin
          dirty_0_98 <= _GEN_13844;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_99 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_99 <= _GEN_3310;
        end else begin
          dirty_0_99 <= _GEN_13845;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_100 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_100 <= _GEN_3311;
        end else begin
          dirty_0_100 <= _GEN_13846;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_101 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_101 <= _GEN_3312;
        end else begin
          dirty_0_101 <= _GEN_13847;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_102 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_102 <= _GEN_3313;
        end else begin
          dirty_0_102 <= _GEN_13848;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_103 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_103 <= _GEN_3314;
        end else begin
          dirty_0_103 <= _GEN_13849;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_104 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_104 <= _GEN_3315;
        end else begin
          dirty_0_104 <= _GEN_13850;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_105 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_105 <= _GEN_3316;
        end else begin
          dirty_0_105 <= _GEN_13851;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_106 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_106 <= _GEN_3317;
        end else begin
          dirty_0_106 <= _GEN_13852;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_107 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_107 <= _GEN_3318;
        end else begin
          dirty_0_107 <= _GEN_13853;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_108 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_108 <= _GEN_3319;
        end else begin
          dirty_0_108 <= _GEN_13854;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_109 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_109 <= _GEN_3320;
        end else begin
          dirty_0_109 <= _GEN_13855;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_110 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_110 <= _GEN_3321;
        end else begin
          dirty_0_110 <= _GEN_13856;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_111 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_111 <= _GEN_3322;
        end else begin
          dirty_0_111 <= _GEN_13857;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_112 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_112 <= _GEN_3323;
        end else begin
          dirty_0_112 <= _GEN_13858;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_113 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_113 <= _GEN_3324;
        end else begin
          dirty_0_113 <= _GEN_13859;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_114 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_114 <= _GEN_3325;
        end else begin
          dirty_0_114 <= _GEN_13860;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_115 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_115 <= _GEN_3326;
        end else begin
          dirty_0_115 <= _GEN_13861;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_116 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_116 <= _GEN_3327;
        end else begin
          dirty_0_116 <= _GEN_13862;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_117 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_117 <= _GEN_3328;
        end else begin
          dirty_0_117 <= _GEN_13863;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_118 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_118 <= _GEN_3329;
        end else begin
          dirty_0_118 <= _GEN_13864;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_119 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_119 <= _GEN_3330;
        end else begin
          dirty_0_119 <= _GEN_13865;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_120 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_120 <= _GEN_3331;
        end else begin
          dirty_0_120 <= _GEN_13866;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_121 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_121 <= _GEN_3332;
        end else begin
          dirty_0_121 <= _GEN_13867;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_122 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_122 <= _GEN_3333;
        end else begin
          dirty_0_122 <= _GEN_13868;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_123 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_123 <= _GEN_3334;
        end else begin
          dirty_0_123 <= _GEN_13869;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_124 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_124 <= _GEN_3335;
        end else begin
          dirty_0_124 <= _GEN_13870;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_125 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_125 <= _GEN_3336;
        end else begin
          dirty_0_125 <= _GEN_13871;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_126 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_126 <= _GEN_3337;
        end else begin
          dirty_0_126 <= _GEN_13872;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      dirty_0_127 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_127 <= _GEN_3338;
        end else begin
          dirty_0_127 <= _GEN_13873;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_0 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_0 <= _GEN_4107;
        end else begin
          dirty_1_0 <= _GEN_13874;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_1 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_1 <= _GEN_4108;
        end else begin
          dirty_1_1 <= _GEN_13875;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_2 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_2 <= _GEN_4109;
        end else begin
          dirty_1_2 <= _GEN_13876;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_3 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_3 <= _GEN_4110;
        end else begin
          dirty_1_3 <= _GEN_13877;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_4 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_4 <= _GEN_4111;
        end else begin
          dirty_1_4 <= _GEN_13878;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_5 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_5 <= _GEN_4112;
        end else begin
          dirty_1_5 <= _GEN_13879;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_6 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_6 <= _GEN_4113;
        end else begin
          dirty_1_6 <= _GEN_13880;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_7 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_7 <= _GEN_4114;
        end else begin
          dirty_1_7 <= _GEN_13881;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_8 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_8 <= _GEN_4115;
        end else begin
          dirty_1_8 <= _GEN_13882;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_9 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_9 <= _GEN_4116;
        end else begin
          dirty_1_9 <= _GEN_13883;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_10 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_10 <= _GEN_4117;
        end else begin
          dirty_1_10 <= _GEN_13884;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_11 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_11 <= _GEN_4118;
        end else begin
          dirty_1_11 <= _GEN_13885;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_12 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_12 <= _GEN_4119;
        end else begin
          dirty_1_12 <= _GEN_13886;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_13 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_13 <= _GEN_4120;
        end else begin
          dirty_1_13 <= _GEN_13887;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_14 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_14 <= _GEN_4121;
        end else begin
          dirty_1_14 <= _GEN_13888;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_15 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_15 <= _GEN_4122;
        end else begin
          dirty_1_15 <= _GEN_13889;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_16 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_16 <= _GEN_4123;
        end else begin
          dirty_1_16 <= _GEN_13890;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_17 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_17 <= _GEN_4124;
        end else begin
          dirty_1_17 <= _GEN_13891;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_18 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_18 <= _GEN_4125;
        end else begin
          dirty_1_18 <= _GEN_13892;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_19 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_19 <= _GEN_4126;
        end else begin
          dirty_1_19 <= _GEN_13893;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_20 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_20 <= _GEN_4127;
        end else begin
          dirty_1_20 <= _GEN_13894;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_21 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_21 <= _GEN_4128;
        end else begin
          dirty_1_21 <= _GEN_13895;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_22 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_22 <= _GEN_4129;
        end else begin
          dirty_1_22 <= _GEN_13896;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_23 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_23 <= _GEN_4130;
        end else begin
          dirty_1_23 <= _GEN_13897;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_24 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_24 <= _GEN_4131;
        end else begin
          dirty_1_24 <= _GEN_13898;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_25 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_25 <= _GEN_4132;
        end else begin
          dirty_1_25 <= _GEN_13899;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_26 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_26 <= _GEN_4133;
        end else begin
          dirty_1_26 <= _GEN_13900;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_27 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_27 <= _GEN_4134;
        end else begin
          dirty_1_27 <= _GEN_13901;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_28 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_28 <= _GEN_4135;
        end else begin
          dirty_1_28 <= _GEN_13902;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_29 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_29 <= _GEN_4136;
        end else begin
          dirty_1_29 <= _GEN_13903;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_30 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_30 <= _GEN_4137;
        end else begin
          dirty_1_30 <= _GEN_13904;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_31 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_31 <= _GEN_4138;
        end else begin
          dirty_1_31 <= _GEN_13905;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_32 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_32 <= _GEN_4139;
        end else begin
          dirty_1_32 <= _GEN_13906;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_33 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_33 <= _GEN_4140;
        end else begin
          dirty_1_33 <= _GEN_13907;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_34 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_34 <= _GEN_4141;
        end else begin
          dirty_1_34 <= _GEN_13908;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_35 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_35 <= _GEN_4142;
        end else begin
          dirty_1_35 <= _GEN_13909;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_36 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_36 <= _GEN_4143;
        end else begin
          dirty_1_36 <= _GEN_13910;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_37 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_37 <= _GEN_4144;
        end else begin
          dirty_1_37 <= _GEN_13911;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_38 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_38 <= _GEN_4145;
        end else begin
          dirty_1_38 <= _GEN_13912;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_39 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_39 <= _GEN_4146;
        end else begin
          dirty_1_39 <= _GEN_13913;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_40 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_40 <= _GEN_4147;
        end else begin
          dirty_1_40 <= _GEN_13914;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_41 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_41 <= _GEN_4148;
        end else begin
          dirty_1_41 <= _GEN_13915;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_42 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_42 <= _GEN_4149;
        end else begin
          dirty_1_42 <= _GEN_13916;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_43 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_43 <= _GEN_4150;
        end else begin
          dirty_1_43 <= _GEN_13917;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_44 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_44 <= _GEN_4151;
        end else begin
          dirty_1_44 <= _GEN_13918;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_45 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_45 <= _GEN_4152;
        end else begin
          dirty_1_45 <= _GEN_13919;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_46 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_46 <= _GEN_4153;
        end else begin
          dirty_1_46 <= _GEN_13920;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_47 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_47 <= _GEN_4154;
        end else begin
          dirty_1_47 <= _GEN_13921;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_48 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_48 <= _GEN_4155;
        end else begin
          dirty_1_48 <= _GEN_13922;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_49 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_49 <= _GEN_4156;
        end else begin
          dirty_1_49 <= _GEN_13923;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_50 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_50 <= _GEN_4157;
        end else begin
          dirty_1_50 <= _GEN_13924;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_51 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_51 <= _GEN_4158;
        end else begin
          dirty_1_51 <= _GEN_13925;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_52 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_52 <= _GEN_4159;
        end else begin
          dirty_1_52 <= _GEN_13926;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_53 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_53 <= _GEN_4160;
        end else begin
          dirty_1_53 <= _GEN_13927;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_54 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_54 <= _GEN_4161;
        end else begin
          dirty_1_54 <= _GEN_13928;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_55 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_55 <= _GEN_4162;
        end else begin
          dirty_1_55 <= _GEN_13929;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_56 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_56 <= _GEN_4163;
        end else begin
          dirty_1_56 <= _GEN_13930;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_57 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_57 <= _GEN_4164;
        end else begin
          dirty_1_57 <= _GEN_13931;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_58 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_58 <= _GEN_4165;
        end else begin
          dirty_1_58 <= _GEN_13932;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_59 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_59 <= _GEN_4166;
        end else begin
          dirty_1_59 <= _GEN_13933;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_60 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_60 <= _GEN_4167;
        end else begin
          dirty_1_60 <= _GEN_13934;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_61 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_61 <= _GEN_4168;
        end else begin
          dirty_1_61 <= _GEN_13935;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_62 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_62 <= _GEN_4169;
        end else begin
          dirty_1_62 <= _GEN_13936;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_63 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_63 <= _GEN_4170;
        end else begin
          dirty_1_63 <= _GEN_13937;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_64 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_64 <= _GEN_4171;
        end else begin
          dirty_1_64 <= _GEN_13938;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_65 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_65 <= _GEN_4172;
        end else begin
          dirty_1_65 <= _GEN_13939;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_66 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_66 <= _GEN_4173;
        end else begin
          dirty_1_66 <= _GEN_13940;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_67 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_67 <= _GEN_4174;
        end else begin
          dirty_1_67 <= _GEN_13941;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_68 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_68 <= _GEN_4175;
        end else begin
          dirty_1_68 <= _GEN_13942;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_69 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_69 <= _GEN_4176;
        end else begin
          dirty_1_69 <= _GEN_13943;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_70 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_70 <= _GEN_4177;
        end else begin
          dirty_1_70 <= _GEN_13944;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_71 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_71 <= _GEN_4178;
        end else begin
          dirty_1_71 <= _GEN_13945;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_72 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_72 <= _GEN_4179;
        end else begin
          dirty_1_72 <= _GEN_13946;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_73 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_73 <= _GEN_4180;
        end else begin
          dirty_1_73 <= _GEN_13947;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_74 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_74 <= _GEN_4181;
        end else begin
          dirty_1_74 <= _GEN_13948;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_75 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_75 <= _GEN_4182;
        end else begin
          dirty_1_75 <= _GEN_13949;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_76 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_76 <= _GEN_4183;
        end else begin
          dirty_1_76 <= _GEN_13950;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_77 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_77 <= _GEN_4184;
        end else begin
          dirty_1_77 <= _GEN_13951;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_78 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_78 <= _GEN_4185;
        end else begin
          dirty_1_78 <= _GEN_13952;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_79 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_79 <= _GEN_4186;
        end else begin
          dirty_1_79 <= _GEN_13953;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_80 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_80 <= _GEN_4187;
        end else begin
          dirty_1_80 <= _GEN_13954;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_81 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_81 <= _GEN_4188;
        end else begin
          dirty_1_81 <= _GEN_13955;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_82 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_82 <= _GEN_4189;
        end else begin
          dirty_1_82 <= _GEN_13956;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_83 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_83 <= _GEN_4190;
        end else begin
          dirty_1_83 <= _GEN_13957;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_84 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_84 <= _GEN_4191;
        end else begin
          dirty_1_84 <= _GEN_13958;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_85 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_85 <= _GEN_4192;
        end else begin
          dirty_1_85 <= _GEN_13959;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_86 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_86 <= _GEN_4193;
        end else begin
          dirty_1_86 <= _GEN_13960;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_87 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_87 <= _GEN_4194;
        end else begin
          dirty_1_87 <= _GEN_13961;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_88 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_88 <= _GEN_4195;
        end else begin
          dirty_1_88 <= _GEN_13962;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_89 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_89 <= _GEN_4196;
        end else begin
          dirty_1_89 <= _GEN_13963;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_90 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_90 <= _GEN_4197;
        end else begin
          dirty_1_90 <= _GEN_13964;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_91 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_91 <= _GEN_4198;
        end else begin
          dirty_1_91 <= _GEN_13965;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_92 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_92 <= _GEN_4199;
        end else begin
          dirty_1_92 <= _GEN_13966;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_93 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_93 <= _GEN_4200;
        end else begin
          dirty_1_93 <= _GEN_13967;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_94 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_94 <= _GEN_4201;
        end else begin
          dirty_1_94 <= _GEN_13968;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_95 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_95 <= _GEN_4202;
        end else begin
          dirty_1_95 <= _GEN_13969;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_96 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_96 <= _GEN_4203;
        end else begin
          dirty_1_96 <= _GEN_13970;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_97 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_97 <= _GEN_4204;
        end else begin
          dirty_1_97 <= _GEN_13971;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_98 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_98 <= _GEN_4205;
        end else begin
          dirty_1_98 <= _GEN_13972;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_99 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_99 <= _GEN_4206;
        end else begin
          dirty_1_99 <= _GEN_13973;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_100 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_100 <= _GEN_4207;
        end else begin
          dirty_1_100 <= _GEN_13974;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_101 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_101 <= _GEN_4208;
        end else begin
          dirty_1_101 <= _GEN_13975;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_102 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_102 <= _GEN_4209;
        end else begin
          dirty_1_102 <= _GEN_13976;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_103 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_103 <= _GEN_4210;
        end else begin
          dirty_1_103 <= _GEN_13977;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_104 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_104 <= _GEN_4211;
        end else begin
          dirty_1_104 <= _GEN_13978;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_105 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_105 <= _GEN_4212;
        end else begin
          dirty_1_105 <= _GEN_13979;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_106 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_106 <= _GEN_4213;
        end else begin
          dirty_1_106 <= _GEN_13980;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_107 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_107 <= _GEN_4214;
        end else begin
          dirty_1_107 <= _GEN_13981;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_108 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_108 <= _GEN_4215;
        end else begin
          dirty_1_108 <= _GEN_13982;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_109 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_109 <= _GEN_4216;
        end else begin
          dirty_1_109 <= _GEN_13983;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_110 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_110 <= _GEN_4217;
        end else begin
          dirty_1_110 <= _GEN_13984;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_111 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_111 <= _GEN_4218;
        end else begin
          dirty_1_111 <= _GEN_13985;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_112 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_112 <= _GEN_4219;
        end else begin
          dirty_1_112 <= _GEN_13986;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_113 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_113 <= _GEN_4220;
        end else begin
          dirty_1_113 <= _GEN_13987;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_114 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_114 <= _GEN_4221;
        end else begin
          dirty_1_114 <= _GEN_13988;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_115 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_115 <= _GEN_4222;
        end else begin
          dirty_1_115 <= _GEN_13989;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_116 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_116 <= _GEN_4223;
        end else begin
          dirty_1_116 <= _GEN_13990;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_117 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_117 <= _GEN_4224;
        end else begin
          dirty_1_117 <= _GEN_13991;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_118 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_118 <= _GEN_4225;
        end else begin
          dirty_1_118 <= _GEN_13992;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_119 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_119 <= _GEN_4226;
        end else begin
          dirty_1_119 <= _GEN_13993;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_120 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_120 <= _GEN_4227;
        end else begin
          dirty_1_120 <= _GEN_13994;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_121 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_121 <= _GEN_4228;
        end else begin
          dirty_1_121 <= _GEN_13995;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_122 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_122 <= _GEN_4229;
        end else begin
          dirty_1_122 <= _GEN_13996;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_123 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_123 <= _GEN_4230;
        end else begin
          dirty_1_123 <= _GEN_13997;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_124 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_124 <= _GEN_4231;
        end else begin
          dirty_1_124 <= _GEN_13998;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_125 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_125 <= _GEN_4232;
        end else begin
          dirty_1_125 <= _GEN_13999;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_126 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_126 <= _GEN_4233;
        end else begin
          dirty_1_126 <= _GEN_14000;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 33:26]
      dirty_1_127 <= 1'h0; // @[d_cache.scala 33:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (3'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_127 <= _GEN_4234;
        end else begin
          dirty_1_127 <= _GEN_14001;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:27]
      way0_hit <= 1'h0; // @[d_cache.scala 34:27]
    end else begin
      way0_hit <= _T_4;
    end
    if (reset) begin // @[d_cache.scala 35:27]
      way1_hit <= 1'h0; // @[d_cache.scala 35:27]
    end else begin
      way1_hit <= _T_7;
    end
    if (reset) begin // @[d_cache.scala 37:34]
      write_back_data <= 64'h0; // @[d_cache.scala 37:34]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          write_back_data <= _GEN_13744;
        end
      end
    end
    write_back_addr <= _GEN_20774[31:0]; // @[d_cache.scala 38:{34,34}]
    if (reset) begin // @[d_cache.scala 41:28]
      unuse_way <= 2'h0; // @[d_cache.scala 41:28]
    end else if (~_GEN_255) begin // @[d_cache.scala 74:31]
      unuse_way <= 2'h1; // @[d_cache.scala 75:19]
    end else if (~_GEN_512) begin // @[d_cache.scala 76:37]
      unuse_way <= 2'h2; // @[d_cache.scala 77:19]
    end else begin
      unuse_way <= 2'h0; // @[d_cache.scala 79:19]
    end
    if (reset) begin // @[d_cache.scala 42:31]
      receive_data <= 64'h0; // @[d_cache.scala 42:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          receive_data <= _GEN_12974;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 43:24]
      quene <= 1'h0; // @[d_cache.scala 43:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 87:18]
          quene <= _GEN_13359;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 82:24]
      state <= 3'h0; // @[d_cache.scala 82:24]
    end else if (3'h0 == state) begin // @[d_cache.scala 87:18]
      if (io_from_lsu_arvalid) begin // @[d_cache.scala 89:38]
        state <= 3'h1; // @[d_cache.scala 90:23]
      end else if (io_from_lsu_awvalid) begin // @[d_cache.scala 91:44]
        state <= 3'h2; // @[d_cache.scala 92:23]
      end
    end else if (3'h1 == state) begin // @[d_cache.scala 87:18]
      if (way0_hit) begin // @[d_cache.scala 97:27]
        state <= _GEN_646;
      end else begin
        state <= _GEN_775;
      end
    end else if (3'h2 == state) begin // @[d_cache.scala 87:18]
      state <= _GEN_3082;
    end else begin
      state <= _GEN_12973;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"read addr : %x  write addr : %x\n",io_from_lsu_araddr,io_from_lsu_awaddr); // @[d_cache.scala 16:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"d_cache state:%d\n",state); // @[d_cache.scala 83:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"receive data:%x\n",receive_data); // @[d_cache.scala 85:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_14 & _T_15 & way0_hit & io_from_lsu_rready & _T_1) begin
          $fwrite(32'h80000002,"dirty_0:%d\n",7'h7f == index ? dirty_0_127 : _GEN_644); // @[d_cache.scala 99:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_20776 & ~way0_hit & way1_hit & io_from_lsu_rready & _T_1) begin
          $fwrite(32'h80000002,"dirty_1:%d\n",7'h7f == index ? dirty_1_127 : _GEN_773); // @[d_cache.scala 105:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"cacheline0:%x   cacheline1:%x\n",_GEN_904,_GEN_1416); // @[d_cache.scala 373:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"record_wdata1:%x  record_wstrb1:%x record_pc:%x record_awaddr:%x record_olddata:%x\n",7'h7f
             == index ? record_wdata1_127 : _GEN_19231,7'h7f == index ? record_wstrb1_127 : _GEN_19359,7'h7f == index ?
            record_pc_127 : _GEN_19487,7'h7f == index ? record_addr_127 : _GEN_19615,7'h7f == index ? record_olddata_127
             : _GEN_19743); // @[d_cache.scala 374:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ram_0_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ram_0_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ram_0_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ram_0_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ram_0_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ram_0_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ram_0_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ram_0_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  ram_0_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  ram_0_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  ram_0_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  ram_0_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  ram_0_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  ram_0_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  ram_0_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  ram_0_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  ram_0_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  ram_0_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  ram_0_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  ram_0_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  ram_0_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  ram_0_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  ram_0_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  ram_0_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  ram_0_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  ram_0_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  ram_0_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  ram_0_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  ram_0_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  ram_0_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  ram_0_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  ram_0_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  ram_0_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  ram_0_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  ram_0_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  ram_0_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  ram_0_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  ram_0_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  ram_0_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  ram_0_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  ram_0_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  ram_0_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  ram_0_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  ram_0_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  ram_0_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  ram_0_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  ram_0_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  ram_0_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  ram_0_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  ram_0_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  ram_0_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  ram_0_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  ram_0_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  ram_0_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  ram_0_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  ram_0_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  ram_0_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  ram_0_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  ram_0_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  ram_0_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  ram_0_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  ram_0_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  ram_0_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  ram_0_63 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  ram_0_64 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  ram_0_65 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  ram_0_66 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  ram_0_67 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  ram_0_68 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  ram_0_69 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  ram_0_70 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  ram_0_71 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  ram_0_72 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  ram_0_73 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  ram_0_74 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  ram_0_75 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  ram_0_76 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  ram_0_77 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  ram_0_78 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  ram_0_79 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  ram_0_80 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  ram_0_81 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  ram_0_82 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  ram_0_83 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  ram_0_84 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  ram_0_85 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  ram_0_86 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  ram_0_87 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  ram_0_88 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  ram_0_89 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  ram_0_90 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  ram_0_91 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  ram_0_92 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  ram_0_93 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  ram_0_94 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  ram_0_95 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  ram_0_96 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  ram_0_97 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  ram_0_98 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  ram_0_99 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  ram_0_100 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  ram_0_101 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  ram_0_102 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  ram_0_103 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  ram_0_104 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  ram_0_105 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  ram_0_106 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  ram_0_107 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  ram_0_108 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  ram_0_109 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  ram_0_110 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  ram_0_111 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  ram_0_112 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  ram_0_113 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  ram_0_114 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  ram_0_115 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  ram_0_116 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  ram_0_117 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  ram_0_118 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  ram_0_119 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  ram_0_120 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  ram_0_121 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  ram_0_122 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  ram_0_123 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  ram_0_124 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  ram_0_125 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  ram_0_126 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  ram_0_127 = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  ram_1_0 = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  ram_1_1 = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  ram_1_2 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  ram_1_3 = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  ram_1_4 = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  ram_1_5 = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  ram_1_6 = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  ram_1_7 = _RAND_135[63:0];
  _RAND_136 = {2{`RANDOM}};
  ram_1_8 = _RAND_136[63:0];
  _RAND_137 = {2{`RANDOM}};
  ram_1_9 = _RAND_137[63:0];
  _RAND_138 = {2{`RANDOM}};
  ram_1_10 = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  ram_1_11 = _RAND_139[63:0];
  _RAND_140 = {2{`RANDOM}};
  ram_1_12 = _RAND_140[63:0];
  _RAND_141 = {2{`RANDOM}};
  ram_1_13 = _RAND_141[63:0];
  _RAND_142 = {2{`RANDOM}};
  ram_1_14 = _RAND_142[63:0];
  _RAND_143 = {2{`RANDOM}};
  ram_1_15 = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  ram_1_16 = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  ram_1_17 = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  ram_1_18 = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  ram_1_19 = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  ram_1_20 = _RAND_148[63:0];
  _RAND_149 = {2{`RANDOM}};
  ram_1_21 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  ram_1_22 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  ram_1_23 = _RAND_151[63:0];
  _RAND_152 = {2{`RANDOM}};
  ram_1_24 = _RAND_152[63:0];
  _RAND_153 = {2{`RANDOM}};
  ram_1_25 = _RAND_153[63:0];
  _RAND_154 = {2{`RANDOM}};
  ram_1_26 = _RAND_154[63:0];
  _RAND_155 = {2{`RANDOM}};
  ram_1_27 = _RAND_155[63:0];
  _RAND_156 = {2{`RANDOM}};
  ram_1_28 = _RAND_156[63:0];
  _RAND_157 = {2{`RANDOM}};
  ram_1_29 = _RAND_157[63:0];
  _RAND_158 = {2{`RANDOM}};
  ram_1_30 = _RAND_158[63:0];
  _RAND_159 = {2{`RANDOM}};
  ram_1_31 = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  ram_1_32 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  ram_1_33 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  ram_1_34 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  ram_1_35 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  ram_1_36 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  ram_1_37 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  ram_1_38 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  ram_1_39 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  ram_1_40 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  ram_1_41 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  ram_1_42 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  ram_1_43 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  ram_1_44 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  ram_1_45 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  ram_1_46 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  ram_1_47 = _RAND_175[63:0];
  _RAND_176 = {2{`RANDOM}};
  ram_1_48 = _RAND_176[63:0];
  _RAND_177 = {2{`RANDOM}};
  ram_1_49 = _RAND_177[63:0];
  _RAND_178 = {2{`RANDOM}};
  ram_1_50 = _RAND_178[63:0];
  _RAND_179 = {2{`RANDOM}};
  ram_1_51 = _RAND_179[63:0];
  _RAND_180 = {2{`RANDOM}};
  ram_1_52 = _RAND_180[63:0];
  _RAND_181 = {2{`RANDOM}};
  ram_1_53 = _RAND_181[63:0];
  _RAND_182 = {2{`RANDOM}};
  ram_1_54 = _RAND_182[63:0];
  _RAND_183 = {2{`RANDOM}};
  ram_1_55 = _RAND_183[63:0];
  _RAND_184 = {2{`RANDOM}};
  ram_1_56 = _RAND_184[63:0];
  _RAND_185 = {2{`RANDOM}};
  ram_1_57 = _RAND_185[63:0];
  _RAND_186 = {2{`RANDOM}};
  ram_1_58 = _RAND_186[63:0];
  _RAND_187 = {2{`RANDOM}};
  ram_1_59 = _RAND_187[63:0];
  _RAND_188 = {2{`RANDOM}};
  ram_1_60 = _RAND_188[63:0];
  _RAND_189 = {2{`RANDOM}};
  ram_1_61 = _RAND_189[63:0];
  _RAND_190 = {2{`RANDOM}};
  ram_1_62 = _RAND_190[63:0];
  _RAND_191 = {2{`RANDOM}};
  ram_1_63 = _RAND_191[63:0];
  _RAND_192 = {2{`RANDOM}};
  ram_1_64 = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  ram_1_65 = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  ram_1_66 = _RAND_194[63:0];
  _RAND_195 = {2{`RANDOM}};
  ram_1_67 = _RAND_195[63:0];
  _RAND_196 = {2{`RANDOM}};
  ram_1_68 = _RAND_196[63:0];
  _RAND_197 = {2{`RANDOM}};
  ram_1_69 = _RAND_197[63:0];
  _RAND_198 = {2{`RANDOM}};
  ram_1_70 = _RAND_198[63:0];
  _RAND_199 = {2{`RANDOM}};
  ram_1_71 = _RAND_199[63:0];
  _RAND_200 = {2{`RANDOM}};
  ram_1_72 = _RAND_200[63:0];
  _RAND_201 = {2{`RANDOM}};
  ram_1_73 = _RAND_201[63:0];
  _RAND_202 = {2{`RANDOM}};
  ram_1_74 = _RAND_202[63:0];
  _RAND_203 = {2{`RANDOM}};
  ram_1_75 = _RAND_203[63:0];
  _RAND_204 = {2{`RANDOM}};
  ram_1_76 = _RAND_204[63:0];
  _RAND_205 = {2{`RANDOM}};
  ram_1_77 = _RAND_205[63:0];
  _RAND_206 = {2{`RANDOM}};
  ram_1_78 = _RAND_206[63:0];
  _RAND_207 = {2{`RANDOM}};
  ram_1_79 = _RAND_207[63:0];
  _RAND_208 = {2{`RANDOM}};
  ram_1_80 = _RAND_208[63:0];
  _RAND_209 = {2{`RANDOM}};
  ram_1_81 = _RAND_209[63:0];
  _RAND_210 = {2{`RANDOM}};
  ram_1_82 = _RAND_210[63:0];
  _RAND_211 = {2{`RANDOM}};
  ram_1_83 = _RAND_211[63:0];
  _RAND_212 = {2{`RANDOM}};
  ram_1_84 = _RAND_212[63:0];
  _RAND_213 = {2{`RANDOM}};
  ram_1_85 = _RAND_213[63:0];
  _RAND_214 = {2{`RANDOM}};
  ram_1_86 = _RAND_214[63:0];
  _RAND_215 = {2{`RANDOM}};
  ram_1_87 = _RAND_215[63:0];
  _RAND_216 = {2{`RANDOM}};
  ram_1_88 = _RAND_216[63:0];
  _RAND_217 = {2{`RANDOM}};
  ram_1_89 = _RAND_217[63:0];
  _RAND_218 = {2{`RANDOM}};
  ram_1_90 = _RAND_218[63:0];
  _RAND_219 = {2{`RANDOM}};
  ram_1_91 = _RAND_219[63:0];
  _RAND_220 = {2{`RANDOM}};
  ram_1_92 = _RAND_220[63:0];
  _RAND_221 = {2{`RANDOM}};
  ram_1_93 = _RAND_221[63:0];
  _RAND_222 = {2{`RANDOM}};
  ram_1_94 = _RAND_222[63:0];
  _RAND_223 = {2{`RANDOM}};
  ram_1_95 = _RAND_223[63:0];
  _RAND_224 = {2{`RANDOM}};
  ram_1_96 = _RAND_224[63:0];
  _RAND_225 = {2{`RANDOM}};
  ram_1_97 = _RAND_225[63:0];
  _RAND_226 = {2{`RANDOM}};
  ram_1_98 = _RAND_226[63:0];
  _RAND_227 = {2{`RANDOM}};
  ram_1_99 = _RAND_227[63:0];
  _RAND_228 = {2{`RANDOM}};
  ram_1_100 = _RAND_228[63:0];
  _RAND_229 = {2{`RANDOM}};
  ram_1_101 = _RAND_229[63:0];
  _RAND_230 = {2{`RANDOM}};
  ram_1_102 = _RAND_230[63:0];
  _RAND_231 = {2{`RANDOM}};
  ram_1_103 = _RAND_231[63:0];
  _RAND_232 = {2{`RANDOM}};
  ram_1_104 = _RAND_232[63:0];
  _RAND_233 = {2{`RANDOM}};
  ram_1_105 = _RAND_233[63:0];
  _RAND_234 = {2{`RANDOM}};
  ram_1_106 = _RAND_234[63:0];
  _RAND_235 = {2{`RANDOM}};
  ram_1_107 = _RAND_235[63:0];
  _RAND_236 = {2{`RANDOM}};
  ram_1_108 = _RAND_236[63:0];
  _RAND_237 = {2{`RANDOM}};
  ram_1_109 = _RAND_237[63:0];
  _RAND_238 = {2{`RANDOM}};
  ram_1_110 = _RAND_238[63:0];
  _RAND_239 = {2{`RANDOM}};
  ram_1_111 = _RAND_239[63:0];
  _RAND_240 = {2{`RANDOM}};
  ram_1_112 = _RAND_240[63:0];
  _RAND_241 = {2{`RANDOM}};
  ram_1_113 = _RAND_241[63:0];
  _RAND_242 = {2{`RANDOM}};
  ram_1_114 = _RAND_242[63:0];
  _RAND_243 = {2{`RANDOM}};
  ram_1_115 = _RAND_243[63:0];
  _RAND_244 = {2{`RANDOM}};
  ram_1_116 = _RAND_244[63:0];
  _RAND_245 = {2{`RANDOM}};
  ram_1_117 = _RAND_245[63:0];
  _RAND_246 = {2{`RANDOM}};
  ram_1_118 = _RAND_246[63:0];
  _RAND_247 = {2{`RANDOM}};
  ram_1_119 = _RAND_247[63:0];
  _RAND_248 = {2{`RANDOM}};
  ram_1_120 = _RAND_248[63:0];
  _RAND_249 = {2{`RANDOM}};
  ram_1_121 = _RAND_249[63:0];
  _RAND_250 = {2{`RANDOM}};
  ram_1_122 = _RAND_250[63:0];
  _RAND_251 = {2{`RANDOM}};
  ram_1_123 = _RAND_251[63:0];
  _RAND_252 = {2{`RANDOM}};
  ram_1_124 = _RAND_252[63:0];
  _RAND_253 = {2{`RANDOM}};
  ram_1_125 = _RAND_253[63:0];
  _RAND_254 = {2{`RANDOM}};
  ram_1_126 = _RAND_254[63:0];
  _RAND_255 = {2{`RANDOM}};
  ram_1_127 = _RAND_255[63:0];
  _RAND_256 = {2{`RANDOM}};
  record_wdata1_0 = _RAND_256[63:0];
  _RAND_257 = {2{`RANDOM}};
  record_wdata1_1 = _RAND_257[63:0];
  _RAND_258 = {2{`RANDOM}};
  record_wdata1_2 = _RAND_258[63:0];
  _RAND_259 = {2{`RANDOM}};
  record_wdata1_3 = _RAND_259[63:0];
  _RAND_260 = {2{`RANDOM}};
  record_wdata1_4 = _RAND_260[63:0];
  _RAND_261 = {2{`RANDOM}};
  record_wdata1_5 = _RAND_261[63:0];
  _RAND_262 = {2{`RANDOM}};
  record_wdata1_6 = _RAND_262[63:0];
  _RAND_263 = {2{`RANDOM}};
  record_wdata1_7 = _RAND_263[63:0];
  _RAND_264 = {2{`RANDOM}};
  record_wdata1_8 = _RAND_264[63:0];
  _RAND_265 = {2{`RANDOM}};
  record_wdata1_9 = _RAND_265[63:0];
  _RAND_266 = {2{`RANDOM}};
  record_wdata1_10 = _RAND_266[63:0];
  _RAND_267 = {2{`RANDOM}};
  record_wdata1_11 = _RAND_267[63:0];
  _RAND_268 = {2{`RANDOM}};
  record_wdata1_12 = _RAND_268[63:0];
  _RAND_269 = {2{`RANDOM}};
  record_wdata1_13 = _RAND_269[63:0];
  _RAND_270 = {2{`RANDOM}};
  record_wdata1_14 = _RAND_270[63:0];
  _RAND_271 = {2{`RANDOM}};
  record_wdata1_15 = _RAND_271[63:0];
  _RAND_272 = {2{`RANDOM}};
  record_wdata1_16 = _RAND_272[63:0];
  _RAND_273 = {2{`RANDOM}};
  record_wdata1_17 = _RAND_273[63:0];
  _RAND_274 = {2{`RANDOM}};
  record_wdata1_18 = _RAND_274[63:0];
  _RAND_275 = {2{`RANDOM}};
  record_wdata1_19 = _RAND_275[63:0];
  _RAND_276 = {2{`RANDOM}};
  record_wdata1_20 = _RAND_276[63:0];
  _RAND_277 = {2{`RANDOM}};
  record_wdata1_21 = _RAND_277[63:0];
  _RAND_278 = {2{`RANDOM}};
  record_wdata1_22 = _RAND_278[63:0];
  _RAND_279 = {2{`RANDOM}};
  record_wdata1_23 = _RAND_279[63:0];
  _RAND_280 = {2{`RANDOM}};
  record_wdata1_24 = _RAND_280[63:0];
  _RAND_281 = {2{`RANDOM}};
  record_wdata1_25 = _RAND_281[63:0];
  _RAND_282 = {2{`RANDOM}};
  record_wdata1_26 = _RAND_282[63:0];
  _RAND_283 = {2{`RANDOM}};
  record_wdata1_27 = _RAND_283[63:0];
  _RAND_284 = {2{`RANDOM}};
  record_wdata1_28 = _RAND_284[63:0];
  _RAND_285 = {2{`RANDOM}};
  record_wdata1_29 = _RAND_285[63:0];
  _RAND_286 = {2{`RANDOM}};
  record_wdata1_30 = _RAND_286[63:0];
  _RAND_287 = {2{`RANDOM}};
  record_wdata1_31 = _RAND_287[63:0];
  _RAND_288 = {2{`RANDOM}};
  record_wdata1_32 = _RAND_288[63:0];
  _RAND_289 = {2{`RANDOM}};
  record_wdata1_33 = _RAND_289[63:0];
  _RAND_290 = {2{`RANDOM}};
  record_wdata1_34 = _RAND_290[63:0];
  _RAND_291 = {2{`RANDOM}};
  record_wdata1_35 = _RAND_291[63:0];
  _RAND_292 = {2{`RANDOM}};
  record_wdata1_36 = _RAND_292[63:0];
  _RAND_293 = {2{`RANDOM}};
  record_wdata1_37 = _RAND_293[63:0];
  _RAND_294 = {2{`RANDOM}};
  record_wdata1_38 = _RAND_294[63:0];
  _RAND_295 = {2{`RANDOM}};
  record_wdata1_39 = _RAND_295[63:0];
  _RAND_296 = {2{`RANDOM}};
  record_wdata1_40 = _RAND_296[63:0];
  _RAND_297 = {2{`RANDOM}};
  record_wdata1_41 = _RAND_297[63:0];
  _RAND_298 = {2{`RANDOM}};
  record_wdata1_42 = _RAND_298[63:0];
  _RAND_299 = {2{`RANDOM}};
  record_wdata1_43 = _RAND_299[63:0];
  _RAND_300 = {2{`RANDOM}};
  record_wdata1_44 = _RAND_300[63:0];
  _RAND_301 = {2{`RANDOM}};
  record_wdata1_45 = _RAND_301[63:0];
  _RAND_302 = {2{`RANDOM}};
  record_wdata1_46 = _RAND_302[63:0];
  _RAND_303 = {2{`RANDOM}};
  record_wdata1_47 = _RAND_303[63:0];
  _RAND_304 = {2{`RANDOM}};
  record_wdata1_48 = _RAND_304[63:0];
  _RAND_305 = {2{`RANDOM}};
  record_wdata1_49 = _RAND_305[63:0];
  _RAND_306 = {2{`RANDOM}};
  record_wdata1_50 = _RAND_306[63:0];
  _RAND_307 = {2{`RANDOM}};
  record_wdata1_51 = _RAND_307[63:0];
  _RAND_308 = {2{`RANDOM}};
  record_wdata1_52 = _RAND_308[63:0];
  _RAND_309 = {2{`RANDOM}};
  record_wdata1_53 = _RAND_309[63:0];
  _RAND_310 = {2{`RANDOM}};
  record_wdata1_54 = _RAND_310[63:0];
  _RAND_311 = {2{`RANDOM}};
  record_wdata1_55 = _RAND_311[63:0];
  _RAND_312 = {2{`RANDOM}};
  record_wdata1_56 = _RAND_312[63:0];
  _RAND_313 = {2{`RANDOM}};
  record_wdata1_57 = _RAND_313[63:0];
  _RAND_314 = {2{`RANDOM}};
  record_wdata1_58 = _RAND_314[63:0];
  _RAND_315 = {2{`RANDOM}};
  record_wdata1_59 = _RAND_315[63:0];
  _RAND_316 = {2{`RANDOM}};
  record_wdata1_60 = _RAND_316[63:0];
  _RAND_317 = {2{`RANDOM}};
  record_wdata1_61 = _RAND_317[63:0];
  _RAND_318 = {2{`RANDOM}};
  record_wdata1_62 = _RAND_318[63:0];
  _RAND_319 = {2{`RANDOM}};
  record_wdata1_63 = _RAND_319[63:0];
  _RAND_320 = {2{`RANDOM}};
  record_wdata1_64 = _RAND_320[63:0];
  _RAND_321 = {2{`RANDOM}};
  record_wdata1_65 = _RAND_321[63:0];
  _RAND_322 = {2{`RANDOM}};
  record_wdata1_66 = _RAND_322[63:0];
  _RAND_323 = {2{`RANDOM}};
  record_wdata1_67 = _RAND_323[63:0];
  _RAND_324 = {2{`RANDOM}};
  record_wdata1_68 = _RAND_324[63:0];
  _RAND_325 = {2{`RANDOM}};
  record_wdata1_69 = _RAND_325[63:0];
  _RAND_326 = {2{`RANDOM}};
  record_wdata1_70 = _RAND_326[63:0];
  _RAND_327 = {2{`RANDOM}};
  record_wdata1_71 = _RAND_327[63:0];
  _RAND_328 = {2{`RANDOM}};
  record_wdata1_72 = _RAND_328[63:0];
  _RAND_329 = {2{`RANDOM}};
  record_wdata1_73 = _RAND_329[63:0];
  _RAND_330 = {2{`RANDOM}};
  record_wdata1_74 = _RAND_330[63:0];
  _RAND_331 = {2{`RANDOM}};
  record_wdata1_75 = _RAND_331[63:0];
  _RAND_332 = {2{`RANDOM}};
  record_wdata1_76 = _RAND_332[63:0];
  _RAND_333 = {2{`RANDOM}};
  record_wdata1_77 = _RAND_333[63:0];
  _RAND_334 = {2{`RANDOM}};
  record_wdata1_78 = _RAND_334[63:0];
  _RAND_335 = {2{`RANDOM}};
  record_wdata1_79 = _RAND_335[63:0];
  _RAND_336 = {2{`RANDOM}};
  record_wdata1_80 = _RAND_336[63:0];
  _RAND_337 = {2{`RANDOM}};
  record_wdata1_81 = _RAND_337[63:0];
  _RAND_338 = {2{`RANDOM}};
  record_wdata1_82 = _RAND_338[63:0];
  _RAND_339 = {2{`RANDOM}};
  record_wdata1_83 = _RAND_339[63:0];
  _RAND_340 = {2{`RANDOM}};
  record_wdata1_84 = _RAND_340[63:0];
  _RAND_341 = {2{`RANDOM}};
  record_wdata1_85 = _RAND_341[63:0];
  _RAND_342 = {2{`RANDOM}};
  record_wdata1_86 = _RAND_342[63:0];
  _RAND_343 = {2{`RANDOM}};
  record_wdata1_87 = _RAND_343[63:0];
  _RAND_344 = {2{`RANDOM}};
  record_wdata1_88 = _RAND_344[63:0];
  _RAND_345 = {2{`RANDOM}};
  record_wdata1_89 = _RAND_345[63:0];
  _RAND_346 = {2{`RANDOM}};
  record_wdata1_90 = _RAND_346[63:0];
  _RAND_347 = {2{`RANDOM}};
  record_wdata1_91 = _RAND_347[63:0];
  _RAND_348 = {2{`RANDOM}};
  record_wdata1_92 = _RAND_348[63:0];
  _RAND_349 = {2{`RANDOM}};
  record_wdata1_93 = _RAND_349[63:0];
  _RAND_350 = {2{`RANDOM}};
  record_wdata1_94 = _RAND_350[63:0];
  _RAND_351 = {2{`RANDOM}};
  record_wdata1_95 = _RAND_351[63:0];
  _RAND_352 = {2{`RANDOM}};
  record_wdata1_96 = _RAND_352[63:0];
  _RAND_353 = {2{`RANDOM}};
  record_wdata1_97 = _RAND_353[63:0];
  _RAND_354 = {2{`RANDOM}};
  record_wdata1_98 = _RAND_354[63:0];
  _RAND_355 = {2{`RANDOM}};
  record_wdata1_99 = _RAND_355[63:0];
  _RAND_356 = {2{`RANDOM}};
  record_wdata1_100 = _RAND_356[63:0];
  _RAND_357 = {2{`RANDOM}};
  record_wdata1_101 = _RAND_357[63:0];
  _RAND_358 = {2{`RANDOM}};
  record_wdata1_102 = _RAND_358[63:0];
  _RAND_359 = {2{`RANDOM}};
  record_wdata1_103 = _RAND_359[63:0];
  _RAND_360 = {2{`RANDOM}};
  record_wdata1_104 = _RAND_360[63:0];
  _RAND_361 = {2{`RANDOM}};
  record_wdata1_105 = _RAND_361[63:0];
  _RAND_362 = {2{`RANDOM}};
  record_wdata1_106 = _RAND_362[63:0];
  _RAND_363 = {2{`RANDOM}};
  record_wdata1_107 = _RAND_363[63:0];
  _RAND_364 = {2{`RANDOM}};
  record_wdata1_108 = _RAND_364[63:0];
  _RAND_365 = {2{`RANDOM}};
  record_wdata1_109 = _RAND_365[63:0];
  _RAND_366 = {2{`RANDOM}};
  record_wdata1_110 = _RAND_366[63:0];
  _RAND_367 = {2{`RANDOM}};
  record_wdata1_111 = _RAND_367[63:0];
  _RAND_368 = {2{`RANDOM}};
  record_wdata1_112 = _RAND_368[63:0];
  _RAND_369 = {2{`RANDOM}};
  record_wdata1_113 = _RAND_369[63:0];
  _RAND_370 = {2{`RANDOM}};
  record_wdata1_114 = _RAND_370[63:0];
  _RAND_371 = {2{`RANDOM}};
  record_wdata1_115 = _RAND_371[63:0];
  _RAND_372 = {2{`RANDOM}};
  record_wdata1_116 = _RAND_372[63:0];
  _RAND_373 = {2{`RANDOM}};
  record_wdata1_117 = _RAND_373[63:0];
  _RAND_374 = {2{`RANDOM}};
  record_wdata1_118 = _RAND_374[63:0];
  _RAND_375 = {2{`RANDOM}};
  record_wdata1_119 = _RAND_375[63:0];
  _RAND_376 = {2{`RANDOM}};
  record_wdata1_120 = _RAND_376[63:0];
  _RAND_377 = {2{`RANDOM}};
  record_wdata1_121 = _RAND_377[63:0];
  _RAND_378 = {2{`RANDOM}};
  record_wdata1_122 = _RAND_378[63:0];
  _RAND_379 = {2{`RANDOM}};
  record_wdata1_123 = _RAND_379[63:0];
  _RAND_380 = {2{`RANDOM}};
  record_wdata1_124 = _RAND_380[63:0];
  _RAND_381 = {2{`RANDOM}};
  record_wdata1_125 = _RAND_381[63:0];
  _RAND_382 = {2{`RANDOM}};
  record_wdata1_126 = _RAND_382[63:0];
  _RAND_383 = {2{`RANDOM}};
  record_wdata1_127 = _RAND_383[63:0];
  _RAND_384 = {1{`RANDOM}};
  record_wstrb1_0 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  record_wstrb1_1 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  record_wstrb1_2 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  record_wstrb1_3 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  record_wstrb1_4 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  record_wstrb1_5 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  record_wstrb1_6 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  record_wstrb1_7 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  record_wstrb1_8 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  record_wstrb1_9 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  record_wstrb1_10 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  record_wstrb1_11 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  record_wstrb1_12 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  record_wstrb1_13 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  record_wstrb1_14 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  record_wstrb1_15 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  record_wstrb1_16 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  record_wstrb1_17 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  record_wstrb1_18 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  record_wstrb1_19 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  record_wstrb1_20 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  record_wstrb1_21 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  record_wstrb1_22 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  record_wstrb1_23 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  record_wstrb1_24 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  record_wstrb1_25 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  record_wstrb1_26 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  record_wstrb1_27 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  record_wstrb1_28 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  record_wstrb1_29 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  record_wstrb1_30 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  record_wstrb1_31 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  record_wstrb1_32 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  record_wstrb1_33 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  record_wstrb1_34 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  record_wstrb1_35 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  record_wstrb1_36 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  record_wstrb1_37 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  record_wstrb1_38 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  record_wstrb1_39 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  record_wstrb1_40 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  record_wstrb1_41 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  record_wstrb1_42 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  record_wstrb1_43 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  record_wstrb1_44 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  record_wstrb1_45 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  record_wstrb1_46 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  record_wstrb1_47 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  record_wstrb1_48 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  record_wstrb1_49 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  record_wstrb1_50 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  record_wstrb1_51 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  record_wstrb1_52 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  record_wstrb1_53 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  record_wstrb1_54 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  record_wstrb1_55 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  record_wstrb1_56 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  record_wstrb1_57 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  record_wstrb1_58 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  record_wstrb1_59 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  record_wstrb1_60 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  record_wstrb1_61 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  record_wstrb1_62 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  record_wstrb1_63 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  record_wstrb1_64 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  record_wstrb1_65 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  record_wstrb1_66 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  record_wstrb1_67 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  record_wstrb1_68 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  record_wstrb1_69 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  record_wstrb1_70 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  record_wstrb1_71 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  record_wstrb1_72 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  record_wstrb1_73 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  record_wstrb1_74 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  record_wstrb1_75 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  record_wstrb1_76 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  record_wstrb1_77 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  record_wstrb1_78 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  record_wstrb1_79 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  record_wstrb1_80 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  record_wstrb1_81 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  record_wstrb1_82 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  record_wstrb1_83 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  record_wstrb1_84 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  record_wstrb1_85 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  record_wstrb1_86 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  record_wstrb1_87 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  record_wstrb1_88 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  record_wstrb1_89 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  record_wstrb1_90 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  record_wstrb1_91 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  record_wstrb1_92 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  record_wstrb1_93 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  record_wstrb1_94 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  record_wstrb1_95 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  record_wstrb1_96 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  record_wstrb1_97 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  record_wstrb1_98 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  record_wstrb1_99 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  record_wstrb1_100 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  record_wstrb1_101 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  record_wstrb1_102 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  record_wstrb1_103 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  record_wstrb1_104 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  record_wstrb1_105 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  record_wstrb1_106 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  record_wstrb1_107 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  record_wstrb1_108 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  record_wstrb1_109 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  record_wstrb1_110 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  record_wstrb1_111 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  record_wstrb1_112 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  record_wstrb1_113 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  record_wstrb1_114 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  record_wstrb1_115 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  record_wstrb1_116 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  record_wstrb1_117 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  record_wstrb1_118 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  record_wstrb1_119 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  record_wstrb1_120 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  record_wstrb1_121 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  record_wstrb1_122 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  record_wstrb1_123 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  record_wstrb1_124 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  record_wstrb1_125 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  record_wstrb1_126 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  record_wstrb1_127 = _RAND_511[7:0];
  _RAND_512 = {2{`RANDOM}};
  record_pc_0 = _RAND_512[63:0];
  _RAND_513 = {2{`RANDOM}};
  record_pc_1 = _RAND_513[63:0];
  _RAND_514 = {2{`RANDOM}};
  record_pc_2 = _RAND_514[63:0];
  _RAND_515 = {2{`RANDOM}};
  record_pc_3 = _RAND_515[63:0];
  _RAND_516 = {2{`RANDOM}};
  record_pc_4 = _RAND_516[63:0];
  _RAND_517 = {2{`RANDOM}};
  record_pc_5 = _RAND_517[63:0];
  _RAND_518 = {2{`RANDOM}};
  record_pc_6 = _RAND_518[63:0];
  _RAND_519 = {2{`RANDOM}};
  record_pc_7 = _RAND_519[63:0];
  _RAND_520 = {2{`RANDOM}};
  record_pc_8 = _RAND_520[63:0];
  _RAND_521 = {2{`RANDOM}};
  record_pc_9 = _RAND_521[63:0];
  _RAND_522 = {2{`RANDOM}};
  record_pc_10 = _RAND_522[63:0];
  _RAND_523 = {2{`RANDOM}};
  record_pc_11 = _RAND_523[63:0];
  _RAND_524 = {2{`RANDOM}};
  record_pc_12 = _RAND_524[63:0];
  _RAND_525 = {2{`RANDOM}};
  record_pc_13 = _RAND_525[63:0];
  _RAND_526 = {2{`RANDOM}};
  record_pc_14 = _RAND_526[63:0];
  _RAND_527 = {2{`RANDOM}};
  record_pc_15 = _RAND_527[63:0];
  _RAND_528 = {2{`RANDOM}};
  record_pc_16 = _RAND_528[63:0];
  _RAND_529 = {2{`RANDOM}};
  record_pc_17 = _RAND_529[63:0];
  _RAND_530 = {2{`RANDOM}};
  record_pc_18 = _RAND_530[63:0];
  _RAND_531 = {2{`RANDOM}};
  record_pc_19 = _RAND_531[63:0];
  _RAND_532 = {2{`RANDOM}};
  record_pc_20 = _RAND_532[63:0];
  _RAND_533 = {2{`RANDOM}};
  record_pc_21 = _RAND_533[63:0];
  _RAND_534 = {2{`RANDOM}};
  record_pc_22 = _RAND_534[63:0];
  _RAND_535 = {2{`RANDOM}};
  record_pc_23 = _RAND_535[63:0];
  _RAND_536 = {2{`RANDOM}};
  record_pc_24 = _RAND_536[63:0];
  _RAND_537 = {2{`RANDOM}};
  record_pc_25 = _RAND_537[63:0];
  _RAND_538 = {2{`RANDOM}};
  record_pc_26 = _RAND_538[63:0];
  _RAND_539 = {2{`RANDOM}};
  record_pc_27 = _RAND_539[63:0];
  _RAND_540 = {2{`RANDOM}};
  record_pc_28 = _RAND_540[63:0];
  _RAND_541 = {2{`RANDOM}};
  record_pc_29 = _RAND_541[63:0];
  _RAND_542 = {2{`RANDOM}};
  record_pc_30 = _RAND_542[63:0];
  _RAND_543 = {2{`RANDOM}};
  record_pc_31 = _RAND_543[63:0];
  _RAND_544 = {2{`RANDOM}};
  record_pc_32 = _RAND_544[63:0];
  _RAND_545 = {2{`RANDOM}};
  record_pc_33 = _RAND_545[63:0];
  _RAND_546 = {2{`RANDOM}};
  record_pc_34 = _RAND_546[63:0];
  _RAND_547 = {2{`RANDOM}};
  record_pc_35 = _RAND_547[63:0];
  _RAND_548 = {2{`RANDOM}};
  record_pc_36 = _RAND_548[63:0];
  _RAND_549 = {2{`RANDOM}};
  record_pc_37 = _RAND_549[63:0];
  _RAND_550 = {2{`RANDOM}};
  record_pc_38 = _RAND_550[63:0];
  _RAND_551 = {2{`RANDOM}};
  record_pc_39 = _RAND_551[63:0];
  _RAND_552 = {2{`RANDOM}};
  record_pc_40 = _RAND_552[63:0];
  _RAND_553 = {2{`RANDOM}};
  record_pc_41 = _RAND_553[63:0];
  _RAND_554 = {2{`RANDOM}};
  record_pc_42 = _RAND_554[63:0];
  _RAND_555 = {2{`RANDOM}};
  record_pc_43 = _RAND_555[63:0];
  _RAND_556 = {2{`RANDOM}};
  record_pc_44 = _RAND_556[63:0];
  _RAND_557 = {2{`RANDOM}};
  record_pc_45 = _RAND_557[63:0];
  _RAND_558 = {2{`RANDOM}};
  record_pc_46 = _RAND_558[63:0];
  _RAND_559 = {2{`RANDOM}};
  record_pc_47 = _RAND_559[63:0];
  _RAND_560 = {2{`RANDOM}};
  record_pc_48 = _RAND_560[63:0];
  _RAND_561 = {2{`RANDOM}};
  record_pc_49 = _RAND_561[63:0];
  _RAND_562 = {2{`RANDOM}};
  record_pc_50 = _RAND_562[63:0];
  _RAND_563 = {2{`RANDOM}};
  record_pc_51 = _RAND_563[63:0];
  _RAND_564 = {2{`RANDOM}};
  record_pc_52 = _RAND_564[63:0];
  _RAND_565 = {2{`RANDOM}};
  record_pc_53 = _RAND_565[63:0];
  _RAND_566 = {2{`RANDOM}};
  record_pc_54 = _RAND_566[63:0];
  _RAND_567 = {2{`RANDOM}};
  record_pc_55 = _RAND_567[63:0];
  _RAND_568 = {2{`RANDOM}};
  record_pc_56 = _RAND_568[63:0];
  _RAND_569 = {2{`RANDOM}};
  record_pc_57 = _RAND_569[63:0];
  _RAND_570 = {2{`RANDOM}};
  record_pc_58 = _RAND_570[63:0];
  _RAND_571 = {2{`RANDOM}};
  record_pc_59 = _RAND_571[63:0];
  _RAND_572 = {2{`RANDOM}};
  record_pc_60 = _RAND_572[63:0];
  _RAND_573 = {2{`RANDOM}};
  record_pc_61 = _RAND_573[63:0];
  _RAND_574 = {2{`RANDOM}};
  record_pc_62 = _RAND_574[63:0];
  _RAND_575 = {2{`RANDOM}};
  record_pc_63 = _RAND_575[63:0];
  _RAND_576 = {2{`RANDOM}};
  record_pc_64 = _RAND_576[63:0];
  _RAND_577 = {2{`RANDOM}};
  record_pc_65 = _RAND_577[63:0];
  _RAND_578 = {2{`RANDOM}};
  record_pc_66 = _RAND_578[63:0];
  _RAND_579 = {2{`RANDOM}};
  record_pc_67 = _RAND_579[63:0];
  _RAND_580 = {2{`RANDOM}};
  record_pc_68 = _RAND_580[63:0];
  _RAND_581 = {2{`RANDOM}};
  record_pc_69 = _RAND_581[63:0];
  _RAND_582 = {2{`RANDOM}};
  record_pc_70 = _RAND_582[63:0];
  _RAND_583 = {2{`RANDOM}};
  record_pc_71 = _RAND_583[63:0];
  _RAND_584 = {2{`RANDOM}};
  record_pc_72 = _RAND_584[63:0];
  _RAND_585 = {2{`RANDOM}};
  record_pc_73 = _RAND_585[63:0];
  _RAND_586 = {2{`RANDOM}};
  record_pc_74 = _RAND_586[63:0];
  _RAND_587 = {2{`RANDOM}};
  record_pc_75 = _RAND_587[63:0];
  _RAND_588 = {2{`RANDOM}};
  record_pc_76 = _RAND_588[63:0];
  _RAND_589 = {2{`RANDOM}};
  record_pc_77 = _RAND_589[63:0];
  _RAND_590 = {2{`RANDOM}};
  record_pc_78 = _RAND_590[63:0];
  _RAND_591 = {2{`RANDOM}};
  record_pc_79 = _RAND_591[63:0];
  _RAND_592 = {2{`RANDOM}};
  record_pc_80 = _RAND_592[63:0];
  _RAND_593 = {2{`RANDOM}};
  record_pc_81 = _RAND_593[63:0];
  _RAND_594 = {2{`RANDOM}};
  record_pc_82 = _RAND_594[63:0];
  _RAND_595 = {2{`RANDOM}};
  record_pc_83 = _RAND_595[63:0];
  _RAND_596 = {2{`RANDOM}};
  record_pc_84 = _RAND_596[63:0];
  _RAND_597 = {2{`RANDOM}};
  record_pc_85 = _RAND_597[63:0];
  _RAND_598 = {2{`RANDOM}};
  record_pc_86 = _RAND_598[63:0];
  _RAND_599 = {2{`RANDOM}};
  record_pc_87 = _RAND_599[63:0];
  _RAND_600 = {2{`RANDOM}};
  record_pc_88 = _RAND_600[63:0];
  _RAND_601 = {2{`RANDOM}};
  record_pc_89 = _RAND_601[63:0];
  _RAND_602 = {2{`RANDOM}};
  record_pc_90 = _RAND_602[63:0];
  _RAND_603 = {2{`RANDOM}};
  record_pc_91 = _RAND_603[63:0];
  _RAND_604 = {2{`RANDOM}};
  record_pc_92 = _RAND_604[63:0];
  _RAND_605 = {2{`RANDOM}};
  record_pc_93 = _RAND_605[63:0];
  _RAND_606 = {2{`RANDOM}};
  record_pc_94 = _RAND_606[63:0];
  _RAND_607 = {2{`RANDOM}};
  record_pc_95 = _RAND_607[63:0];
  _RAND_608 = {2{`RANDOM}};
  record_pc_96 = _RAND_608[63:0];
  _RAND_609 = {2{`RANDOM}};
  record_pc_97 = _RAND_609[63:0];
  _RAND_610 = {2{`RANDOM}};
  record_pc_98 = _RAND_610[63:0];
  _RAND_611 = {2{`RANDOM}};
  record_pc_99 = _RAND_611[63:0];
  _RAND_612 = {2{`RANDOM}};
  record_pc_100 = _RAND_612[63:0];
  _RAND_613 = {2{`RANDOM}};
  record_pc_101 = _RAND_613[63:0];
  _RAND_614 = {2{`RANDOM}};
  record_pc_102 = _RAND_614[63:0];
  _RAND_615 = {2{`RANDOM}};
  record_pc_103 = _RAND_615[63:0];
  _RAND_616 = {2{`RANDOM}};
  record_pc_104 = _RAND_616[63:0];
  _RAND_617 = {2{`RANDOM}};
  record_pc_105 = _RAND_617[63:0];
  _RAND_618 = {2{`RANDOM}};
  record_pc_106 = _RAND_618[63:0];
  _RAND_619 = {2{`RANDOM}};
  record_pc_107 = _RAND_619[63:0];
  _RAND_620 = {2{`RANDOM}};
  record_pc_108 = _RAND_620[63:0];
  _RAND_621 = {2{`RANDOM}};
  record_pc_109 = _RAND_621[63:0];
  _RAND_622 = {2{`RANDOM}};
  record_pc_110 = _RAND_622[63:0];
  _RAND_623 = {2{`RANDOM}};
  record_pc_111 = _RAND_623[63:0];
  _RAND_624 = {2{`RANDOM}};
  record_pc_112 = _RAND_624[63:0];
  _RAND_625 = {2{`RANDOM}};
  record_pc_113 = _RAND_625[63:0];
  _RAND_626 = {2{`RANDOM}};
  record_pc_114 = _RAND_626[63:0];
  _RAND_627 = {2{`RANDOM}};
  record_pc_115 = _RAND_627[63:0];
  _RAND_628 = {2{`RANDOM}};
  record_pc_116 = _RAND_628[63:0];
  _RAND_629 = {2{`RANDOM}};
  record_pc_117 = _RAND_629[63:0];
  _RAND_630 = {2{`RANDOM}};
  record_pc_118 = _RAND_630[63:0];
  _RAND_631 = {2{`RANDOM}};
  record_pc_119 = _RAND_631[63:0];
  _RAND_632 = {2{`RANDOM}};
  record_pc_120 = _RAND_632[63:0];
  _RAND_633 = {2{`RANDOM}};
  record_pc_121 = _RAND_633[63:0];
  _RAND_634 = {2{`RANDOM}};
  record_pc_122 = _RAND_634[63:0];
  _RAND_635 = {2{`RANDOM}};
  record_pc_123 = _RAND_635[63:0];
  _RAND_636 = {2{`RANDOM}};
  record_pc_124 = _RAND_636[63:0];
  _RAND_637 = {2{`RANDOM}};
  record_pc_125 = _RAND_637[63:0];
  _RAND_638 = {2{`RANDOM}};
  record_pc_126 = _RAND_638[63:0];
  _RAND_639 = {2{`RANDOM}};
  record_pc_127 = _RAND_639[63:0];
  _RAND_640 = {1{`RANDOM}};
  record_addr_0 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  record_addr_1 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  record_addr_2 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  record_addr_3 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  record_addr_4 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  record_addr_5 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  record_addr_6 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  record_addr_7 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  record_addr_8 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  record_addr_9 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  record_addr_10 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  record_addr_11 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  record_addr_12 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  record_addr_13 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  record_addr_14 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  record_addr_15 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  record_addr_16 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  record_addr_17 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  record_addr_18 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  record_addr_19 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  record_addr_20 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  record_addr_21 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  record_addr_22 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  record_addr_23 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  record_addr_24 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  record_addr_25 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  record_addr_26 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  record_addr_27 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  record_addr_28 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  record_addr_29 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  record_addr_30 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  record_addr_31 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  record_addr_32 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  record_addr_33 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  record_addr_34 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  record_addr_35 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  record_addr_36 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  record_addr_37 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  record_addr_38 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  record_addr_39 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  record_addr_40 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  record_addr_41 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  record_addr_42 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  record_addr_43 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  record_addr_44 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  record_addr_45 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  record_addr_46 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  record_addr_47 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  record_addr_48 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  record_addr_49 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  record_addr_50 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  record_addr_51 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  record_addr_52 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  record_addr_53 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  record_addr_54 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  record_addr_55 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  record_addr_56 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  record_addr_57 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  record_addr_58 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  record_addr_59 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  record_addr_60 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  record_addr_61 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  record_addr_62 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  record_addr_63 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  record_addr_64 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  record_addr_65 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  record_addr_66 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  record_addr_67 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  record_addr_68 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  record_addr_69 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  record_addr_70 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  record_addr_71 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  record_addr_72 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  record_addr_73 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  record_addr_74 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  record_addr_75 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  record_addr_76 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  record_addr_77 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  record_addr_78 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  record_addr_79 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  record_addr_80 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  record_addr_81 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  record_addr_82 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  record_addr_83 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  record_addr_84 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  record_addr_85 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  record_addr_86 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  record_addr_87 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  record_addr_88 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  record_addr_89 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  record_addr_90 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  record_addr_91 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  record_addr_92 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  record_addr_93 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  record_addr_94 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  record_addr_95 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  record_addr_96 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  record_addr_97 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  record_addr_98 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  record_addr_99 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  record_addr_100 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  record_addr_101 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  record_addr_102 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  record_addr_103 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  record_addr_104 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  record_addr_105 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  record_addr_106 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  record_addr_107 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  record_addr_108 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  record_addr_109 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  record_addr_110 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  record_addr_111 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  record_addr_112 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  record_addr_113 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  record_addr_114 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  record_addr_115 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  record_addr_116 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  record_addr_117 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  record_addr_118 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  record_addr_119 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  record_addr_120 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  record_addr_121 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  record_addr_122 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  record_addr_123 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  record_addr_124 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  record_addr_125 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  record_addr_126 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  record_addr_127 = _RAND_767[31:0];
  _RAND_768 = {2{`RANDOM}};
  record_olddata_0 = _RAND_768[63:0];
  _RAND_769 = {2{`RANDOM}};
  record_olddata_1 = _RAND_769[63:0];
  _RAND_770 = {2{`RANDOM}};
  record_olddata_2 = _RAND_770[63:0];
  _RAND_771 = {2{`RANDOM}};
  record_olddata_3 = _RAND_771[63:0];
  _RAND_772 = {2{`RANDOM}};
  record_olddata_4 = _RAND_772[63:0];
  _RAND_773 = {2{`RANDOM}};
  record_olddata_5 = _RAND_773[63:0];
  _RAND_774 = {2{`RANDOM}};
  record_olddata_6 = _RAND_774[63:0];
  _RAND_775 = {2{`RANDOM}};
  record_olddata_7 = _RAND_775[63:0];
  _RAND_776 = {2{`RANDOM}};
  record_olddata_8 = _RAND_776[63:0];
  _RAND_777 = {2{`RANDOM}};
  record_olddata_9 = _RAND_777[63:0];
  _RAND_778 = {2{`RANDOM}};
  record_olddata_10 = _RAND_778[63:0];
  _RAND_779 = {2{`RANDOM}};
  record_olddata_11 = _RAND_779[63:0];
  _RAND_780 = {2{`RANDOM}};
  record_olddata_12 = _RAND_780[63:0];
  _RAND_781 = {2{`RANDOM}};
  record_olddata_13 = _RAND_781[63:0];
  _RAND_782 = {2{`RANDOM}};
  record_olddata_14 = _RAND_782[63:0];
  _RAND_783 = {2{`RANDOM}};
  record_olddata_15 = _RAND_783[63:0];
  _RAND_784 = {2{`RANDOM}};
  record_olddata_16 = _RAND_784[63:0];
  _RAND_785 = {2{`RANDOM}};
  record_olddata_17 = _RAND_785[63:0];
  _RAND_786 = {2{`RANDOM}};
  record_olddata_18 = _RAND_786[63:0];
  _RAND_787 = {2{`RANDOM}};
  record_olddata_19 = _RAND_787[63:0];
  _RAND_788 = {2{`RANDOM}};
  record_olddata_20 = _RAND_788[63:0];
  _RAND_789 = {2{`RANDOM}};
  record_olddata_21 = _RAND_789[63:0];
  _RAND_790 = {2{`RANDOM}};
  record_olddata_22 = _RAND_790[63:0];
  _RAND_791 = {2{`RANDOM}};
  record_olddata_23 = _RAND_791[63:0];
  _RAND_792 = {2{`RANDOM}};
  record_olddata_24 = _RAND_792[63:0];
  _RAND_793 = {2{`RANDOM}};
  record_olddata_25 = _RAND_793[63:0];
  _RAND_794 = {2{`RANDOM}};
  record_olddata_26 = _RAND_794[63:0];
  _RAND_795 = {2{`RANDOM}};
  record_olddata_27 = _RAND_795[63:0];
  _RAND_796 = {2{`RANDOM}};
  record_olddata_28 = _RAND_796[63:0];
  _RAND_797 = {2{`RANDOM}};
  record_olddata_29 = _RAND_797[63:0];
  _RAND_798 = {2{`RANDOM}};
  record_olddata_30 = _RAND_798[63:0];
  _RAND_799 = {2{`RANDOM}};
  record_olddata_31 = _RAND_799[63:0];
  _RAND_800 = {2{`RANDOM}};
  record_olddata_32 = _RAND_800[63:0];
  _RAND_801 = {2{`RANDOM}};
  record_olddata_33 = _RAND_801[63:0];
  _RAND_802 = {2{`RANDOM}};
  record_olddata_34 = _RAND_802[63:0];
  _RAND_803 = {2{`RANDOM}};
  record_olddata_35 = _RAND_803[63:0];
  _RAND_804 = {2{`RANDOM}};
  record_olddata_36 = _RAND_804[63:0];
  _RAND_805 = {2{`RANDOM}};
  record_olddata_37 = _RAND_805[63:0];
  _RAND_806 = {2{`RANDOM}};
  record_olddata_38 = _RAND_806[63:0];
  _RAND_807 = {2{`RANDOM}};
  record_olddata_39 = _RAND_807[63:0];
  _RAND_808 = {2{`RANDOM}};
  record_olddata_40 = _RAND_808[63:0];
  _RAND_809 = {2{`RANDOM}};
  record_olddata_41 = _RAND_809[63:0];
  _RAND_810 = {2{`RANDOM}};
  record_olddata_42 = _RAND_810[63:0];
  _RAND_811 = {2{`RANDOM}};
  record_olddata_43 = _RAND_811[63:0];
  _RAND_812 = {2{`RANDOM}};
  record_olddata_44 = _RAND_812[63:0];
  _RAND_813 = {2{`RANDOM}};
  record_olddata_45 = _RAND_813[63:0];
  _RAND_814 = {2{`RANDOM}};
  record_olddata_46 = _RAND_814[63:0];
  _RAND_815 = {2{`RANDOM}};
  record_olddata_47 = _RAND_815[63:0];
  _RAND_816 = {2{`RANDOM}};
  record_olddata_48 = _RAND_816[63:0];
  _RAND_817 = {2{`RANDOM}};
  record_olddata_49 = _RAND_817[63:0];
  _RAND_818 = {2{`RANDOM}};
  record_olddata_50 = _RAND_818[63:0];
  _RAND_819 = {2{`RANDOM}};
  record_olddata_51 = _RAND_819[63:0];
  _RAND_820 = {2{`RANDOM}};
  record_olddata_52 = _RAND_820[63:0];
  _RAND_821 = {2{`RANDOM}};
  record_olddata_53 = _RAND_821[63:0];
  _RAND_822 = {2{`RANDOM}};
  record_olddata_54 = _RAND_822[63:0];
  _RAND_823 = {2{`RANDOM}};
  record_olddata_55 = _RAND_823[63:0];
  _RAND_824 = {2{`RANDOM}};
  record_olddata_56 = _RAND_824[63:0];
  _RAND_825 = {2{`RANDOM}};
  record_olddata_57 = _RAND_825[63:0];
  _RAND_826 = {2{`RANDOM}};
  record_olddata_58 = _RAND_826[63:0];
  _RAND_827 = {2{`RANDOM}};
  record_olddata_59 = _RAND_827[63:0];
  _RAND_828 = {2{`RANDOM}};
  record_olddata_60 = _RAND_828[63:0];
  _RAND_829 = {2{`RANDOM}};
  record_olddata_61 = _RAND_829[63:0];
  _RAND_830 = {2{`RANDOM}};
  record_olddata_62 = _RAND_830[63:0];
  _RAND_831 = {2{`RANDOM}};
  record_olddata_63 = _RAND_831[63:0];
  _RAND_832 = {2{`RANDOM}};
  record_olddata_64 = _RAND_832[63:0];
  _RAND_833 = {2{`RANDOM}};
  record_olddata_65 = _RAND_833[63:0];
  _RAND_834 = {2{`RANDOM}};
  record_olddata_66 = _RAND_834[63:0];
  _RAND_835 = {2{`RANDOM}};
  record_olddata_67 = _RAND_835[63:0];
  _RAND_836 = {2{`RANDOM}};
  record_olddata_68 = _RAND_836[63:0];
  _RAND_837 = {2{`RANDOM}};
  record_olddata_69 = _RAND_837[63:0];
  _RAND_838 = {2{`RANDOM}};
  record_olddata_70 = _RAND_838[63:0];
  _RAND_839 = {2{`RANDOM}};
  record_olddata_71 = _RAND_839[63:0];
  _RAND_840 = {2{`RANDOM}};
  record_olddata_72 = _RAND_840[63:0];
  _RAND_841 = {2{`RANDOM}};
  record_olddata_73 = _RAND_841[63:0];
  _RAND_842 = {2{`RANDOM}};
  record_olddata_74 = _RAND_842[63:0];
  _RAND_843 = {2{`RANDOM}};
  record_olddata_75 = _RAND_843[63:0];
  _RAND_844 = {2{`RANDOM}};
  record_olddata_76 = _RAND_844[63:0];
  _RAND_845 = {2{`RANDOM}};
  record_olddata_77 = _RAND_845[63:0];
  _RAND_846 = {2{`RANDOM}};
  record_olddata_78 = _RAND_846[63:0];
  _RAND_847 = {2{`RANDOM}};
  record_olddata_79 = _RAND_847[63:0];
  _RAND_848 = {2{`RANDOM}};
  record_olddata_80 = _RAND_848[63:0];
  _RAND_849 = {2{`RANDOM}};
  record_olddata_81 = _RAND_849[63:0];
  _RAND_850 = {2{`RANDOM}};
  record_olddata_82 = _RAND_850[63:0];
  _RAND_851 = {2{`RANDOM}};
  record_olddata_83 = _RAND_851[63:0];
  _RAND_852 = {2{`RANDOM}};
  record_olddata_84 = _RAND_852[63:0];
  _RAND_853 = {2{`RANDOM}};
  record_olddata_85 = _RAND_853[63:0];
  _RAND_854 = {2{`RANDOM}};
  record_olddata_86 = _RAND_854[63:0];
  _RAND_855 = {2{`RANDOM}};
  record_olddata_87 = _RAND_855[63:0];
  _RAND_856 = {2{`RANDOM}};
  record_olddata_88 = _RAND_856[63:0];
  _RAND_857 = {2{`RANDOM}};
  record_olddata_89 = _RAND_857[63:0];
  _RAND_858 = {2{`RANDOM}};
  record_olddata_90 = _RAND_858[63:0];
  _RAND_859 = {2{`RANDOM}};
  record_olddata_91 = _RAND_859[63:0];
  _RAND_860 = {2{`RANDOM}};
  record_olddata_92 = _RAND_860[63:0];
  _RAND_861 = {2{`RANDOM}};
  record_olddata_93 = _RAND_861[63:0];
  _RAND_862 = {2{`RANDOM}};
  record_olddata_94 = _RAND_862[63:0];
  _RAND_863 = {2{`RANDOM}};
  record_olddata_95 = _RAND_863[63:0];
  _RAND_864 = {2{`RANDOM}};
  record_olddata_96 = _RAND_864[63:0];
  _RAND_865 = {2{`RANDOM}};
  record_olddata_97 = _RAND_865[63:0];
  _RAND_866 = {2{`RANDOM}};
  record_olddata_98 = _RAND_866[63:0];
  _RAND_867 = {2{`RANDOM}};
  record_olddata_99 = _RAND_867[63:0];
  _RAND_868 = {2{`RANDOM}};
  record_olddata_100 = _RAND_868[63:0];
  _RAND_869 = {2{`RANDOM}};
  record_olddata_101 = _RAND_869[63:0];
  _RAND_870 = {2{`RANDOM}};
  record_olddata_102 = _RAND_870[63:0];
  _RAND_871 = {2{`RANDOM}};
  record_olddata_103 = _RAND_871[63:0];
  _RAND_872 = {2{`RANDOM}};
  record_olddata_104 = _RAND_872[63:0];
  _RAND_873 = {2{`RANDOM}};
  record_olddata_105 = _RAND_873[63:0];
  _RAND_874 = {2{`RANDOM}};
  record_olddata_106 = _RAND_874[63:0];
  _RAND_875 = {2{`RANDOM}};
  record_olddata_107 = _RAND_875[63:0];
  _RAND_876 = {2{`RANDOM}};
  record_olddata_108 = _RAND_876[63:0];
  _RAND_877 = {2{`RANDOM}};
  record_olddata_109 = _RAND_877[63:0];
  _RAND_878 = {2{`RANDOM}};
  record_olddata_110 = _RAND_878[63:0];
  _RAND_879 = {2{`RANDOM}};
  record_olddata_111 = _RAND_879[63:0];
  _RAND_880 = {2{`RANDOM}};
  record_olddata_112 = _RAND_880[63:0];
  _RAND_881 = {2{`RANDOM}};
  record_olddata_113 = _RAND_881[63:0];
  _RAND_882 = {2{`RANDOM}};
  record_olddata_114 = _RAND_882[63:0];
  _RAND_883 = {2{`RANDOM}};
  record_olddata_115 = _RAND_883[63:0];
  _RAND_884 = {2{`RANDOM}};
  record_olddata_116 = _RAND_884[63:0];
  _RAND_885 = {2{`RANDOM}};
  record_olddata_117 = _RAND_885[63:0];
  _RAND_886 = {2{`RANDOM}};
  record_olddata_118 = _RAND_886[63:0];
  _RAND_887 = {2{`RANDOM}};
  record_olddata_119 = _RAND_887[63:0];
  _RAND_888 = {2{`RANDOM}};
  record_olddata_120 = _RAND_888[63:0];
  _RAND_889 = {2{`RANDOM}};
  record_olddata_121 = _RAND_889[63:0];
  _RAND_890 = {2{`RANDOM}};
  record_olddata_122 = _RAND_890[63:0];
  _RAND_891 = {2{`RANDOM}};
  record_olddata_123 = _RAND_891[63:0];
  _RAND_892 = {2{`RANDOM}};
  record_olddata_124 = _RAND_892[63:0];
  _RAND_893 = {2{`RANDOM}};
  record_olddata_125 = _RAND_893[63:0];
  _RAND_894 = {2{`RANDOM}};
  record_olddata_126 = _RAND_894[63:0];
  _RAND_895 = {2{`RANDOM}};
  record_olddata_127 = _RAND_895[63:0];
  _RAND_896 = {1{`RANDOM}};
  tag_0_0 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  tag_0_1 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  tag_0_2 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  tag_0_3 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  tag_0_4 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  tag_0_5 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  tag_0_6 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  tag_0_7 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  tag_0_8 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  tag_0_9 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  tag_0_10 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  tag_0_11 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  tag_0_12 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  tag_0_13 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  tag_0_14 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  tag_0_15 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  tag_0_16 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  tag_0_17 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  tag_0_18 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  tag_0_19 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  tag_0_20 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  tag_0_21 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  tag_0_22 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  tag_0_23 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  tag_0_24 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  tag_0_25 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  tag_0_26 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  tag_0_27 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  tag_0_28 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  tag_0_29 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  tag_0_30 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  tag_0_31 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  tag_0_32 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  tag_0_33 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  tag_0_34 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  tag_0_35 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  tag_0_36 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  tag_0_37 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  tag_0_38 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  tag_0_39 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  tag_0_40 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  tag_0_41 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  tag_0_42 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  tag_0_43 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  tag_0_44 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  tag_0_45 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  tag_0_46 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  tag_0_47 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  tag_0_48 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  tag_0_49 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  tag_0_50 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  tag_0_51 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  tag_0_52 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  tag_0_53 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  tag_0_54 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  tag_0_55 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  tag_0_56 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  tag_0_57 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  tag_0_58 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  tag_0_59 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  tag_0_60 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  tag_0_61 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  tag_0_62 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  tag_0_63 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  tag_0_64 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  tag_0_65 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  tag_0_66 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  tag_0_67 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  tag_0_68 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  tag_0_69 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  tag_0_70 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  tag_0_71 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  tag_0_72 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  tag_0_73 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  tag_0_74 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  tag_0_75 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  tag_0_76 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  tag_0_77 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  tag_0_78 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  tag_0_79 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  tag_0_80 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  tag_0_81 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  tag_0_82 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  tag_0_83 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  tag_0_84 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  tag_0_85 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  tag_0_86 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  tag_0_87 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  tag_0_88 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  tag_0_89 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  tag_0_90 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  tag_0_91 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  tag_0_92 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  tag_0_93 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  tag_0_94 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  tag_0_95 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  tag_0_96 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  tag_0_97 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  tag_0_98 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  tag_0_99 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  tag_0_100 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  tag_0_101 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  tag_0_102 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  tag_0_103 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  tag_0_104 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  tag_0_105 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  tag_0_106 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  tag_0_107 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  tag_0_108 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  tag_0_109 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  tag_0_110 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  tag_0_111 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  tag_0_112 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  tag_0_113 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  tag_0_114 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  tag_0_115 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  tag_0_116 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  tag_0_117 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  tag_0_118 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  tag_0_119 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  tag_0_120 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  tag_0_121 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  tag_0_122 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  tag_0_123 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  tag_0_124 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  tag_0_125 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  tag_0_126 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  tag_0_127 = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  tag_1_0 = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  tag_1_1 = _RAND_1025[31:0];
  _RAND_1026 = {1{`RANDOM}};
  tag_1_2 = _RAND_1026[31:0];
  _RAND_1027 = {1{`RANDOM}};
  tag_1_3 = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  tag_1_4 = _RAND_1028[31:0];
  _RAND_1029 = {1{`RANDOM}};
  tag_1_5 = _RAND_1029[31:0];
  _RAND_1030 = {1{`RANDOM}};
  tag_1_6 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  tag_1_7 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  tag_1_8 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  tag_1_9 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  tag_1_10 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  tag_1_11 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  tag_1_12 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  tag_1_13 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  tag_1_14 = _RAND_1038[31:0];
  _RAND_1039 = {1{`RANDOM}};
  tag_1_15 = _RAND_1039[31:0];
  _RAND_1040 = {1{`RANDOM}};
  tag_1_16 = _RAND_1040[31:0];
  _RAND_1041 = {1{`RANDOM}};
  tag_1_17 = _RAND_1041[31:0];
  _RAND_1042 = {1{`RANDOM}};
  tag_1_18 = _RAND_1042[31:0];
  _RAND_1043 = {1{`RANDOM}};
  tag_1_19 = _RAND_1043[31:0];
  _RAND_1044 = {1{`RANDOM}};
  tag_1_20 = _RAND_1044[31:0];
  _RAND_1045 = {1{`RANDOM}};
  tag_1_21 = _RAND_1045[31:0];
  _RAND_1046 = {1{`RANDOM}};
  tag_1_22 = _RAND_1046[31:0];
  _RAND_1047 = {1{`RANDOM}};
  tag_1_23 = _RAND_1047[31:0];
  _RAND_1048 = {1{`RANDOM}};
  tag_1_24 = _RAND_1048[31:0];
  _RAND_1049 = {1{`RANDOM}};
  tag_1_25 = _RAND_1049[31:0];
  _RAND_1050 = {1{`RANDOM}};
  tag_1_26 = _RAND_1050[31:0];
  _RAND_1051 = {1{`RANDOM}};
  tag_1_27 = _RAND_1051[31:0];
  _RAND_1052 = {1{`RANDOM}};
  tag_1_28 = _RAND_1052[31:0];
  _RAND_1053 = {1{`RANDOM}};
  tag_1_29 = _RAND_1053[31:0];
  _RAND_1054 = {1{`RANDOM}};
  tag_1_30 = _RAND_1054[31:0];
  _RAND_1055 = {1{`RANDOM}};
  tag_1_31 = _RAND_1055[31:0];
  _RAND_1056 = {1{`RANDOM}};
  tag_1_32 = _RAND_1056[31:0];
  _RAND_1057 = {1{`RANDOM}};
  tag_1_33 = _RAND_1057[31:0];
  _RAND_1058 = {1{`RANDOM}};
  tag_1_34 = _RAND_1058[31:0];
  _RAND_1059 = {1{`RANDOM}};
  tag_1_35 = _RAND_1059[31:0];
  _RAND_1060 = {1{`RANDOM}};
  tag_1_36 = _RAND_1060[31:0];
  _RAND_1061 = {1{`RANDOM}};
  tag_1_37 = _RAND_1061[31:0];
  _RAND_1062 = {1{`RANDOM}};
  tag_1_38 = _RAND_1062[31:0];
  _RAND_1063 = {1{`RANDOM}};
  tag_1_39 = _RAND_1063[31:0];
  _RAND_1064 = {1{`RANDOM}};
  tag_1_40 = _RAND_1064[31:0];
  _RAND_1065 = {1{`RANDOM}};
  tag_1_41 = _RAND_1065[31:0];
  _RAND_1066 = {1{`RANDOM}};
  tag_1_42 = _RAND_1066[31:0];
  _RAND_1067 = {1{`RANDOM}};
  tag_1_43 = _RAND_1067[31:0];
  _RAND_1068 = {1{`RANDOM}};
  tag_1_44 = _RAND_1068[31:0];
  _RAND_1069 = {1{`RANDOM}};
  tag_1_45 = _RAND_1069[31:0];
  _RAND_1070 = {1{`RANDOM}};
  tag_1_46 = _RAND_1070[31:0];
  _RAND_1071 = {1{`RANDOM}};
  tag_1_47 = _RAND_1071[31:0];
  _RAND_1072 = {1{`RANDOM}};
  tag_1_48 = _RAND_1072[31:0];
  _RAND_1073 = {1{`RANDOM}};
  tag_1_49 = _RAND_1073[31:0];
  _RAND_1074 = {1{`RANDOM}};
  tag_1_50 = _RAND_1074[31:0];
  _RAND_1075 = {1{`RANDOM}};
  tag_1_51 = _RAND_1075[31:0];
  _RAND_1076 = {1{`RANDOM}};
  tag_1_52 = _RAND_1076[31:0];
  _RAND_1077 = {1{`RANDOM}};
  tag_1_53 = _RAND_1077[31:0];
  _RAND_1078 = {1{`RANDOM}};
  tag_1_54 = _RAND_1078[31:0];
  _RAND_1079 = {1{`RANDOM}};
  tag_1_55 = _RAND_1079[31:0];
  _RAND_1080 = {1{`RANDOM}};
  tag_1_56 = _RAND_1080[31:0];
  _RAND_1081 = {1{`RANDOM}};
  tag_1_57 = _RAND_1081[31:0];
  _RAND_1082 = {1{`RANDOM}};
  tag_1_58 = _RAND_1082[31:0];
  _RAND_1083 = {1{`RANDOM}};
  tag_1_59 = _RAND_1083[31:0];
  _RAND_1084 = {1{`RANDOM}};
  tag_1_60 = _RAND_1084[31:0];
  _RAND_1085 = {1{`RANDOM}};
  tag_1_61 = _RAND_1085[31:0];
  _RAND_1086 = {1{`RANDOM}};
  tag_1_62 = _RAND_1086[31:0];
  _RAND_1087 = {1{`RANDOM}};
  tag_1_63 = _RAND_1087[31:0];
  _RAND_1088 = {1{`RANDOM}};
  tag_1_64 = _RAND_1088[31:0];
  _RAND_1089 = {1{`RANDOM}};
  tag_1_65 = _RAND_1089[31:0];
  _RAND_1090 = {1{`RANDOM}};
  tag_1_66 = _RAND_1090[31:0];
  _RAND_1091 = {1{`RANDOM}};
  tag_1_67 = _RAND_1091[31:0];
  _RAND_1092 = {1{`RANDOM}};
  tag_1_68 = _RAND_1092[31:0];
  _RAND_1093 = {1{`RANDOM}};
  tag_1_69 = _RAND_1093[31:0];
  _RAND_1094 = {1{`RANDOM}};
  tag_1_70 = _RAND_1094[31:0];
  _RAND_1095 = {1{`RANDOM}};
  tag_1_71 = _RAND_1095[31:0];
  _RAND_1096 = {1{`RANDOM}};
  tag_1_72 = _RAND_1096[31:0];
  _RAND_1097 = {1{`RANDOM}};
  tag_1_73 = _RAND_1097[31:0];
  _RAND_1098 = {1{`RANDOM}};
  tag_1_74 = _RAND_1098[31:0];
  _RAND_1099 = {1{`RANDOM}};
  tag_1_75 = _RAND_1099[31:0];
  _RAND_1100 = {1{`RANDOM}};
  tag_1_76 = _RAND_1100[31:0];
  _RAND_1101 = {1{`RANDOM}};
  tag_1_77 = _RAND_1101[31:0];
  _RAND_1102 = {1{`RANDOM}};
  tag_1_78 = _RAND_1102[31:0];
  _RAND_1103 = {1{`RANDOM}};
  tag_1_79 = _RAND_1103[31:0];
  _RAND_1104 = {1{`RANDOM}};
  tag_1_80 = _RAND_1104[31:0];
  _RAND_1105 = {1{`RANDOM}};
  tag_1_81 = _RAND_1105[31:0];
  _RAND_1106 = {1{`RANDOM}};
  tag_1_82 = _RAND_1106[31:0];
  _RAND_1107 = {1{`RANDOM}};
  tag_1_83 = _RAND_1107[31:0];
  _RAND_1108 = {1{`RANDOM}};
  tag_1_84 = _RAND_1108[31:0];
  _RAND_1109 = {1{`RANDOM}};
  tag_1_85 = _RAND_1109[31:0];
  _RAND_1110 = {1{`RANDOM}};
  tag_1_86 = _RAND_1110[31:0];
  _RAND_1111 = {1{`RANDOM}};
  tag_1_87 = _RAND_1111[31:0];
  _RAND_1112 = {1{`RANDOM}};
  tag_1_88 = _RAND_1112[31:0];
  _RAND_1113 = {1{`RANDOM}};
  tag_1_89 = _RAND_1113[31:0];
  _RAND_1114 = {1{`RANDOM}};
  tag_1_90 = _RAND_1114[31:0];
  _RAND_1115 = {1{`RANDOM}};
  tag_1_91 = _RAND_1115[31:0];
  _RAND_1116 = {1{`RANDOM}};
  tag_1_92 = _RAND_1116[31:0];
  _RAND_1117 = {1{`RANDOM}};
  tag_1_93 = _RAND_1117[31:0];
  _RAND_1118 = {1{`RANDOM}};
  tag_1_94 = _RAND_1118[31:0];
  _RAND_1119 = {1{`RANDOM}};
  tag_1_95 = _RAND_1119[31:0];
  _RAND_1120 = {1{`RANDOM}};
  tag_1_96 = _RAND_1120[31:0];
  _RAND_1121 = {1{`RANDOM}};
  tag_1_97 = _RAND_1121[31:0];
  _RAND_1122 = {1{`RANDOM}};
  tag_1_98 = _RAND_1122[31:0];
  _RAND_1123 = {1{`RANDOM}};
  tag_1_99 = _RAND_1123[31:0];
  _RAND_1124 = {1{`RANDOM}};
  tag_1_100 = _RAND_1124[31:0];
  _RAND_1125 = {1{`RANDOM}};
  tag_1_101 = _RAND_1125[31:0];
  _RAND_1126 = {1{`RANDOM}};
  tag_1_102 = _RAND_1126[31:0];
  _RAND_1127 = {1{`RANDOM}};
  tag_1_103 = _RAND_1127[31:0];
  _RAND_1128 = {1{`RANDOM}};
  tag_1_104 = _RAND_1128[31:0];
  _RAND_1129 = {1{`RANDOM}};
  tag_1_105 = _RAND_1129[31:0];
  _RAND_1130 = {1{`RANDOM}};
  tag_1_106 = _RAND_1130[31:0];
  _RAND_1131 = {1{`RANDOM}};
  tag_1_107 = _RAND_1131[31:0];
  _RAND_1132 = {1{`RANDOM}};
  tag_1_108 = _RAND_1132[31:0];
  _RAND_1133 = {1{`RANDOM}};
  tag_1_109 = _RAND_1133[31:0];
  _RAND_1134 = {1{`RANDOM}};
  tag_1_110 = _RAND_1134[31:0];
  _RAND_1135 = {1{`RANDOM}};
  tag_1_111 = _RAND_1135[31:0];
  _RAND_1136 = {1{`RANDOM}};
  tag_1_112 = _RAND_1136[31:0];
  _RAND_1137 = {1{`RANDOM}};
  tag_1_113 = _RAND_1137[31:0];
  _RAND_1138 = {1{`RANDOM}};
  tag_1_114 = _RAND_1138[31:0];
  _RAND_1139 = {1{`RANDOM}};
  tag_1_115 = _RAND_1139[31:0];
  _RAND_1140 = {1{`RANDOM}};
  tag_1_116 = _RAND_1140[31:0];
  _RAND_1141 = {1{`RANDOM}};
  tag_1_117 = _RAND_1141[31:0];
  _RAND_1142 = {1{`RANDOM}};
  tag_1_118 = _RAND_1142[31:0];
  _RAND_1143 = {1{`RANDOM}};
  tag_1_119 = _RAND_1143[31:0];
  _RAND_1144 = {1{`RANDOM}};
  tag_1_120 = _RAND_1144[31:0];
  _RAND_1145 = {1{`RANDOM}};
  tag_1_121 = _RAND_1145[31:0];
  _RAND_1146 = {1{`RANDOM}};
  tag_1_122 = _RAND_1146[31:0];
  _RAND_1147 = {1{`RANDOM}};
  tag_1_123 = _RAND_1147[31:0];
  _RAND_1148 = {1{`RANDOM}};
  tag_1_124 = _RAND_1148[31:0];
  _RAND_1149 = {1{`RANDOM}};
  tag_1_125 = _RAND_1149[31:0];
  _RAND_1150 = {1{`RANDOM}};
  tag_1_126 = _RAND_1150[31:0];
  _RAND_1151 = {1{`RANDOM}};
  tag_1_127 = _RAND_1151[31:0];
  _RAND_1152 = {1{`RANDOM}};
  valid_0_0 = _RAND_1152[0:0];
  _RAND_1153 = {1{`RANDOM}};
  valid_0_1 = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  valid_0_2 = _RAND_1154[0:0];
  _RAND_1155 = {1{`RANDOM}};
  valid_0_3 = _RAND_1155[0:0];
  _RAND_1156 = {1{`RANDOM}};
  valid_0_4 = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  valid_0_5 = _RAND_1157[0:0];
  _RAND_1158 = {1{`RANDOM}};
  valid_0_6 = _RAND_1158[0:0];
  _RAND_1159 = {1{`RANDOM}};
  valid_0_7 = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  valid_0_8 = _RAND_1160[0:0];
  _RAND_1161 = {1{`RANDOM}};
  valid_0_9 = _RAND_1161[0:0];
  _RAND_1162 = {1{`RANDOM}};
  valid_0_10 = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  valid_0_11 = _RAND_1163[0:0];
  _RAND_1164 = {1{`RANDOM}};
  valid_0_12 = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  valid_0_13 = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  valid_0_14 = _RAND_1166[0:0];
  _RAND_1167 = {1{`RANDOM}};
  valid_0_15 = _RAND_1167[0:0];
  _RAND_1168 = {1{`RANDOM}};
  valid_0_16 = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  valid_0_17 = _RAND_1169[0:0];
  _RAND_1170 = {1{`RANDOM}};
  valid_0_18 = _RAND_1170[0:0];
  _RAND_1171 = {1{`RANDOM}};
  valid_0_19 = _RAND_1171[0:0];
  _RAND_1172 = {1{`RANDOM}};
  valid_0_20 = _RAND_1172[0:0];
  _RAND_1173 = {1{`RANDOM}};
  valid_0_21 = _RAND_1173[0:0];
  _RAND_1174 = {1{`RANDOM}};
  valid_0_22 = _RAND_1174[0:0];
  _RAND_1175 = {1{`RANDOM}};
  valid_0_23 = _RAND_1175[0:0];
  _RAND_1176 = {1{`RANDOM}};
  valid_0_24 = _RAND_1176[0:0];
  _RAND_1177 = {1{`RANDOM}};
  valid_0_25 = _RAND_1177[0:0];
  _RAND_1178 = {1{`RANDOM}};
  valid_0_26 = _RAND_1178[0:0];
  _RAND_1179 = {1{`RANDOM}};
  valid_0_27 = _RAND_1179[0:0];
  _RAND_1180 = {1{`RANDOM}};
  valid_0_28 = _RAND_1180[0:0];
  _RAND_1181 = {1{`RANDOM}};
  valid_0_29 = _RAND_1181[0:0];
  _RAND_1182 = {1{`RANDOM}};
  valid_0_30 = _RAND_1182[0:0];
  _RAND_1183 = {1{`RANDOM}};
  valid_0_31 = _RAND_1183[0:0];
  _RAND_1184 = {1{`RANDOM}};
  valid_0_32 = _RAND_1184[0:0];
  _RAND_1185 = {1{`RANDOM}};
  valid_0_33 = _RAND_1185[0:0];
  _RAND_1186 = {1{`RANDOM}};
  valid_0_34 = _RAND_1186[0:0];
  _RAND_1187 = {1{`RANDOM}};
  valid_0_35 = _RAND_1187[0:0];
  _RAND_1188 = {1{`RANDOM}};
  valid_0_36 = _RAND_1188[0:0];
  _RAND_1189 = {1{`RANDOM}};
  valid_0_37 = _RAND_1189[0:0];
  _RAND_1190 = {1{`RANDOM}};
  valid_0_38 = _RAND_1190[0:0];
  _RAND_1191 = {1{`RANDOM}};
  valid_0_39 = _RAND_1191[0:0];
  _RAND_1192 = {1{`RANDOM}};
  valid_0_40 = _RAND_1192[0:0];
  _RAND_1193 = {1{`RANDOM}};
  valid_0_41 = _RAND_1193[0:0];
  _RAND_1194 = {1{`RANDOM}};
  valid_0_42 = _RAND_1194[0:0];
  _RAND_1195 = {1{`RANDOM}};
  valid_0_43 = _RAND_1195[0:0];
  _RAND_1196 = {1{`RANDOM}};
  valid_0_44 = _RAND_1196[0:0];
  _RAND_1197 = {1{`RANDOM}};
  valid_0_45 = _RAND_1197[0:0];
  _RAND_1198 = {1{`RANDOM}};
  valid_0_46 = _RAND_1198[0:0];
  _RAND_1199 = {1{`RANDOM}};
  valid_0_47 = _RAND_1199[0:0];
  _RAND_1200 = {1{`RANDOM}};
  valid_0_48 = _RAND_1200[0:0];
  _RAND_1201 = {1{`RANDOM}};
  valid_0_49 = _RAND_1201[0:0];
  _RAND_1202 = {1{`RANDOM}};
  valid_0_50 = _RAND_1202[0:0];
  _RAND_1203 = {1{`RANDOM}};
  valid_0_51 = _RAND_1203[0:0];
  _RAND_1204 = {1{`RANDOM}};
  valid_0_52 = _RAND_1204[0:0];
  _RAND_1205 = {1{`RANDOM}};
  valid_0_53 = _RAND_1205[0:0];
  _RAND_1206 = {1{`RANDOM}};
  valid_0_54 = _RAND_1206[0:0];
  _RAND_1207 = {1{`RANDOM}};
  valid_0_55 = _RAND_1207[0:0];
  _RAND_1208 = {1{`RANDOM}};
  valid_0_56 = _RAND_1208[0:0];
  _RAND_1209 = {1{`RANDOM}};
  valid_0_57 = _RAND_1209[0:0];
  _RAND_1210 = {1{`RANDOM}};
  valid_0_58 = _RAND_1210[0:0];
  _RAND_1211 = {1{`RANDOM}};
  valid_0_59 = _RAND_1211[0:0];
  _RAND_1212 = {1{`RANDOM}};
  valid_0_60 = _RAND_1212[0:0];
  _RAND_1213 = {1{`RANDOM}};
  valid_0_61 = _RAND_1213[0:0];
  _RAND_1214 = {1{`RANDOM}};
  valid_0_62 = _RAND_1214[0:0];
  _RAND_1215 = {1{`RANDOM}};
  valid_0_63 = _RAND_1215[0:0];
  _RAND_1216 = {1{`RANDOM}};
  valid_0_64 = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  valid_0_65 = _RAND_1217[0:0];
  _RAND_1218 = {1{`RANDOM}};
  valid_0_66 = _RAND_1218[0:0];
  _RAND_1219 = {1{`RANDOM}};
  valid_0_67 = _RAND_1219[0:0];
  _RAND_1220 = {1{`RANDOM}};
  valid_0_68 = _RAND_1220[0:0];
  _RAND_1221 = {1{`RANDOM}};
  valid_0_69 = _RAND_1221[0:0];
  _RAND_1222 = {1{`RANDOM}};
  valid_0_70 = _RAND_1222[0:0];
  _RAND_1223 = {1{`RANDOM}};
  valid_0_71 = _RAND_1223[0:0];
  _RAND_1224 = {1{`RANDOM}};
  valid_0_72 = _RAND_1224[0:0];
  _RAND_1225 = {1{`RANDOM}};
  valid_0_73 = _RAND_1225[0:0];
  _RAND_1226 = {1{`RANDOM}};
  valid_0_74 = _RAND_1226[0:0];
  _RAND_1227 = {1{`RANDOM}};
  valid_0_75 = _RAND_1227[0:0];
  _RAND_1228 = {1{`RANDOM}};
  valid_0_76 = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  valid_0_77 = _RAND_1229[0:0];
  _RAND_1230 = {1{`RANDOM}};
  valid_0_78 = _RAND_1230[0:0];
  _RAND_1231 = {1{`RANDOM}};
  valid_0_79 = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  valid_0_80 = _RAND_1232[0:0];
  _RAND_1233 = {1{`RANDOM}};
  valid_0_81 = _RAND_1233[0:0];
  _RAND_1234 = {1{`RANDOM}};
  valid_0_82 = _RAND_1234[0:0];
  _RAND_1235 = {1{`RANDOM}};
  valid_0_83 = _RAND_1235[0:0];
  _RAND_1236 = {1{`RANDOM}};
  valid_0_84 = _RAND_1236[0:0];
  _RAND_1237 = {1{`RANDOM}};
  valid_0_85 = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  valid_0_86 = _RAND_1238[0:0];
  _RAND_1239 = {1{`RANDOM}};
  valid_0_87 = _RAND_1239[0:0];
  _RAND_1240 = {1{`RANDOM}};
  valid_0_88 = _RAND_1240[0:0];
  _RAND_1241 = {1{`RANDOM}};
  valid_0_89 = _RAND_1241[0:0];
  _RAND_1242 = {1{`RANDOM}};
  valid_0_90 = _RAND_1242[0:0];
  _RAND_1243 = {1{`RANDOM}};
  valid_0_91 = _RAND_1243[0:0];
  _RAND_1244 = {1{`RANDOM}};
  valid_0_92 = _RAND_1244[0:0];
  _RAND_1245 = {1{`RANDOM}};
  valid_0_93 = _RAND_1245[0:0];
  _RAND_1246 = {1{`RANDOM}};
  valid_0_94 = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  valid_0_95 = _RAND_1247[0:0];
  _RAND_1248 = {1{`RANDOM}};
  valid_0_96 = _RAND_1248[0:0];
  _RAND_1249 = {1{`RANDOM}};
  valid_0_97 = _RAND_1249[0:0];
  _RAND_1250 = {1{`RANDOM}};
  valid_0_98 = _RAND_1250[0:0];
  _RAND_1251 = {1{`RANDOM}};
  valid_0_99 = _RAND_1251[0:0];
  _RAND_1252 = {1{`RANDOM}};
  valid_0_100 = _RAND_1252[0:0];
  _RAND_1253 = {1{`RANDOM}};
  valid_0_101 = _RAND_1253[0:0];
  _RAND_1254 = {1{`RANDOM}};
  valid_0_102 = _RAND_1254[0:0];
  _RAND_1255 = {1{`RANDOM}};
  valid_0_103 = _RAND_1255[0:0];
  _RAND_1256 = {1{`RANDOM}};
  valid_0_104 = _RAND_1256[0:0];
  _RAND_1257 = {1{`RANDOM}};
  valid_0_105 = _RAND_1257[0:0];
  _RAND_1258 = {1{`RANDOM}};
  valid_0_106 = _RAND_1258[0:0];
  _RAND_1259 = {1{`RANDOM}};
  valid_0_107 = _RAND_1259[0:0];
  _RAND_1260 = {1{`RANDOM}};
  valid_0_108 = _RAND_1260[0:0];
  _RAND_1261 = {1{`RANDOM}};
  valid_0_109 = _RAND_1261[0:0];
  _RAND_1262 = {1{`RANDOM}};
  valid_0_110 = _RAND_1262[0:0];
  _RAND_1263 = {1{`RANDOM}};
  valid_0_111 = _RAND_1263[0:0];
  _RAND_1264 = {1{`RANDOM}};
  valid_0_112 = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  valid_0_113 = _RAND_1265[0:0];
  _RAND_1266 = {1{`RANDOM}};
  valid_0_114 = _RAND_1266[0:0];
  _RAND_1267 = {1{`RANDOM}};
  valid_0_115 = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  valid_0_116 = _RAND_1268[0:0];
  _RAND_1269 = {1{`RANDOM}};
  valid_0_117 = _RAND_1269[0:0];
  _RAND_1270 = {1{`RANDOM}};
  valid_0_118 = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  valid_0_119 = _RAND_1271[0:0];
  _RAND_1272 = {1{`RANDOM}};
  valid_0_120 = _RAND_1272[0:0];
  _RAND_1273 = {1{`RANDOM}};
  valid_0_121 = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  valid_0_122 = _RAND_1274[0:0];
  _RAND_1275 = {1{`RANDOM}};
  valid_0_123 = _RAND_1275[0:0];
  _RAND_1276 = {1{`RANDOM}};
  valid_0_124 = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  valid_0_125 = _RAND_1277[0:0];
  _RAND_1278 = {1{`RANDOM}};
  valid_0_126 = _RAND_1278[0:0];
  _RAND_1279 = {1{`RANDOM}};
  valid_0_127 = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  valid_1_0 = _RAND_1280[0:0];
  _RAND_1281 = {1{`RANDOM}};
  valid_1_1 = _RAND_1281[0:0];
  _RAND_1282 = {1{`RANDOM}};
  valid_1_2 = _RAND_1282[0:0];
  _RAND_1283 = {1{`RANDOM}};
  valid_1_3 = _RAND_1283[0:0];
  _RAND_1284 = {1{`RANDOM}};
  valid_1_4 = _RAND_1284[0:0];
  _RAND_1285 = {1{`RANDOM}};
  valid_1_5 = _RAND_1285[0:0];
  _RAND_1286 = {1{`RANDOM}};
  valid_1_6 = _RAND_1286[0:0];
  _RAND_1287 = {1{`RANDOM}};
  valid_1_7 = _RAND_1287[0:0];
  _RAND_1288 = {1{`RANDOM}};
  valid_1_8 = _RAND_1288[0:0];
  _RAND_1289 = {1{`RANDOM}};
  valid_1_9 = _RAND_1289[0:0];
  _RAND_1290 = {1{`RANDOM}};
  valid_1_10 = _RAND_1290[0:0];
  _RAND_1291 = {1{`RANDOM}};
  valid_1_11 = _RAND_1291[0:0];
  _RAND_1292 = {1{`RANDOM}};
  valid_1_12 = _RAND_1292[0:0];
  _RAND_1293 = {1{`RANDOM}};
  valid_1_13 = _RAND_1293[0:0];
  _RAND_1294 = {1{`RANDOM}};
  valid_1_14 = _RAND_1294[0:0];
  _RAND_1295 = {1{`RANDOM}};
  valid_1_15 = _RAND_1295[0:0];
  _RAND_1296 = {1{`RANDOM}};
  valid_1_16 = _RAND_1296[0:0];
  _RAND_1297 = {1{`RANDOM}};
  valid_1_17 = _RAND_1297[0:0];
  _RAND_1298 = {1{`RANDOM}};
  valid_1_18 = _RAND_1298[0:0];
  _RAND_1299 = {1{`RANDOM}};
  valid_1_19 = _RAND_1299[0:0];
  _RAND_1300 = {1{`RANDOM}};
  valid_1_20 = _RAND_1300[0:0];
  _RAND_1301 = {1{`RANDOM}};
  valid_1_21 = _RAND_1301[0:0];
  _RAND_1302 = {1{`RANDOM}};
  valid_1_22 = _RAND_1302[0:0];
  _RAND_1303 = {1{`RANDOM}};
  valid_1_23 = _RAND_1303[0:0];
  _RAND_1304 = {1{`RANDOM}};
  valid_1_24 = _RAND_1304[0:0];
  _RAND_1305 = {1{`RANDOM}};
  valid_1_25 = _RAND_1305[0:0];
  _RAND_1306 = {1{`RANDOM}};
  valid_1_26 = _RAND_1306[0:0];
  _RAND_1307 = {1{`RANDOM}};
  valid_1_27 = _RAND_1307[0:0];
  _RAND_1308 = {1{`RANDOM}};
  valid_1_28 = _RAND_1308[0:0];
  _RAND_1309 = {1{`RANDOM}};
  valid_1_29 = _RAND_1309[0:0];
  _RAND_1310 = {1{`RANDOM}};
  valid_1_30 = _RAND_1310[0:0];
  _RAND_1311 = {1{`RANDOM}};
  valid_1_31 = _RAND_1311[0:0];
  _RAND_1312 = {1{`RANDOM}};
  valid_1_32 = _RAND_1312[0:0];
  _RAND_1313 = {1{`RANDOM}};
  valid_1_33 = _RAND_1313[0:0];
  _RAND_1314 = {1{`RANDOM}};
  valid_1_34 = _RAND_1314[0:0];
  _RAND_1315 = {1{`RANDOM}};
  valid_1_35 = _RAND_1315[0:0];
  _RAND_1316 = {1{`RANDOM}};
  valid_1_36 = _RAND_1316[0:0];
  _RAND_1317 = {1{`RANDOM}};
  valid_1_37 = _RAND_1317[0:0];
  _RAND_1318 = {1{`RANDOM}};
  valid_1_38 = _RAND_1318[0:0];
  _RAND_1319 = {1{`RANDOM}};
  valid_1_39 = _RAND_1319[0:0];
  _RAND_1320 = {1{`RANDOM}};
  valid_1_40 = _RAND_1320[0:0];
  _RAND_1321 = {1{`RANDOM}};
  valid_1_41 = _RAND_1321[0:0];
  _RAND_1322 = {1{`RANDOM}};
  valid_1_42 = _RAND_1322[0:0];
  _RAND_1323 = {1{`RANDOM}};
  valid_1_43 = _RAND_1323[0:0];
  _RAND_1324 = {1{`RANDOM}};
  valid_1_44 = _RAND_1324[0:0];
  _RAND_1325 = {1{`RANDOM}};
  valid_1_45 = _RAND_1325[0:0];
  _RAND_1326 = {1{`RANDOM}};
  valid_1_46 = _RAND_1326[0:0];
  _RAND_1327 = {1{`RANDOM}};
  valid_1_47 = _RAND_1327[0:0];
  _RAND_1328 = {1{`RANDOM}};
  valid_1_48 = _RAND_1328[0:0];
  _RAND_1329 = {1{`RANDOM}};
  valid_1_49 = _RAND_1329[0:0];
  _RAND_1330 = {1{`RANDOM}};
  valid_1_50 = _RAND_1330[0:0];
  _RAND_1331 = {1{`RANDOM}};
  valid_1_51 = _RAND_1331[0:0];
  _RAND_1332 = {1{`RANDOM}};
  valid_1_52 = _RAND_1332[0:0];
  _RAND_1333 = {1{`RANDOM}};
  valid_1_53 = _RAND_1333[0:0];
  _RAND_1334 = {1{`RANDOM}};
  valid_1_54 = _RAND_1334[0:0];
  _RAND_1335 = {1{`RANDOM}};
  valid_1_55 = _RAND_1335[0:0];
  _RAND_1336 = {1{`RANDOM}};
  valid_1_56 = _RAND_1336[0:0];
  _RAND_1337 = {1{`RANDOM}};
  valid_1_57 = _RAND_1337[0:0];
  _RAND_1338 = {1{`RANDOM}};
  valid_1_58 = _RAND_1338[0:0];
  _RAND_1339 = {1{`RANDOM}};
  valid_1_59 = _RAND_1339[0:0];
  _RAND_1340 = {1{`RANDOM}};
  valid_1_60 = _RAND_1340[0:0];
  _RAND_1341 = {1{`RANDOM}};
  valid_1_61 = _RAND_1341[0:0];
  _RAND_1342 = {1{`RANDOM}};
  valid_1_62 = _RAND_1342[0:0];
  _RAND_1343 = {1{`RANDOM}};
  valid_1_63 = _RAND_1343[0:0];
  _RAND_1344 = {1{`RANDOM}};
  valid_1_64 = _RAND_1344[0:0];
  _RAND_1345 = {1{`RANDOM}};
  valid_1_65 = _RAND_1345[0:0];
  _RAND_1346 = {1{`RANDOM}};
  valid_1_66 = _RAND_1346[0:0];
  _RAND_1347 = {1{`RANDOM}};
  valid_1_67 = _RAND_1347[0:0];
  _RAND_1348 = {1{`RANDOM}};
  valid_1_68 = _RAND_1348[0:0];
  _RAND_1349 = {1{`RANDOM}};
  valid_1_69 = _RAND_1349[0:0];
  _RAND_1350 = {1{`RANDOM}};
  valid_1_70 = _RAND_1350[0:0];
  _RAND_1351 = {1{`RANDOM}};
  valid_1_71 = _RAND_1351[0:0];
  _RAND_1352 = {1{`RANDOM}};
  valid_1_72 = _RAND_1352[0:0];
  _RAND_1353 = {1{`RANDOM}};
  valid_1_73 = _RAND_1353[0:0];
  _RAND_1354 = {1{`RANDOM}};
  valid_1_74 = _RAND_1354[0:0];
  _RAND_1355 = {1{`RANDOM}};
  valid_1_75 = _RAND_1355[0:0];
  _RAND_1356 = {1{`RANDOM}};
  valid_1_76 = _RAND_1356[0:0];
  _RAND_1357 = {1{`RANDOM}};
  valid_1_77 = _RAND_1357[0:0];
  _RAND_1358 = {1{`RANDOM}};
  valid_1_78 = _RAND_1358[0:0];
  _RAND_1359 = {1{`RANDOM}};
  valid_1_79 = _RAND_1359[0:0];
  _RAND_1360 = {1{`RANDOM}};
  valid_1_80 = _RAND_1360[0:0];
  _RAND_1361 = {1{`RANDOM}};
  valid_1_81 = _RAND_1361[0:0];
  _RAND_1362 = {1{`RANDOM}};
  valid_1_82 = _RAND_1362[0:0];
  _RAND_1363 = {1{`RANDOM}};
  valid_1_83 = _RAND_1363[0:0];
  _RAND_1364 = {1{`RANDOM}};
  valid_1_84 = _RAND_1364[0:0];
  _RAND_1365 = {1{`RANDOM}};
  valid_1_85 = _RAND_1365[0:0];
  _RAND_1366 = {1{`RANDOM}};
  valid_1_86 = _RAND_1366[0:0];
  _RAND_1367 = {1{`RANDOM}};
  valid_1_87 = _RAND_1367[0:0];
  _RAND_1368 = {1{`RANDOM}};
  valid_1_88 = _RAND_1368[0:0];
  _RAND_1369 = {1{`RANDOM}};
  valid_1_89 = _RAND_1369[0:0];
  _RAND_1370 = {1{`RANDOM}};
  valid_1_90 = _RAND_1370[0:0];
  _RAND_1371 = {1{`RANDOM}};
  valid_1_91 = _RAND_1371[0:0];
  _RAND_1372 = {1{`RANDOM}};
  valid_1_92 = _RAND_1372[0:0];
  _RAND_1373 = {1{`RANDOM}};
  valid_1_93 = _RAND_1373[0:0];
  _RAND_1374 = {1{`RANDOM}};
  valid_1_94 = _RAND_1374[0:0];
  _RAND_1375 = {1{`RANDOM}};
  valid_1_95 = _RAND_1375[0:0];
  _RAND_1376 = {1{`RANDOM}};
  valid_1_96 = _RAND_1376[0:0];
  _RAND_1377 = {1{`RANDOM}};
  valid_1_97 = _RAND_1377[0:0];
  _RAND_1378 = {1{`RANDOM}};
  valid_1_98 = _RAND_1378[0:0];
  _RAND_1379 = {1{`RANDOM}};
  valid_1_99 = _RAND_1379[0:0];
  _RAND_1380 = {1{`RANDOM}};
  valid_1_100 = _RAND_1380[0:0];
  _RAND_1381 = {1{`RANDOM}};
  valid_1_101 = _RAND_1381[0:0];
  _RAND_1382 = {1{`RANDOM}};
  valid_1_102 = _RAND_1382[0:0];
  _RAND_1383 = {1{`RANDOM}};
  valid_1_103 = _RAND_1383[0:0];
  _RAND_1384 = {1{`RANDOM}};
  valid_1_104 = _RAND_1384[0:0];
  _RAND_1385 = {1{`RANDOM}};
  valid_1_105 = _RAND_1385[0:0];
  _RAND_1386 = {1{`RANDOM}};
  valid_1_106 = _RAND_1386[0:0];
  _RAND_1387 = {1{`RANDOM}};
  valid_1_107 = _RAND_1387[0:0];
  _RAND_1388 = {1{`RANDOM}};
  valid_1_108 = _RAND_1388[0:0];
  _RAND_1389 = {1{`RANDOM}};
  valid_1_109 = _RAND_1389[0:0];
  _RAND_1390 = {1{`RANDOM}};
  valid_1_110 = _RAND_1390[0:0];
  _RAND_1391 = {1{`RANDOM}};
  valid_1_111 = _RAND_1391[0:0];
  _RAND_1392 = {1{`RANDOM}};
  valid_1_112 = _RAND_1392[0:0];
  _RAND_1393 = {1{`RANDOM}};
  valid_1_113 = _RAND_1393[0:0];
  _RAND_1394 = {1{`RANDOM}};
  valid_1_114 = _RAND_1394[0:0];
  _RAND_1395 = {1{`RANDOM}};
  valid_1_115 = _RAND_1395[0:0];
  _RAND_1396 = {1{`RANDOM}};
  valid_1_116 = _RAND_1396[0:0];
  _RAND_1397 = {1{`RANDOM}};
  valid_1_117 = _RAND_1397[0:0];
  _RAND_1398 = {1{`RANDOM}};
  valid_1_118 = _RAND_1398[0:0];
  _RAND_1399 = {1{`RANDOM}};
  valid_1_119 = _RAND_1399[0:0];
  _RAND_1400 = {1{`RANDOM}};
  valid_1_120 = _RAND_1400[0:0];
  _RAND_1401 = {1{`RANDOM}};
  valid_1_121 = _RAND_1401[0:0];
  _RAND_1402 = {1{`RANDOM}};
  valid_1_122 = _RAND_1402[0:0];
  _RAND_1403 = {1{`RANDOM}};
  valid_1_123 = _RAND_1403[0:0];
  _RAND_1404 = {1{`RANDOM}};
  valid_1_124 = _RAND_1404[0:0];
  _RAND_1405 = {1{`RANDOM}};
  valid_1_125 = _RAND_1405[0:0];
  _RAND_1406 = {1{`RANDOM}};
  valid_1_126 = _RAND_1406[0:0];
  _RAND_1407 = {1{`RANDOM}};
  valid_1_127 = _RAND_1407[0:0];
  _RAND_1408 = {1{`RANDOM}};
  dirty_0_0 = _RAND_1408[0:0];
  _RAND_1409 = {1{`RANDOM}};
  dirty_0_1 = _RAND_1409[0:0];
  _RAND_1410 = {1{`RANDOM}};
  dirty_0_2 = _RAND_1410[0:0];
  _RAND_1411 = {1{`RANDOM}};
  dirty_0_3 = _RAND_1411[0:0];
  _RAND_1412 = {1{`RANDOM}};
  dirty_0_4 = _RAND_1412[0:0];
  _RAND_1413 = {1{`RANDOM}};
  dirty_0_5 = _RAND_1413[0:0];
  _RAND_1414 = {1{`RANDOM}};
  dirty_0_6 = _RAND_1414[0:0];
  _RAND_1415 = {1{`RANDOM}};
  dirty_0_7 = _RAND_1415[0:0];
  _RAND_1416 = {1{`RANDOM}};
  dirty_0_8 = _RAND_1416[0:0];
  _RAND_1417 = {1{`RANDOM}};
  dirty_0_9 = _RAND_1417[0:0];
  _RAND_1418 = {1{`RANDOM}};
  dirty_0_10 = _RAND_1418[0:0];
  _RAND_1419 = {1{`RANDOM}};
  dirty_0_11 = _RAND_1419[0:0];
  _RAND_1420 = {1{`RANDOM}};
  dirty_0_12 = _RAND_1420[0:0];
  _RAND_1421 = {1{`RANDOM}};
  dirty_0_13 = _RAND_1421[0:0];
  _RAND_1422 = {1{`RANDOM}};
  dirty_0_14 = _RAND_1422[0:0];
  _RAND_1423 = {1{`RANDOM}};
  dirty_0_15 = _RAND_1423[0:0];
  _RAND_1424 = {1{`RANDOM}};
  dirty_0_16 = _RAND_1424[0:0];
  _RAND_1425 = {1{`RANDOM}};
  dirty_0_17 = _RAND_1425[0:0];
  _RAND_1426 = {1{`RANDOM}};
  dirty_0_18 = _RAND_1426[0:0];
  _RAND_1427 = {1{`RANDOM}};
  dirty_0_19 = _RAND_1427[0:0];
  _RAND_1428 = {1{`RANDOM}};
  dirty_0_20 = _RAND_1428[0:0];
  _RAND_1429 = {1{`RANDOM}};
  dirty_0_21 = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  dirty_0_22 = _RAND_1430[0:0];
  _RAND_1431 = {1{`RANDOM}};
  dirty_0_23 = _RAND_1431[0:0];
  _RAND_1432 = {1{`RANDOM}};
  dirty_0_24 = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  dirty_0_25 = _RAND_1433[0:0];
  _RAND_1434 = {1{`RANDOM}};
  dirty_0_26 = _RAND_1434[0:0];
  _RAND_1435 = {1{`RANDOM}};
  dirty_0_27 = _RAND_1435[0:0];
  _RAND_1436 = {1{`RANDOM}};
  dirty_0_28 = _RAND_1436[0:0];
  _RAND_1437 = {1{`RANDOM}};
  dirty_0_29 = _RAND_1437[0:0];
  _RAND_1438 = {1{`RANDOM}};
  dirty_0_30 = _RAND_1438[0:0];
  _RAND_1439 = {1{`RANDOM}};
  dirty_0_31 = _RAND_1439[0:0];
  _RAND_1440 = {1{`RANDOM}};
  dirty_0_32 = _RAND_1440[0:0];
  _RAND_1441 = {1{`RANDOM}};
  dirty_0_33 = _RAND_1441[0:0];
  _RAND_1442 = {1{`RANDOM}};
  dirty_0_34 = _RAND_1442[0:0];
  _RAND_1443 = {1{`RANDOM}};
  dirty_0_35 = _RAND_1443[0:0];
  _RAND_1444 = {1{`RANDOM}};
  dirty_0_36 = _RAND_1444[0:0];
  _RAND_1445 = {1{`RANDOM}};
  dirty_0_37 = _RAND_1445[0:0];
  _RAND_1446 = {1{`RANDOM}};
  dirty_0_38 = _RAND_1446[0:0];
  _RAND_1447 = {1{`RANDOM}};
  dirty_0_39 = _RAND_1447[0:0];
  _RAND_1448 = {1{`RANDOM}};
  dirty_0_40 = _RAND_1448[0:0];
  _RAND_1449 = {1{`RANDOM}};
  dirty_0_41 = _RAND_1449[0:0];
  _RAND_1450 = {1{`RANDOM}};
  dirty_0_42 = _RAND_1450[0:0];
  _RAND_1451 = {1{`RANDOM}};
  dirty_0_43 = _RAND_1451[0:0];
  _RAND_1452 = {1{`RANDOM}};
  dirty_0_44 = _RAND_1452[0:0];
  _RAND_1453 = {1{`RANDOM}};
  dirty_0_45 = _RAND_1453[0:0];
  _RAND_1454 = {1{`RANDOM}};
  dirty_0_46 = _RAND_1454[0:0];
  _RAND_1455 = {1{`RANDOM}};
  dirty_0_47 = _RAND_1455[0:0];
  _RAND_1456 = {1{`RANDOM}};
  dirty_0_48 = _RAND_1456[0:0];
  _RAND_1457 = {1{`RANDOM}};
  dirty_0_49 = _RAND_1457[0:0];
  _RAND_1458 = {1{`RANDOM}};
  dirty_0_50 = _RAND_1458[0:0];
  _RAND_1459 = {1{`RANDOM}};
  dirty_0_51 = _RAND_1459[0:0];
  _RAND_1460 = {1{`RANDOM}};
  dirty_0_52 = _RAND_1460[0:0];
  _RAND_1461 = {1{`RANDOM}};
  dirty_0_53 = _RAND_1461[0:0];
  _RAND_1462 = {1{`RANDOM}};
  dirty_0_54 = _RAND_1462[0:0];
  _RAND_1463 = {1{`RANDOM}};
  dirty_0_55 = _RAND_1463[0:0];
  _RAND_1464 = {1{`RANDOM}};
  dirty_0_56 = _RAND_1464[0:0];
  _RAND_1465 = {1{`RANDOM}};
  dirty_0_57 = _RAND_1465[0:0];
  _RAND_1466 = {1{`RANDOM}};
  dirty_0_58 = _RAND_1466[0:0];
  _RAND_1467 = {1{`RANDOM}};
  dirty_0_59 = _RAND_1467[0:0];
  _RAND_1468 = {1{`RANDOM}};
  dirty_0_60 = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  dirty_0_61 = _RAND_1469[0:0];
  _RAND_1470 = {1{`RANDOM}};
  dirty_0_62 = _RAND_1470[0:0];
  _RAND_1471 = {1{`RANDOM}};
  dirty_0_63 = _RAND_1471[0:0];
  _RAND_1472 = {1{`RANDOM}};
  dirty_0_64 = _RAND_1472[0:0];
  _RAND_1473 = {1{`RANDOM}};
  dirty_0_65 = _RAND_1473[0:0];
  _RAND_1474 = {1{`RANDOM}};
  dirty_0_66 = _RAND_1474[0:0];
  _RAND_1475 = {1{`RANDOM}};
  dirty_0_67 = _RAND_1475[0:0];
  _RAND_1476 = {1{`RANDOM}};
  dirty_0_68 = _RAND_1476[0:0];
  _RAND_1477 = {1{`RANDOM}};
  dirty_0_69 = _RAND_1477[0:0];
  _RAND_1478 = {1{`RANDOM}};
  dirty_0_70 = _RAND_1478[0:0];
  _RAND_1479 = {1{`RANDOM}};
  dirty_0_71 = _RAND_1479[0:0];
  _RAND_1480 = {1{`RANDOM}};
  dirty_0_72 = _RAND_1480[0:0];
  _RAND_1481 = {1{`RANDOM}};
  dirty_0_73 = _RAND_1481[0:0];
  _RAND_1482 = {1{`RANDOM}};
  dirty_0_74 = _RAND_1482[0:0];
  _RAND_1483 = {1{`RANDOM}};
  dirty_0_75 = _RAND_1483[0:0];
  _RAND_1484 = {1{`RANDOM}};
  dirty_0_76 = _RAND_1484[0:0];
  _RAND_1485 = {1{`RANDOM}};
  dirty_0_77 = _RAND_1485[0:0];
  _RAND_1486 = {1{`RANDOM}};
  dirty_0_78 = _RAND_1486[0:0];
  _RAND_1487 = {1{`RANDOM}};
  dirty_0_79 = _RAND_1487[0:0];
  _RAND_1488 = {1{`RANDOM}};
  dirty_0_80 = _RAND_1488[0:0];
  _RAND_1489 = {1{`RANDOM}};
  dirty_0_81 = _RAND_1489[0:0];
  _RAND_1490 = {1{`RANDOM}};
  dirty_0_82 = _RAND_1490[0:0];
  _RAND_1491 = {1{`RANDOM}};
  dirty_0_83 = _RAND_1491[0:0];
  _RAND_1492 = {1{`RANDOM}};
  dirty_0_84 = _RAND_1492[0:0];
  _RAND_1493 = {1{`RANDOM}};
  dirty_0_85 = _RAND_1493[0:0];
  _RAND_1494 = {1{`RANDOM}};
  dirty_0_86 = _RAND_1494[0:0];
  _RAND_1495 = {1{`RANDOM}};
  dirty_0_87 = _RAND_1495[0:0];
  _RAND_1496 = {1{`RANDOM}};
  dirty_0_88 = _RAND_1496[0:0];
  _RAND_1497 = {1{`RANDOM}};
  dirty_0_89 = _RAND_1497[0:0];
  _RAND_1498 = {1{`RANDOM}};
  dirty_0_90 = _RAND_1498[0:0];
  _RAND_1499 = {1{`RANDOM}};
  dirty_0_91 = _RAND_1499[0:0];
  _RAND_1500 = {1{`RANDOM}};
  dirty_0_92 = _RAND_1500[0:0];
  _RAND_1501 = {1{`RANDOM}};
  dirty_0_93 = _RAND_1501[0:0];
  _RAND_1502 = {1{`RANDOM}};
  dirty_0_94 = _RAND_1502[0:0];
  _RAND_1503 = {1{`RANDOM}};
  dirty_0_95 = _RAND_1503[0:0];
  _RAND_1504 = {1{`RANDOM}};
  dirty_0_96 = _RAND_1504[0:0];
  _RAND_1505 = {1{`RANDOM}};
  dirty_0_97 = _RAND_1505[0:0];
  _RAND_1506 = {1{`RANDOM}};
  dirty_0_98 = _RAND_1506[0:0];
  _RAND_1507 = {1{`RANDOM}};
  dirty_0_99 = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  dirty_0_100 = _RAND_1508[0:0];
  _RAND_1509 = {1{`RANDOM}};
  dirty_0_101 = _RAND_1509[0:0];
  _RAND_1510 = {1{`RANDOM}};
  dirty_0_102 = _RAND_1510[0:0];
  _RAND_1511 = {1{`RANDOM}};
  dirty_0_103 = _RAND_1511[0:0];
  _RAND_1512 = {1{`RANDOM}};
  dirty_0_104 = _RAND_1512[0:0];
  _RAND_1513 = {1{`RANDOM}};
  dirty_0_105 = _RAND_1513[0:0];
  _RAND_1514 = {1{`RANDOM}};
  dirty_0_106 = _RAND_1514[0:0];
  _RAND_1515 = {1{`RANDOM}};
  dirty_0_107 = _RAND_1515[0:0];
  _RAND_1516 = {1{`RANDOM}};
  dirty_0_108 = _RAND_1516[0:0];
  _RAND_1517 = {1{`RANDOM}};
  dirty_0_109 = _RAND_1517[0:0];
  _RAND_1518 = {1{`RANDOM}};
  dirty_0_110 = _RAND_1518[0:0];
  _RAND_1519 = {1{`RANDOM}};
  dirty_0_111 = _RAND_1519[0:0];
  _RAND_1520 = {1{`RANDOM}};
  dirty_0_112 = _RAND_1520[0:0];
  _RAND_1521 = {1{`RANDOM}};
  dirty_0_113 = _RAND_1521[0:0];
  _RAND_1522 = {1{`RANDOM}};
  dirty_0_114 = _RAND_1522[0:0];
  _RAND_1523 = {1{`RANDOM}};
  dirty_0_115 = _RAND_1523[0:0];
  _RAND_1524 = {1{`RANDOM}};
  dirty_0_116 = _RAND_1524[0:0];
  _RAND_1525 = {1{`RANDOM}};
  dirty_0_117 = _RAND_1525[0:0];
  _RAND_1526 = {1{`RANDOM}};
  dirty_0_118 = _RAND_1526[0:0];
  _RAND_1527 = {1{`RANDOM}};
  dirty_0_119 = _RAND_1527[0:0];
  _RAND_1528 = {1{`RANDOM}};
  dirty_0_120 = _RAND_1528[0:0];
  _RAND_1529 = {1{`RANDOM}};
  dirty_0_121 = _RAND_1529[0:0];
  _RAND_1530 = {1{`RANDOM}};
  dirty_0_122 = _RAND_1530[0:0];
  _RAND_1531 = {1{`RANDOM}};
  dirty_0_123 = _RAND_1531[0:0];
  _RAND_1532 = {1{`RANDOM}};
  dirty_0_124 = _RAND_1532[0:0];
  _RAND_1533 = {1{`RANDOM}};
  dirty_0_125 = _RAND_1533[0:0];
  _RAND_1534 = {1{`RANDOM}};
  dirty_0_126 = _RAND_1534[0:0];
  _RAND_1535 = {1{`RANDOM}};
  dirty_0_127 = _RAND_1535[0:0];
  _RAND_1536 = {1{`RANDOM}};
  dirty_1_0 = _RAND_1536[0:0];
  _RAND_1537 = {1{`RANDOM}};
  dirty_1_1 = _RAND_1537[0:0];
  _RAND_1538 = {1{`RANDOM}};
  dirty_1_2 = _RAND_1538[0:0];
  _RAND_1539 = {1{`RANDOM}};
  dirty_1_3 = _RAND_1539[0:0];
  _RAND_1540 = {1{`RANDOM}};
  dirty_1_4 = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  dirty_1_5 = _RAND_1541[0:0];
  _RAND_1542 = {1{`RANDOM}};
  dirty_1_6 = _RAND_1542[0:0];
  _RAND_1543 = {1{`RANDOM}};
  dirty_1_7 = _RAND_1543[0:0];
  _RAND_1544 = {1{`RANDOM}};
  dirty_1_8 = _RAND_1544[0:0];
  _RAND_1545 = {1{`RANDOM}};
  dirty_1_9 = _RAND_1545[0:0];
  _RAND_1546 = {1{`RANDOM}};
  dirty_1_10 = _RAND_1546[0:0];
  _RAND_1547 = {1{`RANDOM}};
  dirty_1_11 = _RAND_1547[0:0];
  _RAND_1548 = {1{`RANDOM}};
  dirty_1_12 = _RAND_1548[0:0];
  _RAND_1549 = {1{`RANDOM}};
  dirty_1_13 = _RAND_1549[0:0];
  _RAND_1550 = {1{`RANDOM}};
  dirty_1_14 = _RAND_1550[0:0];
  _RAND_1551 = {1{`RANDOM}};
  dirty_1_15 = _RAND_1551[0:0];
  _RAND_1552 = {1{`RANDOM}};
  dirty_1_16 = _RAND_1552[0:0];
  _RAND_1553 = {1{`RANDOM}};
  dirty_1_17 = _RAND_1553[0:0];
  _RAND_1554 = {1{`RANDOM}};
  dirty_1_18 = _RAND_1554[0:0];
  _RAND_1555 = {1{`RANDOM}};
  dirty_1_19 = _RAND_1555[0:0];
  _RAND_1556 = {1{`RANDOM}};
  dirty_1_20 = _RAND_1556[0:0];
  _RAND_1557 = {1{`RANDOM}};
  dirty_1_21 = _RAND_1557[0:0];
  _RAND_1558 = {1{`RANDOM}};
  dirty_1_22 = _RAND_1558[0:0];
  _RAND_1559 = {1{`RANDOM}};
  dirty_1_23 = _RAND_1559[0:0];
  _RAND_1560 = {1{`RANDOM}};
  dirty_1_24 = _RAND_1560[0:0];
  _RAND_1561 = {1{`RANDOM}};
  dirty_1_25 = _RAND_1561[0:0];
  _RAND_1562 = {1{`RANDOM}};
  dirty_1_26 = _RAND_1562[0:0];
  _RAND_1563 = {1{`RANDOM}};
  dirty_1_27 = _RAND_1563[0:0];
  _RAND_1564 = {1{`RANDOM}};
  dirty_1_28 = _RAND_1564[0:0];
  _RAND_1565 = {1{`RANDOM}};
  dirty_1_29 = _RAND_1565[0:0];
  _RAND_1566 = {1{`RANDOM}};
  dirty_1_30 = _RAND_1566[0:0];
  _RAND_1567 = {1{`RANDOM}};
  dirty_1_31 = _RAND_1567[0:0];
  _RAND_1568 = {1{`RANDOM}};
  dirty_1_32 = _RAND_1568[0:0];
  _RAND_1569 = {1{`RANDOM}};
  dirty_1_33 = _RAND_1569[0:0];
  _RAND_1570 = {1{`RANDOM}};
  dirty_1_34 = _RAND_1570[0:0];
  _RAND_1571 = {1{`RANDOM}};
  dirty_1_35 = _RAND_1571[0:0];
  _RAND_1572 = {1{`RANDOM}};
  dirty_1_36 = _RAND_1572[0:0];
  _RAND_1573 = {1{`RANDOM}};
  dirty_1_37 = _RAND_1573[0:0];
  _RAND_1574 = {1{`RANDOM}};
  dirty_1_38 = _RAND_1574[0:0];
  _RAND_1575 = {1{`RANDOM}};
  dirty_1_39 = _RAND_1575[0:0];
  _RAND_1576 = {1{`RANDOM}};
  dirty_1_40 = _RAND_1576[0:0];
  _RAND_1577 = {1{`RANDOM}};
  dirty_1_41 = _RAND_1577[0:0];
  _RAND_1578 = {1{`RANDOM}};
  dirty_1_42 = _RAND_1578[0:0];
  _RAND_1579 = {1{`RANDOM}};
  dirty_1_43 = _RAND_1579[0:0];
  _RAND_1580 = {1{`RANDOM}};
  dirty_1_44 = _RAND_1580[0:0];
  _RAND_1581 = {1{`RANDOM}};
  dirty_1_45 = _RAND_1581[0:0];
  _RAND_1582 = {1{`RANDOM}};
  dirty_1_46 = _RAND_1582[0:0];
  _RAND_1583 = {1{`RANDOM}};
  dirty_1_47 = _RAND_1583[0:0];
  _RAND_1584 = {1{`RANDOM}};
  dirty_1_48 = _RAND_1584[0:0];
  _RAND_1585 = {1{`RANDOM}};
  dirty_1_49 = _RAND_1585[0:0];
  _RAND_1586 = {1{`RANDOM}};
  dirty_1_50 = _RAND_1586[0:0];
  _RAND_1587 = {1{`RANDOM}};
  dirty_1_51 = _RAND_1587[0:0];
  _RAND_1588 = {1{`RANDOM}};
  dirty_1_52 = _RAND_1588[0:0];
  _RAND_1589 = {1{`RANDOM}};
  dirty_1_53 = _RAND_1589[0:0];
  _RAND_1590 = {1{`RANDOM}};
  dirty_1_54 = _RAND_1590[0:0];
  _RAND_1591 = {1{`RANDOM}};
  dirty_1_55 = _RAND_1591[0:0];
  _RAND_1592 = {1{`RANDOM}};
  dirty_1_56 = _RAND_1592[0:0];
  _RAND_1593 = {1{`RANDOM}};
  dirty_1_57 = _RAND_1593[0:0];
  _RAND_1594 = {1{`RANDOM}};
  dirty_1_58 = _RAND_1594[0:0];
  _RAND_1595 = {1{`RANDOM}};
  dirty_1_59 = _RAND_1595[0:0];
  _RAND_1596 = {1{`RANDOM}};
  dirty_1_60 = _RAND_1596[0:0];
  _RAND_1597 = {1{`RANDOM}};
  dirty_1_61 = _RAND_1597[0:0];
  _RAND_1598 = {1{`RANDOM}};
  dirty_1_62 = _RAND_1598[0:0];
  _RAND_1599 = {1{`RANDOM}};
  dirty_1_63 = _RAND_1599[0:0];
  _RAND_1600 = {1{`RANDOM}};
  dirty_1_64 = _RAND_1600[0:0];
  _RAND_1601 = {1{`RANDOM}};
  dirty_1_65 = _RAND_1601[0:0];
  _RAND_1602 = {1{`RANDOM}};
  dirty_1_66 = _RAND_1602[0:0];
  _RAND_1603 = {1{`RANDOM}};
  dirty_1_67 = _RAND_1603[0:0];
  _RAND_1604 = {1{`RANDOM}};
  dirty_1_68 = _RAND_1604[0:0];
  _RAND_1605 = {1{`RANDOM}};
  dirty_1_69 = _RAND_1605[0:0];
  _RAND_1606 = {1{`RANDOM}};
  dirty_1_70 = _RAND_1606[0:0];
  _RAND_1607 = {1{`RANDOM}};
  dirty_1_71 = _RAND_1607[0:0];
  _RAND_1608 = {1{`RANDOM}};
  dirty_1_72 = _RAND_1608[0:0];
  _RAND_1609 = {1{`RANDOM}};
  dirty_1_73 = _RAND_1609[0:0];
  _RAND_1610 = {1{`RANDOM}};
  dirty_1_74 = _RAND_1610[0:0];
  _RAND_1611 = {1{`RANDOM}};
  dirty_1_75 = _RAND_1611[0:0];
  _RAND_1612 = {1{`RANDOM}};
  dirty_1_76 = _RAND_1612[0:0];
  _RAND_1613 = {1{`RANDOM}};
  dirty_1_77 = _RAND_1613[0:0];
  _RAND_1614 = {1{`RANDOM}};
  dirty_1_78 = _RAND_1614[0:0];
  _RAND_1615 = {1{`RANDOM}};
  dirty_1_79 = _RAND_1615[0:0];
  _RAND_1616 = {1{`RANDOM}};
  dirty_1_80 = _RAND_1616[0:0];
  _RAND_1617 = {1{`RANDOM}};
  dirty_1_81 = _RAND_1617[0:0];
  _RAND_1618 = {1{`RANDOM}};
  dirty_1_82 = _RAND_1618[0:0];
  _RAND_1619 = {1{`RANDOM}};
  dirty_1_83 = _RAND_1619[0:0];
  _RAND_1620 = {1{`RANDOM}};
  dirty_1_84 = _RAND_1620[0:0];
  _RAND_1621 = {1{`RANDOM}};
  dirty_1_85 = _RAND_1621[0:0];
  _RAND_1622 = {1{`RANDOM}};
  dirty_1_86 = _RAND_1622[0:0];
  _RAND_1623 = {1{`RANDOM}};
  dirty_1_87 = _RAND_1623[0:0];
  _RAND_1624 = {1{`RANDOM}};
  dirty_1_88 = _RAND_1624[0:0];
  _RAND_1625 = {1{`RANDOM}};
  dirty_1_89 = _RAND_1625[0:0];
  _RAND_1626 = {1{`RANDOM}};
  dirty_1_90 = _RAND_1626[0:0];
  _RAND_1627 = {1{`RANDOM}};
  dirty_1_91 = _RAND_1627[0:0];
  _RAND_1628 = {1{`RANDOM}};
  dirty_1_92 = _RAND_1628[0:0];
  _RAND_1629 = {1{`RANDOM}};
  dirty_1_93 = _RAND_1629[0:0];
  _RAND_1630 = {1{`RANDOM}};
  dirty_1_94 = _RAND_1630[0:0];
  _RAND_1631 = {1{`RANDOM}};
  dirty_1_95 = _RAND_1631[0:0];
  _RAND_1632 = {1{`RANDOM}};
  dirty_1_96 = _RAND_1632[0:0];
  _RAND_1633 = {1{`RANDOM}};
  dirty_1_97 = _RAND_1633[0:0];
  _RAND_1634 = {1{`RANDOM}};
  dirty_1_98 = _RAND_1634[0:0];
  _RAND_1635 = {1{`RANDOM}};
  dirty_1_99 = _RAND_1635[0:0];
  _RAND_1636 = {1{`RANDOM}};
  dirty_1_100 = _RAND_1636[0:0];
  _RAND_1637 = {1{`RANDOM}};
  dirty_1_101 = _RAND_1637[0:0];
  _RAND_1638 = {1{`RANDOM}};
  dirty_1_102 = _RAND_1638[0:0];
  _RAND_1639 = {1{`RANDOM}};
  dirty_1_103 = _RAND_1639[0:0];
  _RAND_1640 = {1{`RANDOM}};
  dirty_1_104 = _RAND_1640[0:0];
  _RAND_1641 = {1{`RANDOM}};
  dirty_1_105 = _RAND_1641[0:0];
  _RAND_1642 = {1{`RANDOM}};
  dirty_1_106 = _RAND_1642[0:0];
  _RAND_1643 = {1{`RANDOM}};
  dirty_1_107 = _RAND_1643[0:0];
  _RAND_1644 = {1{`RANDOM}};
  dirty_1_108 = _RAND_1644[0:0];
  _RAND_1645 = {1{`RANDOM}};
  dirty_1_109 = _RAND_1645[0:0];
  _RAND_1646 = {1{`RANDOM}};
  dirty_1_110 = _RAND_1646[0:0];
  _RAND_1647 = {1{`RANDOM}};
  dirty_1_111 = _RAND_1647[0:0];
  _RAND_1648 = {1{`RANDOM}};
  dirty_1_112 = _RAND_1648[0:0];
  _RAND_1649 = {1{`RANDOM}};
  dirty_1_113 = _RAND_1649[0:0];
  _RAND_1650 = {1{`RANDOM}};
  dirty_1_114 = _RAND_1650[0:0];
  _RAND_1651 = {1{`RANDOM}};
  dirty_1_115 = _RAND_1651[0:0];
  _RAND_1652 = {1{`RANDOM}};
  dirty_1_116 = _RAND_1652[0:0];
  _RAND_1653 = {1{`RANDOM}};
  dirty_1_117 = _RAND_1653[0:0];
  _RAND_1654 = {1{`RANDOM}};
  dirty_1_118 = _RAND_1654[0:0];
  _RAND_1655 = {1{`RANDOM}};
  dirty_1_119 = _RAND_1655[0:0];
  _RAND_1656 = {1{`RANDOM}};
  dirty_1_120 = _RAND_1656[0:0];
  _RAND_1657 = {1{`RANDOM}};
  dirty_1_121 = _RAND_1657[0:0];
  _RAND_1658 = {1{`RANDOM}};
  dirty_1_122 = _RAND_1658[0:0];
  _RAND_1659 = {1{`RANDOM}};
  dirty_1_123 = _RAND_1659[0:0];
  _RAND_1660 = {1{`RANDOM}};
  dirty_1_124 = _RAND_1660[0:0];
  _RAND_1661 = {1{`RANDOM}};
  dirty_1_125 = _RAND_1661[0:0];
  _RAND_1662 = {1{`RANDOM}};
  dirty_1_126 = _RAND_1662[0:0];
  _RAND_1663 = {1{`RANDOM}};
  dirty_1_127 = _RAND_1663[0:0];
  _RAND_1664 = {1{`RANDOM}};
  way0_hit = _RAND_1664[0:0];
  _RAND_1665 = {1{`RANDOM}};
  way1_hit = _RAND_1665[0:0];
  _RAND_1666 = {2{`RANDOM}};
  write_back_data = _RAND_1666[63:0];
  _RAND_1667 = {1{`RANDOM}};
  write_back_addr = _RAND_1667[31:0];
  _RAND_1668 = {1{`RANDOM}};
  unuse_way = _RAND_1668[1:0];
  _RAND_1669 = {2{`RANDOM}};
  receive_data = _RAND_1669[63:0];
  _RAND_1670 = {1{`RANDOM}};
  quene = _RAND_1670[0:0];
  _RAND_1671 = {1{`RANDOM}};
  state = _RAND_1671[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IDU(
  input  [31:0] io_inst,
  output [31:0] io_inst_now,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2,
  output [4:0]  io_rd,
  output [63:0] io_imm,
  output        io_ctrl_sign_reg_write,
  output        io_ctrl_sign_csr_write,
  output        io_ctrl_sign_src2_is_imm,
  output        io_ctrl_sign_src1_is_pc,
  output        io_ctrl_sign_Writemem_en,
  output        io_ctrl_sign_Readmem_en,
  output [7:0]  io_ctrl_sign_Wmask
);
  wire [4:0] rd = io_inst[11:7]; // @[IDU.scala 150:15]
  wire [31:0] _inst_type_T = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_1 = 32'h13 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_2 = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_3 = 32'h17 == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_5 = 32'h37 == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_7 = 32'h6f == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_9 = 32'h67 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_11 = 32'h3023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_13 = 32'h3013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_15 = 32'h2003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_16 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_17 = 32'h3b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_19 = 32'h40000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_21 = 32'h1063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_23 = 32'h63 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_25 = 32'h3003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_27 = 32'h1b == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_29 = 32'h33 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_30 = io_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_31 = 32'h40005013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_33 = 32'h4003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_35 = 32'h1023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_37 = 32'h23 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_39 = 32'h6033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_41 = 32'h4013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_43 = 32'h7033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_45 = 32'h7013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_47 = 32'h4000003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_49 = 32'h103b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_51 = 32'h1013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_53 = 32'h5013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_55 = 32'h101b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_57 = 32'h4000501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_59 = 32'h501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_61 = 32'h4000503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_63 = 32'h503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_65 = 32'h3033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_67 = 32'h2033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_69 = 32'h5063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_71 = 32'h4063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_73 = 32'h6063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_75 = 32'h2023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_77 = 32'h1003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_79 = 32'h5003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_81 = 32'h2000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_83 = 32'h200003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_85 = 32'h200403b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_87 = 32'h200603b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_89 = 32'h4033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_91 = 32'h6013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_93 = 32'h2005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_95 = 32'h2004033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_97 = 32'h200503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_99 = 32'h200703b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_101 = 32'h2007033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_103 = 32'h2006033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_105 = 32'h1033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_107 = 32'h5033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_109 = 32'h40005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_111 = 32'h2013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_113 = 32'h6003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_115 = 32'h3 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_117 = 32'h7063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_119 = 32'h73 == io_inst; // @[Lookup.scala 31:38]
  wire  _inst_type_T_121 = 32'h1073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_123 = 32'h2073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_125 = 32'h3073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [6:0] _inst_type_T_126 = _inst_type_T_125 ? 7'h40 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_127 = _inst_type_T_123 ? 7'h40 : _inst_type_T_126; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_128 = _inst_type_T_121 ? 7'h40 : _inst_type_T_127; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_129 = _inst_type_T_119 ? 7'h40 : _inst_type_T_128; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_130 = _inst_type_T_117 ? 7'h45 : _inst_type_T_129; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_131 = _inst_type_T_115 ? 7'h40 : _inst_type_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_132 = _inst_type_T_113 ? 7'h40 : _inst_type_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_133 = _inst_type_T_111 ? 7'h40 : _inst_type_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_134 = _inst_type_T_109 ? 7'h41 : _inst_type_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_135 = _inst_type_T_107 ? 7'h41 : _inst_type_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_136 = _inst_type_T_105 ? 7'h41 : _inst_type_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_137 = _inst_type_T_103 ? 7'h41 : _inst_type_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_138 = _inst_type_T_101 ? 7'h41 : _inst_type_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_139 = _inst_type_T_99 ? 7'h41 : _inst_type_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_140 = _inst_type_T_97 ? 7'h41 : _inst_type_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_141 = _inst_type_T_95 ? 7'h41 : _inst_type_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_142 = _inst_type_T_93 ? 7'h41 : _inst_type_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_143 = _inst_type_T_91 ? 7'h40 : _inst_type_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_144 = _inst_type_T_89 ? 7'h41 : _inst_type_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_145 = _inst_type_T_87 ? 7'h41 : _inst_type_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_146 = _inst_type_T_85 ? 7'h41 : _inst_type_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_147 = _inst_type_T_83 ? 7'h41 : _inst_type_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_148 = _inst_type_T_81 ? 7'h41 : _inst_type_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_149 = _inst_type_T_79 ? 7'h40 : _inst_type_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_150 = _inst_type_T_77 ? 7'h40 : _inst_type_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_151 = _inst_type_T_75 ? 7'h44 : _inst_type_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_152 = _inst_type_T_73 ? 7'h45 : _inst_type_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_153 = _inst_type_T_71 ? 7'h45 : _inst_type_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_154 = _inst_type_T_69 ? 7'h45 : _inst_type_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_155 = _inst_type_T_67 ? 7'h41 : _inst_type_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_156 = _inst_type_T_65 ? 7'h41 : _inst_type_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_157 = _inst_type_T_63 ? 7'h41 : _inst_type_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_158 = _inst_type_T_61 ? 7'h41 : _inst_type_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_159 = _inst_type_T_59 ? 7'h40 : _inst_type_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_160 = _inst_type_T_57 ? 7'h40 : _inst_type_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_161 = _inst_type_T_55 ? 7'h40 : _inst_type_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_162 = _inst_type_T_53 ? 7'h40 : _inst_type_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_163 = _inst_type_T_51 ? 7'h40 : _inst_type_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_164 = _inst_type_T_49 ? 7'h41 : _inst_type_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_165 = _inst_type_T_47 ? 7'h41 : _inst_type_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_166 = _inst_type_T_45 ? 7'h40 : _inst_type_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_167 = _inst_type_T_43 ? 7'h41 : _inst_type_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_168 = _inst_type_T_41 ? 7'h40 : _inst_type_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_169 = _inst_type_T_39 ? 7'h41 : _inst_type_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_170 = _inst_type_T_37 ? 7'h44 : _inst_type_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_171 = _inst_type_T_35 ? 7'h44 : _inst_type_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_172 = _inst_type_T_33 ? 7'h40 : _inst_type_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_173 = _inst_type_T_31 ? 7'h40 : _inst_type_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_174 = _inst_type_T_29 ? 7'h41 : _inst_type_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_175 = _inst_type_T_27 ? 7'h40 : _inst_type_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_176 = _inst_type_T_25 ? 7'h40 : _inst_type_T_175; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_177 = _inst_type_T_23 ? 7'h45 : _inst_type_T_176; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_178 = _inst_type_T_21 ? 7'h45 : _inst_type_T_177; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_179 = _inst_type_T_19 ? 7'h41 : _inst_type_T_178; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_180 = _inst_type_T_17 ? 7'h41 : _inst_type_T_179; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_181 = _inst_type_T_15 ? 7'h40 : _inst_type_T_180; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_182 = _inst_type_T_13 ? 7'h40 : _inst_type_T_181; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_183 = _inst_type_T_11 ? 7'h44 : _inst_type_T_182; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_184 = _inst_type_T_9 ? 7'h40 : _inst_type_T_183; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_185 = _inst_type_T_7 ? 7'h43 : _inst_type_T_184; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_186 = _inst_type_T_5 ? 7'h42 : _inst_type_T_185; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_187 = _inst_type_T_3 ? 7'h42 : _inst_type_T_186; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_188 = _inst_type_T_1 ? 7'h40 : _inst_type_T_187; // @[Lookup.scala 34:39]
  wire [11:0] imm_imm = io_inst[31:20]; // @[IDU.scala 24:23]
  wire [51:0] _imm_T_2 = imm_imm[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_3 = {_imm_T_2,imm_imm}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_1 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21]}; // @[Cat.scala 31:58]
  wire [42:0] _imm_T_6 = imm_imm_1[19] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_7 = {_imm_T_6,io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_2 = io_inst[31:12]; // @[IDU.scala 28:23]
  wire [31:0] _imm_T_10 = imm_imm_2[19] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_12 = {_imm_T_10,imm_imm_2,12'h0}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_3 = {io_inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [51:0] _imm_T_15 = imm_imm_3[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_16 = {_imm_T_15,io_inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_4 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8]}; // @[Cat.scala 31:58]
  wire [50:0] _imm_T_19 = imm_imm_4[11] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_20 = {_imm_T_19,io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] inst_type = {{25'd0}, _inst_type_T_188}; // @[IDU.scala 133:25 152:15]
  wire [63:0] _imm_T_22 = 32'h40 == inst_type ? _imm_T_3 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_24 = 32'h43 == inst_type ? _imm_T_7 : _imm_T_22; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_26 = 32'h42 == inst_type ? _imm_T_12 : _imm_T_24; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_28 = 32'h44 == inst_type ? _imm_T_16 : _imm_T_26; // @[Mux.scala 81:58]
  wire  _inst_now_T_3 = 32'h100073 == io_inst; // @[Lookup.scala 31:38]
  wire  _inst_now_T_123 = 32'h30200073 == io_inst; // @[Lookup.scala 31:38]
  wire [6:0] _inst_now_T_130 = _inst_type_T_125 ? 7'h47 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_131 = _inst_type_T_123 ? 7'h46 : _inst_now_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_132 = _inst_type_T_121 ? 7'h3f : _inst_now_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_133 = _inst_now_T_123 ? 7'h3e : _inst_now_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_134 = _inst_type_T_119 ? 7'h3d : _inst_now_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_135 = _inst_type_T_117 ? 7'h3c : _inst_now_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_136 = _inst_type_T_115 ? 7'h3b : _inst_now_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_137 = _inst_type_T_113 ? 7'h3a : _inst_now_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_138 = _inst_type_T_111 ? 7'h36 : _inst_now_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_139 = _inst_type_T_109 ? 7'h39 : _inst_now_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_140 = _inst_type_T_107 ? 7'h38 : _inst_now_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_141 = _inst_type_T_105 ? 7'h37 : _inst_now_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_142 = _inst_type_T_103 ? 7'h34 : _inst_now_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_143 = _inst_type_T_101 ? 7'h33 : _inst_now_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_144 = _inst_type_T_99 ? 7'h32 : _inst_now_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_145 = _inst_type_T_97 ? 7'h35 : _inst_now_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_146 = _inst_type_T_95 ? 7'h31 : _inst_now_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_147 = _inst_type_T_93 ? 7'h30 : _inst_now_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_148 = _inst_type_T_91 ? 7'h2f : _inst_now_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_149 = _inst_type_T_89 ? 7'h2e : _inst_now_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_150 = _inst_type_T_87 ? 7'h14 : _inst_now_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_151 = _inst_type_T_85 ? 7'h13 : _inst_now_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_152 = _inst_type_T_83 ? 7'h12 : _inst_now_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_153 = _inst_type_T_81 ? 7'h11 : _inst_now_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_154 = _inst_type_T_79 ? 7'h25 : _inst_now_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_155 = _inst_type_T_77 ? 7'h24 : _inst_now_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_156 = _inst_type_T_75 ? 7'h27 : _inst_now_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_157 = _inst_type_T_73 ? 7'h2d : _inst_now_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_158 = _inst_type_T_71 ? 7'h2c : _inst_now_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_159 = _inst_type_T_69 ? 7'h2b : _inst_now_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_160 = _inst_type_T_67 ? 7'h1f : _inst_now_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_161 = _inst_type_T_65 ? 7'h1e : _inst_now_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_162 = _inst_type_T_63 ? 7'h1d : _inst_now_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_163 = _inst_type_T_61 ? 7'h1c : _inst_now_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_164 = _inst_type_T_59 ? 7'h1b : _inst_now_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_165 = _inst_type_T_57 ? 7'h1a : _inst_now_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_166 = _inst_type_T_55 ? 7'h19 : _inst_now_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_167 = _inst_type_T_53 ? 7'h18 : _inst_now_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_168 = _inst_type_T_51 ? 7'h17 : _inst_now_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_169 = _inst_type_T_49 ? 7'h16 : _inst_now_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_170 = _inst_type_T_47 ? 7'hd : _inst_now_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_171 = _inst_type_T_45 ? 7'h9 : _inst_now_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_172 = _inst_type_T_43 ? 7'h8 : _inst_now_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_173 = _inst_type_T_41 ? 7'ha : _inst_now_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_174 = _inst_type_T_39 ? 7'hb : _inst_now_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_175 = _inst_type_T_37 ? 7'h28 : _inst_now_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_176 = _inst_type_T_35 ? 7'h26 : _inst_now_T_175; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_177 = _inst_type_T_33 ? 7'h23 : _inst_now_T_176; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_178 = _inst_type_T_31 ? 7'h15 : _inst_now_T_177; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_179 = _inst_type_T_29 ? 7'hf : _inst_now_T_178; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_180 = _inst_type_T_27 ? 7'h10 : _inst_now_T_179; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_181 = _inst_type_T_25 ? 7'h22 : _inst_now_T_180; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_182 = _inst_type_T_23 ? 7'h29 : _inst_now_T_181; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_183 = _inst_type_T_21 ? 7'h2a : _inst_now_T_182; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_184 = _inst_type_T_19 ? 7'he : _inst_now_T_183; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_185 = _inst_type_T_17 ? 7'hc : _inst_now_T_184; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_186 = _inst_type_T_15 ? 7'h21 : _inst_now_T_185; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_187 = _inst_type_T_13 ? 7'h20 : _inst_now_T_186; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_188 = _inst_type_T_11 ? 7'h7 : _inst_now_T_187; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_189 = _inst_type_T_9 ? 7'h6 : _inst_now_T_188; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_190 = _inst_type_T_7 ? 7'h5 : _inst_now_T_189; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_191 = _inst_type_T_5 ? 7'h4 : _inst_now_T_190; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_192 = _inst_type_T_3 ? 7'h3 : _inst_now_T_191; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_193 = _inst_now_T_3 ? 7'h2 : _inst_now_T_192; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_194 = _inst_type_T_1 ? 7'h1 : _inst_now_T_193; // @[Lookup.scala 34:39]
  wire  _reg_write_T_26 = _inst_now_T_123 ? 1'h0 : 1'h1; // @[Lookup.scala 34:39]
  wire  _reg_write_T_27 = _inst_type_T_119 ? 1'h0 : _reg_write_T_26; // @[Lookup.scala 34:39]
  wire  _reg_write_T_28 = _inst_type_T_117 ? 1'h0 : _reg_write_T_27; // @[Lookup.scala 34:39]
  wire  _reg_write_T_29 = _inst_type_T_73 ? 1'h0 : _reg_write_T_28; // @[Lookup.scala 34:39]
  wire  _reg_write_T_30 = _inst_type_T_71 ? 1'h0 : _reg_write_T_29; // @[Lookup.scala 34:39]
  wire  _reg_write_T_31 = _inst_type_T_69 ? 1'h0 : _reg_write_T_30; // @[Lookup.scala 34:39]
  wire  _reg_write_T_32 = _inst_type_T_23 ? 1'h0 : _reg_write_T_31; // @[Lookup.scala 34:39]
  wire  _reg_write_T_33 = _inst_type_T_21 ? 1'h0 : _reg_write_T_32; // @[Lookup.scala 34:39]
  wire  _reg_write_T_34 = _inst_type_T_75 ? 1'h0 : _reg_write_T_33; // @[Lookup.scala 34:39]
  wire  _reg_write_T_35 = _inst_type_T_37 ? 1'h0 : _reg_write_T_34; // @[Lookup.scala 34:39]
  wire  _reg_write_T_36 = _inst_type_T_35 ? 1'h0 : _reg_write_T_35; // @[Lookup.scala 34:39]
  wire  _reg_write_T_37 = _inst_type_T_11 ? 1'h0 : _reg_write_T_36; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_8 = _inst_type_T_75 ? 4'hf : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_9 = _inst_type_T_37 ? 4'h1 : _Wmask_T_8; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_10 = _inst_type_T_35 ? 4'h3 : _Wmask_T_9; // @[Lookup.scala 34:39]
  assign io_inst_now = {{25'd0}, _inst_now_T_194}; // @[IDU.scala 132:24 226:14]
  assign io_rs1 = io_inst[19:15]; // @[IDU.scala 149:16]
  assign io_rs2 = io_inst[24:20]; // @[IDU.scala 148:16]
  assign io_rd = io_inst[11:7]; // @[IDU.scala 150:15]
  assign io_imm = 32'h45 == inst_type ? _imm_T_20 : _imm_T_28; // @[Mux.scala 81:58]
  assign io_ctrl_sign_reg_write = _inst_now_T_3 ? 1'h0 : _reg_write_T_37; // @[Lookup.scala 34:39]
  assign io_ctrl_sign_csr_write = _inst_type_T_121 | (_inst_type_T_123 | _inst_type_T_125); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_src2_is_imm = 32'h45 == inst_type | (32'h43 == inst_type | (32'h44 == inst_type | (32'h42 ==
    inst_type | 32'h40 == inst_type))); // @[Mux.scala 81:58]
  assign io_ctrl_sign_src1_is_pc = _inst_type_T_7 | (_inst_type_T_3 | (_inst_type_T_21 | (_inst_type_T_23 | (
    _inst_type_T_69 | (_inst_type_T_71 | (_inst_type_T_73 | _inst_type_T_117)))))); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Writemem_en = 32'h44 == inst_type; // @[Mux.scala 81:61]
  assign io_ctrl_sign_Readmem_en = _inst_type_T_25 | (_inst_type_T_15 | (_inst_type_T_113 | (_inst_type_T_77 | (
    _inst_type_T_79 | (_inst_type_T_115 | _inst_type_T_33))))); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Wmask = _inst_type_T_11 ? 8'hff : {{4'd0}, _Wmask_T_10}; // @[Lookup.scala 34:39]
endmodule
module EXU_AXI(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  output [63:0] io_pc_next,
  input  [31:0] io_inst_now,
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [4:0]  io_rd,
  input  [63:0] io_imm,
  input         io_ctrl_sign_reg_write,
  input         io_ctrl_sign_csr_write,
  input         io_ctrl_sign_src2_is_imm,
  input         io_ctrl_sign_src1_is_pc,
  input         io_ctrl_sign_Writemem_en,
  input         io_ctrl_sign_Readmem_en,
  input  [7:0]  io_ctrl_sign_Wmask,
  output [63:0] io_res2rd,
  input         io_inst_valid,
  output        io_inst_store,
  output        io_inst_load,
  output [31:0] io_Mem_addr,
  input  [63:0] io_Mem_rdata,
  output [63:0] io_Mem_wdata,
  output [7:0]  io_Mem_wstrb,
  input         io_rdata_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] Regfile [0:31]; // @[EXU_AXI.scala 37:22]
  wire  Regfile_src1_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_src1_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_src1_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_src2_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_src2_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_src2_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_4_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_MPORT_4_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_MPORT_4_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_1_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_1_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_1_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_2_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_2_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_2_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_3_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_3_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_3_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_4_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_4_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_4_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_5_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_5_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_5_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_6_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_6_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_6_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_7_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_7_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_7_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_8_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_8_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_8_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_9_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_9_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_9_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_10_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_10_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_10_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_11_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_11_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_11_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_0_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_0_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_0_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_1_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_1_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_1_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_2_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_2_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_2_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_3_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_3_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_3_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_4_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_4_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_4_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_5_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_5_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_5_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_6_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_6_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_6_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_7_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_7_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_7_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_8_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_8_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_8_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_9_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_9_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_9_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_10_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_10_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_10_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_11_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_11_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_11_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_12_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_12_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_12_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_13_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_13_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_13_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_14_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_14_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_14_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_15_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_15_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_15_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_16_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_16_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_16_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_17_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_17_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_17_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_18_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_18_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_18_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_19_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_19_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_19_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_20_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_20_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_20_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_21_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_21_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_21_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_22_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_22_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_22_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_23_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_23_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_23_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_24_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_24_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_24_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_25_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_25_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_25_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_26_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_26_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_26_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_27_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_27_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_27_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_28_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_28_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_28_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_29_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_29_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_29_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_30_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_30_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_30_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_31_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_31_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_31_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_1_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_1_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_1_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_2_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_2_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_2_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_3_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_3_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_3_data; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_mask; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_en; // @[EXU_AXI.scala 37:22]
  reg [63:0] CSR_Reg [0:3]; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_2_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_2_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_2_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_csr_wdata_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_csr_wdata_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_csr_wdata_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_csr_wdata_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_csr_wdata_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_csr_wdata_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_2_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_2_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_2_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_5_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_5_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_5_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_7_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_7_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_7_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_j_pc_MPORT_12_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_j_pc_MPORT_12_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_j_pc_MPORT_12_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_j_pc_MPORT_13_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_j_pc_MPORT_13_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_j_pc_MPORT_13_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_0_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_1_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_2_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_1_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_3_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_3_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_3_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_3_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_6_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_6_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_6_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_6_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] reg_trace_input_reg_0; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_1; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_2; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_3; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_4; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_5; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_6; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_7; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_8; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_9; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_10; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_11; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_12; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_13; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_14; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_15; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_16; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_17; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_18; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_19; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_20; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_21; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_22; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_23; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_24; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_25; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_26; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_27; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_28; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_29; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_30; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_31; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_0; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_1; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_2; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_3; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_pc; // @[EXU_AXI.scala 163:27]
  wire [11:0] csr_addr = io_imm[11:0]; // @[EXU_AXI.scala 39:26]
  wire [1:0] _csr_index_T_5 = 12'h300 == csr_addr ? 2'h2 : {{1'd0}, 12'h341 == csr_addr}; // @[Mux.scala 81:58]
  wire  _csr_index_T_6 = 12'h342 == csr_addr; // @[Mux.scala 81:61]
  wire [63:0] _src1_value_T_1 = io_rs1 == 5'h0 ? 64'h0 : Regfile_src1_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] src1_value = io_ctrl_sign_src1_is_pc ? io_pc : _src1_value_T_1; // @[EXU_AXI.scala 49:25]
  wire [63:0] _src2_value_T_1 = io_rs2 == 5'h0 ? 64'h0 : Regfile_src2_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] src2_value = io_ctrl_sign_src2_is_imm ? io_imm : _src2_value_T_1; // @[EXU_AXI.scala 50:25]
  wire [63:0] add_res = src1_value + src2_value; // @[EXU_AXI.scala 51:30]
  wire [63:0] sub_res = src1_value - src2_value; // @[EXU_AXI.scala 52:30]
  wire [63:0] _sra_res_T = io_ctrl_sign_src1_is_pc ? io_pc : _src1_value_T_1; // @[EXU_AXI.scala 53:37]
  wire [63:0] sra_res = $signed(_sra_res_T) >>> src2_value[5:0]; // @[EXU_AXI.scala 53:60]
  wire [63:0] srl_res = src1_value >> src2_value[5:0]; // @[EXU_AXI.scala 54:30]
  wire [126:0] _GEN_1 = {{63'd0}, src1_value}; // @[EXU_AXI.scala 55:30]
  wire [126:0] sll_res = _GEN_1 << src2_value[5:0]; // @[EXU_AXI.scala 55:30]
  wire [31:0] _sraw_res_T_1 = src1_value[31:0]; // @[EXU_AXI.scala 56:43]
  wire [31:0] sraw_res = $signed(_sraw_res_T_1) >>> src2_value[4:0]; // @[EXU_AXI.scala 56:46]
  wire [31:0] srlw_res = src1_value[31:0] >> src2_value[4:0]; // @[EXU_AXI.scala 57:37]
  wire [62:0] _GEN_2 = {{31'd0}, src1_value[31:0]}; // @[EXU_AXI.scala 58:37]
  wire [62:0] sllw_res = _GEN_2 << src2_value[4:0]; // @[EXU_AXI.scala 58:37]
  wire [63:0] or_res = src1_value | src2_value; // @[EXU_AXI.scala 59:29]
  wire [63:0] xor_res = src1_value ^ src2_value; // @[EXU_AXI.scala 60:30]
  wire [63:0] and_res = src1_value & src2_value; // @[EXU_AXI.scala 61:30]
  wire [127:0] _mlu_res_T = src1_value * src2_value; // @[EXU_AXI.scala 62:31]
  wire [63:0] mlu_res = _mlu_res_T[63:0]; // @[EXU_AXI.scala 62:44]
  wire [63:0] _mluw_res_T_2 = src1_value[31:0] * src2_value[31:0]; // @[EXU_AXI.scala 63:38]
  wire [31:0] mluw_res = _mluw_res_T_2[31:0]; // @[EXU_AXI.scala 63:57]
  wire [31:0] _divw_res_T_3 = src2_value[31:0]; // @[EXU_AXI.scala 64:64]
  wire [32:0] _divw_res_T_4 = $signed(_sraw_res_T_1) / $signed(_divw_res_T_3); // @[EXU_AXI.scala 64:45]
  wire [31:0] divw_res = _divw_res_T_4[31:0]; // @[EXU_AXI.scala 64:71]
  wire [31:0] divuw_res = src1_value[31:0] / src2_value[31:0]; // @[EXU_AXI.scala 65:39]
  wire [31:0] remw_res = $signed(_sraw_res_T_1) % $signed(_divw_res_T_3); // @[EXU_AXI.scala 66:71]
  wire [31:0] remuw_res = src1_value[31:0] % src2_value[31:0]; // @[EXU_AXI.scala 67:39]
  wire [63:0] _div_res_T_1 = io_ctrl_sign_src2_is_imm ? io_imm : _src2_value_T_1; // @[EXU_AXI.scala 68:51]
  wire [64:0] div_res = $signed(_sra_res_T) / $signed(_div_res_T_1); // @[EXU_AXI.scala 68:59]
  wire [63:0] divu_res = src1_value / src2_value; // @[EXU_AXI.scala 69:31]
  wire [63:0] rem_res = $signed(_sra_res_T) % $signed(_div_res_T_1); // @[EXU_AXI.scala 70:59]
  wire [63:0] remu_res = src1_value % src2_value; // @[EXU_AXI.scala 71:31]
  wire [63:0] _io_res2rd_T_1 = io_pc + 64'h4; // @[EXU_AXI.scala 76:24]
  wire  _io_res2rd_T_4 = src1_value < src2_value; // @[EXU_AXI.scala 78:34]
  wire  _io_res2rd_T_10 = $signed(_sra_res_T) < $signed(_div_res_T_1); // @[EXU_AXI.scala 80:42]
  wire [31:0] _io_res2rd_T_18 = io_Mem_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_20 = {_io_res2rd_T_18,io_Mem_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_23 = {56'h0,io_Mem_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_26 = {32'h0,io_Mem_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [47:0] _io_res2rd_T_29 = io_Mem_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_31 = {_io_res2rd_T_29,io_Mem_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [55:0] _io_res2rd_T_34 = io_Mem_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_36 = {_io_res2rd_T_34,io_Mem_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_39 = {48'h0,io_Mem_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_42 = add_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_44 = {_io_res2rd_T_42,add_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_52 = sub_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_54 = {_io_res2rd_T_52,sub_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_57 = sllw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_59 = {_io_res2rd_T_57,sllw_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_67 = sraw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _io_res2rd_T_68 = $signed(_sraw_res_T_1) >>> src2_value[4:0]; // @[EXU_AXI.scala 105:56]
  wire [63:0] _io_res2rd_T_69 = {_io_res2rd_T_67,_io_res2rd_T_68}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_72 = srlw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_74 = {_io_res2rd_T_72,srlw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_87 = mluw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_88 = {_io_res2rd_T_87,mluw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_91 = divw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_92 = {_io_res2rd_T_91,divw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_95 = divuw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_96 = {_io_res2rd_T_95,divuw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_99 = remw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_100 = {_io_res2rd_T_99,remw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_103 = remuw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_104 = {_io_res2rd_T_103,remuw_res}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_106 = 32'h1 == io_inst_now ? add_res : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_108 = 32'h3 == io_inst_now ? add_res : _io_res2rd_T_106; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_110 = 32'h4 == io_inst_now ? io_imm : _io_res2rd_T_108; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_112 = 32'h5 == io_inst_now ? _io_res2rd_T_1 : _io_res2rd_T_110; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_114 = 32'h6 == io_inst_now ? _io_res2rd_T_1 : _io_res2rd_T_112; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_116 = 32'h20 == io_inst_now ? {{63'd0}, _io_res2rd_T_4} : _io_res2rd_T_114; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_118 = 32'h1e == io_inst_now ? {{63'd0}, _io_res2rd_T_4} : _io_res2rd_T_116; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_120 = 32'h36 == io_inst_now ? {{63'd0}, _io_res2rd_T_10} : _io_res2rd_T_118; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_122 = 32'h1f == io_inst_now ? {{63'd0}, _io_res2rd_T_10} : _io_res2rd_T_120; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_124 = 32'h21 == io_inst_now ? _io_res2rd_T_20 : _io_res2rd_T_122; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_126 = 32'h22 == io_inst_now ? io_Mem_rdata : _io_res2rd_T_124; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_128 = 32'h23 == io_inst_now ? _io_res2rd_T_23 : _io_res2rd_T_126; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_130 = 32'h3a == io_inst_now ? _io_res2rd_T_26 : _io_res2rd_T_128; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_132 = 32'h24 == io_inst_now ? _io_res2rd_T_31 : _io_res2rd_T_130; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_134 = 32'h3b == io_inst_now ? _io_res2rd_T_36 : _io_res2rd_T_132; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_136 = 32'h25 == io_inst_now ? _io_res2rd_T_39 : _io_res2rd_T_134; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_138 = 32'hc == io_inst_now ? _io_res2rd_T_44 : _io_res2rd_T_136; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_140 = 32'he == io_inst_now ? sub_res : _io_res2rd_T_138; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_142 = 32'h10 == io_inst_now ? _io_res2rd_T_44 : _io_res2rd_T_140; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_144 = 32'hf == io_inst_now ? add_res : _io_res2rd_T_142; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_146 = 32'h15 == io_inst_now ? sra_res : _io_res2rd_T_144; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_148 = 32'hb == io_inst_now ? or_res : _io_res2rd_T_146; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_150 = 32'h2f == io_inst_now ? or_res : _io_res2rd_T_148; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_152 = 32'h2e == io_inst_now ? xor_res : _io_res2rd_T_150; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_154 = 32'ha == io_inst_now ? xor_res : _io_res2rd_T_152; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_156 = 32'h8 == io_inst_now ? and_res : _io_res2rd_T_154; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_158 = 32'h9 == io_inst_now ? and_res : _io_res2rd_T_156; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_160 = 32'hd == io_inst_now ? _io_res2rd_T_54 : _io_res2rd_T_158; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_162 = 32'h16 == io_inst_now ? _io_res2rd_T_59 : _io_res2rd_T_160; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_164 = 32'h17 == io_inst_now ? sll_res : {{63'd0}, _io_res2rd_T_162}; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_166 = 32'h18 == io_inst_now ? {{63'd0}, srl_res} : _io_res2rd_T_164; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_168 = 32'h19 == io_inst_now ? {{63'd0}, _io_res2rd_T_59} : _io_res2rd_T_166; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_170 = 32'h1a == io_inst_now ? {{63'd0}, _io_res2rd_T_69} : _io_res2rd_T_168; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_172 = 32'h1b == io_inst_now ? {{63'd0}, _io_res2rd_T_74} : _io_res2rd_T_170; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_174 = 32'h1c == io_inst_now ? {{63'd0}, _io_res2rd_T_69} : _io_res2rd_T_172; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_176 = 32'h1d == io_inst_now ? {{63'd0}, _io_res2rd_T_74} : _io_res2rd_T_174; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_178 = 32'h11 == io_inst_now ? {{63'd0}, mlu_res} : _io_res2rd_T_176; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_180 = 32'h12 == io_inst_now ? {{63'd0}, _io_res2rd_T_88} : _io_res2rd_T_178; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_182 = 32'h13 == io_inst_now ? {{63'd0}, _io_res2rd_T_92} : _io_res2rd_T_180; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_184 = 32'h30 == io_inst_now ? {{63'd0}, divu_res} : _io_res2rd_T_182; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_186 = 32'h31 == io_inst_now ? {{62'd0}, div_res} : _io_res2rd_T_184; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_188 = 32'h35 == io_inst_now ? {{63'd0}, _io_res2rd_T_96} : _io_res2rd_T_186; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_190 = 32'h14 == io_inst_now ? {{63'd0}, _io_res2rd_T_100} : _io_res2rd_T_188; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_192 = 32'h32 == io_inst_now ? {{63'd0}, _io_res2rd_T_104} : _io_res2rd_T_190; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_194 = 32'h33 == io_inst_now ? {{63'd0}, remu_res} : _io_res2rd_T_192; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_196 = 32'h34 == io_inst_now ? {{63'd0}, rem_res} : _io_res2rd_T_194; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_198 = 32'h37 == io_inst_now ? sll_res : _io_res2rd_T_196; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_200 = 32'h39 == io_inst_now ? {{63'd0}, sra_res} : _io_res2rd_T_198; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_202 = 32'h38 == io_inst_now ? {{63'd0}, srl_res} : _io_res2rd_T_200; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_204 = 32'h3f == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_data} : _io_res2rd_T_202; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_206 = 32'h46 == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_1_data} : _io_res2rd_T_204; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_208 = 32'h47 == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_2_data} : _io_res2rd_T_206; // @[Mux.scala 81:58]
  wire [63:0] reg_value = io_rd == 5'h0 ? 64'h0 : Regfile_reg_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire  _T_6 = io_ctrl_sign_reg_write & io_rd != 5'h0 & (io_inst_valid & ~io_ctrl_sign_Readmem_en |
    io_ctrl_sign_Readmem_en & io_rdata_valid); // @[EXU_AXI.scala 129:63]
  wire [63:0] _csr_wdata_T = src1_value | CSR_Reg_csr_wdata_MPORT_data; // @[EXU_AXI.scala 134:32]
  wire [63:0] _csr_wdata_T_1 = ~CSR_Reg_csr_wdata_MPORT_1_data; // @[EXU_AXI.scala 135:35]
  wire [63:0] _csr_wdata_T_2 = src1_value & _csr_wdata_T_1; // @[EXU_AXI.scala 135:32]
  wire [63:0] _csr_wdata_T_4 = 32'h3f == io_inst_now ? src1_value : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _csr_wdata_T_6 = 32'h46 == io_inst_now ? _csr_wdata_T : _csr_wdata_T_4; // @[Mux.scala 81:58]
  wire [63:0] csr_wdata = 32'h47 == io_inst_now ? _csr_wdata_T_2 : _csr_wdata_T_6; // @[Mux.scala 81:58]
  wire  _T_9 = io_inst_now == 32'h3d & io_inst_valid; // @[EXU_AXI.scala 138:48]
  wire  _T_14 = io_ctrl_sign_csr_write & io_inst_valid; // @[EXU_AXI.scala 141:53]
  wire [63:0] _j_pc_T = add_res & 64'hfffffffffffffffe; // @[EXU_AXI.scala 148:28]
  wire [63:0] _j_pc_T_3 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_data; // @[EXU_AXI.scala 149:39]
  wire [63:0] _j_pc_T_6 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_1_data; // @[EXU_AXI.scala 149:67]
  wire [63:0] _j_pc_T_8 = $signed(_j_pc_T_3) != $signed(_j_pc_T_6) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 149:21]
  wire [63:0] _j_pc_T_11 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_2_data; // @[EXU_AXI.scala 150:39]
  wire [63:0] _j_pc_T_14 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_3_data; // @[EXU_AXI.scala 150:67]
  wire [63:0] _j_pc_T_16 = $signed(_j_pc_T_11) == $signed(_j_pc_T_14) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 150:21]
  wire [63:0] _j_pc_T_19 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_4_data; // @[EXU_AXI.scala 151:39]
  wire [63:0] _j_pc_T_22 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_5_data; // @[EXU_AXI.scala 151:66]
  wire [63:0] _j_pc_T_24 = $signed(_j_pc_T_19) >= $signed(_j_pc_T_22) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 151:21]
  wire [63:0] _j_pc_T_27 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_6_data; // @[EXU_AXI.scala 152:39]
  wire [63:0] _j_pc_T_30 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_7_data; // @[EXU_AXI.scala 152:65]
  wire [63:0] _j_pc_T_32 = $signed(_j_pc_T_27) < $signed(_j_pc_T_30) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 152:21]
  wire [63:0] _j_pc_T_34 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_8_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_36 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_9_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_38 = _j_pc_T_34 < _j_pc_T_36 ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 153:22]
  wire [63:0] _j_pc_T_40 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_10_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_42 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_11_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_44 = _j_pc_T_40 >= _j_pc_T_42 ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 154:22]
  wire [63:0] _j_pc_T_46 = CSR_Reg_j_pc_MPORT_13_data + 64'h4; // @[EXU_AXI.scala 156:33]
  wire [63:0] _j_pc_T_48 = 32'h5 == io_inst_now ? add_res : _io_res2rd_T_1; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_50 = 32'h6 == io_inst_now ? _j_pc_T : _j_pc_T_48; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_52 = 32'h2a == io_inst_now ? _j_pc_T_8 : _j_pc_T_50; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_54 = 32'h29 == io_inst_now ? _j_pc_T_16 : _j_pc_T_52; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_56 = 32'h2b == io_inst_now ? _j_pc_T_24 : _j_pc_T_54; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_58 = 32'h2c == io_inst_now ? _j_pc_T_32 : _j_pc_T_56; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_60 = 32'h2d == io_inst_now ? _j_pc_T_38 : _j_pc_T_58; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_62 = 32'h3c == io_inst_now ? _j_pc_T_44 : _j_pc_T_60; // @[Mux.scala 81:58]
  reg [63:0] pc_next; // @[EXU_AXI.scala 158:26]
  wire [63:0] _mem_wdata_T_1 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_3 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_1_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_6 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_2_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_9 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_3_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_12 = 32'h7 == io_inst_now ? _mem_wdata_T_1 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _mem_wdata_T_14 = 32'h26 == io_inst_now ? {{48'd0}, _mem_wdata_T_3[15:0]} : _mem_wdata_T_12; // @[Mux.scala 81:58]
  wire [63:0] _mem_wdata_T_16 = 32'h28 == io_inst_now ? {{56'd0}, _mem_wdata_T_6[7:0]} : _mem_wdata_T_14; // @[Mux.scala 81:58]
  traceregs reg_trace ( // @[EXU_AXI.scala 163:27]
    .input_reg_0(reg_trace_input_reg_0),
    .input_reg_1(reg_trace_input_reg_1),
    .input_reg_2(reg_trace_input_reg_2),
    .input_reg_3(reg_trace_input_reg_3),
    .input_reg_4(reg_trace_input_reg_4),
    .input_reg_5(reg_trace_input_reg_5),
    .input_reg_6(reg_trace_input_reg_6),
    .input_reg_7(reg_trace_input_reg_7),
    .input_reg_8(reg_trace_input_reg_8),
    .input_reg_9(reg_trace_input_reg_9),
    .input_reg_10(reg_trace_input_reg_10),
    .input_reg_11(reg_trace_input_reg_11),
    .input_reg_12(reg_trace_input_reg_12),
    .input_reg_13(reg_trace_input_reg_13),
    .input_reg_14(reg_trace_input_reg_14),
    .input_reg_15(reg_trace_input_reg_15),
    .input_reg_16(reg_trace_input_reg_16),
    .input_reg_17(reg_trace_input_reg_17),
    .input_reg_18(reg_trace_input_reg_18),
    .input_reg_19(reg_trace_input_reg_19),
    .input_reg_20(reg_trace_input_reg_20),
    .input_reg_21(reg_trace_input_reg_21),
    .input_reg_22(reg_trace_input_reg_22),
    .input_reg_23(reg_trace_input_reg_23),
    .input_reg_24(reg_trace_input_reg_24),
    .input_reg_25(reg_trace_input_reg_25),
    .input_reg_26(reg_trace_input_reg_26),
    .input_reg_27(reg_trace_input_reg_27),
    .input_reg_28(reg_trace_input_reg_28),
    .input_reg_29(reg_trace_input_reg_29),
    .input_reg_30(reg_trace_input_reg_30),
    .input_reg_31(reg_trace_input_reg_31),
    .csr_reg_0(reg_trace_csr_reg_0),
    .csr_reg_1(reg_trace_csr_reg_1),
    .csr_reg_2(reg_trace_csr_reg_2),
    .csr_reg_3(reg_trace_csr_reg_3),
    .pc(reg_trace_pc)
  );
  assign Regfile_src1_value_MPORT_en = 1'h1;
  assign Regfile_src1_value_MPORT_addr = io_rs1;
  assign Regfile_src1_value_MPORT_data = Regfile[Regfile_src1_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_src2_value_MPORT_en = 1'h1;
  assign Regfile_src2_value_MPORT_addr = io_rs2;
  assign Regfile_src2_value_MPORT_data = Regfile[Regfile_src2_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_value_MPORT_en = 1'h1;
  assign Regfile_reg_value_MPORT_addr = io_rd;
  assign Regfile_reg_value_MPORT_data = Regfile[Regfile_reg_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_MPORT_4_en = 1'h1;
  assign Regfile_MPORT_4_addr = 5'h11;
  assign Regfile_MPORT_4_data = Regfile[Regfile_MPORT_4_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_en = 1'h1;
  assign Regfile_j_pc_MPORT_addr = io_rs1;
  assign Regfile_j_pc_MPORT_data = Regfile[Regfile_j_pc_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_1_en = 1'h1;
  assign Regfile_j_pc_MPORT_1_addr = io_rs2;
  assign Regfile_j_pc_MPORT_1_data = Regfile[Regfile_j_pc_MPORT_1_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_2_en = 1'h1;
  assign Regfile_j_pc_MPORT_2_addr = io_rs1;
  assign Regfile_j_pc_MPORT_2_data = Regfile[Regfile_j_pc_MPORT_2_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_3_en = 1'h1;
  assign Regfile_j_pc_MPORT_3_addr = io_rs2;
  assign Regfile_j_pc_MPORT_3_data = Regfile[Regfile_j_pc_MPORT_3_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_4_en = 1'h1;
  assign Regfile_j_pc_MPORT_4_addr = io_rs1;
  assign Regfile_j_pc_MPORT_4_data = Regfile[Regfile_j_pc_MPORT_4_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_5_en = 1'h1;
  assign Regfile_j_pc_MPORT_5_addr = io_rs2;
  assign Regfile_j_pc_MPORT_5_data = Regfile[Regfile_j_pc_MPORT_5_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_6_en = 1'h1;
  assign Regfile_j_pc_MPORT_6_addr = io_rs1;
  assign Regfile_j_pc_MPORT_6_data = Regfile[Regfile_j_pc_MPORT_6_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_7_en = 1'h1;
  assign Regfile_j_pc_MPORT_7_addr = io_rs2;
  assign Regfile_j_pc_MPORT_7_data = Regfile[Regfile_j_pc_MPORT_7_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_8_en = 1'h1;
  assign Regfile_j_pc_MPORT_8_addr = io_rs1;
  assign Regfile_j_pc_MPORT_8_data = Regfile[Regfile_j_pc_MPORT_8_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_9_en = 1'h1;
  assign Regfile_j_pc_MPORT_9_addr = io_rs2;
  assign Regfile_j_pc_MPORT_9_data = Regfile[Regfile_j_pc_MPORT_9_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_10_en = 1'h1;
  assign Regfile_j_pc_MPORT_10_addr = io_rs1;
  assign Regfile_j_pc_MPORT_10_data = Regfile[Regfile_j_pc_MPORT_10_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_11_en = 1'h1;
  assign Regfile_j_pc_MPORT_11_addr = io_rs2;
  assign Regfile_j_pc_MPORT_11_data = Regfile[Regfile_j_pc_MPORT_11_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_0_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_0_MPORT_addr = 5'h0;
  assign Regfile_reg_trace_io_input_reg_0_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_0_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_1_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_1_MPORT_addr = 5'h1;
  assign Regfile_reg_trace_io_input_reg_1_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_1_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_2_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_2_MPORT_addr = 5'h2;
  assign Regfile_reg_trace_io_input_reg_2_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_2_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_3_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_3_MPORT_addr = 5'h3;
  assign Regfile_reg_trace_io_input_reg_3_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_3_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_4_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_4_MPORT_addr = 5'h4;
  assign Regfile_reg_trace_io_input_reg_4_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_4_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_5_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_5_MPORT_addr = 5'h5;
  assign Regfile_reg_trace_io_input_reg_5_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_5_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_6_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_6_MPORT_addr = 5'h6;
  assign Regfile_reg_trace_io_input_reg_6_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_6_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_7_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_7_MPORT_addr = 5'h7;
  assign Regfile_reg_trace_io_input_reg_7_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_7_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_8_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_8_MPORT_addr = 5'h8;
  assign Regfile_reg_trace_io_input_reg_8_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_8_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_9_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_9_MPORT_addr = 5'h9;
  assign Regfile_reg_trace_io_input_reg_9_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_9_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_10_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_10_MPORT_addr = 5'ha;
  assign Regfile_reg_trace_io_input_reg_10_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_10_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_11_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_11_MPORT_addr = 5'hb;
  assign Regfile_reg_trace_io_input_reg_11_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_11_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_12_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_12_MPORT_addr = 5'hc;
  assign Regfile_reg_trace_io_input_reg_12_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_12_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_13_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_13_MPORT_addr = 5'hd;
  assign Regfile_reg_trace_io_input_reg_13_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_13_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_14_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_14_MPORT_addr = 5'he;
  assign Regfile_reg_trace_io_input_reg_14_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_14_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_15_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_15_MPORT_addr = 5'hf;
  assign Regfile_reg_trace_io_input_reg_15_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_15_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_16_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_16_MPORT_addr = 5'h10;
  assign Regfile_reg_trace_io_input_reg_16_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_16_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_17_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_17_MPORT_addr = 5'h11;
  assign Regfile_reg_trace_io_input_reg_17_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_17_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_18_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_18_MPORT_addr = 5'h12;
  assign Regfile_reg_trace_io_input_reg_18_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_18_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_19_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_19_MPORT_addr = 5'h13;
  assign Regfile_reg_trace_io_input_reg_19_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_19_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_20_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_20_MPORT_addr = 5'h14;
  assign Regfile_reg_trace_io_input_reg_20_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_20_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_21_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_21_MPORT_addr = 5'h15;
  assign Regfile_reg_trace_io_input_reg_21_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_21_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_22_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_22_MPORT_addr = 5'h16;
  assign Regfile_reg_trace_io_input_reg_22_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_22_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_23_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_23_MPORT_addr = 5'h17;
  assign Regfile_reg_trace_io_input_reg_23_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_23_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_24_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_24_MPORT_addr = 5'h18;
  assign Regfile_reg_trace_io_input_reg_24_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_24_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_25_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_25_MPORT_addr = 5'h19;
  assign Regfile_reg_trace_io_input_reg_25_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_25_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_26_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_26_MPORT_addr = 5'h1a;
  assign Regfile_reg_trace_io_input_reg_26_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_26_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_27_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_27_MPORT_addr = 5'h1b;
  assign Regfile_reg_trace_io_input_reg_27_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_27_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_28_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_28_MPORT_addr = 5'h1c;
  assign Regfile_reg_trace_io_input_reg_28_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_28_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_29_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_29_MPORT_addr = 5'h1d;
  assign Regfile_reg_trace_io_input_reg_29_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_29_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_30_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_30_MPORT_addr = 5'h1e;
  assign Regfile_reg_trace_io_input_reg_30_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_30_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_31_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_31_MPORT_addr = 5'h1f;
  assign Regfile_reg_trace_io_input_reg_31_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_31_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_data = Regfile[Regfile_mem_wdata_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_1_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_1_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_1_data = Regfile[Regfile_mem_wdata_MPORT_1_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_2_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_2_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_2_data = Regfile[Regfile_mem_wdata_MPORT_2_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_3_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_3_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_3_data = Regfile[Regfile_mem_wdata_MPORT_3_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_MPORT_data = _T_6 ? io_res2rd : reg_value;
  assign Regfile_MPORT_addr = io_rd;
  assign Regfile_MPORT_mask = 1'h1;
  assign Regfile_MPORT_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_io_res2rd_MPORT_1_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_1_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_1_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_1_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_io_res2rd_MPORT_2_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_2_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_2_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_2_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_csr_wdata_MPORT_en = 1'h1;
  assign CSR_Reg_csr_wdata_MPORT_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_csr_wdata_MPORT_data = CSR_Reg[CSR_Reg_csr_wdata_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_csr_wdata_MPORT_1_en = 1'h1;
  assign CSR_Reg_csr_wdata_MPORT_1_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_csr_wdata_MPORT_1_data = CSR_Reg[CSR_Reg_csr_wdata_MPORT_1_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_2_en = 1'h1;
  assign CSR_Reg_MPORT_2_addr = 2'h1;
  assign CSR_Reg_MPORT_2_data = CSR_Reg[CSR_Reg_MPORT_2_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_5_en = 1'h1;
  assign CSR_Reg_MPORT_5_addr = 2'h3;
  assign CSR_Reg_MPORT_5_data = CSR_Reg[CSR_Reg_MPORT_5_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_7_en = 1'h1;
  assign CSR_Reg_MPORT_7_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_MPORT_7_data = CSR_Reg[CSR_Reg_MPORT_7_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_j_pc_MPORT_12_en = 1'h1;
  assign CSR_Reg_j_pc_MPORT_12_addr = 2'h0;
  assign CSR_Reg_j_pc_MPORT_12_data = CSR_Reg[CSR_Reg_j_pc_MPORT_12_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_j_pc_MPORT_13_en = 1'h1;
  assign CSR_Reg_j_pc_MPORT_13_addr = 2'h1;
  assign CSR_Reg_j_pc_MPORT_13_data = CSR_Reg[CSR_Reg_j_pc_MPORT_13_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr = 2'h0;
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr = 2'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr = 2'h2;
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_1_data = _T_9 ? io_pc : CSR_Reg_MPORT_2_data;
  assign CSR_Reg_MPORT_1_addr = 2'h1;
  assign CSR_Reg_MPORT_1_mask = 1'h1;
  assign CSR_Reg_MPORT_1_en = 1'h1;
  assign CSR_Reg_MPORT_3_data = _T_9 ? Regfile_MPORT_4_data : CSR_Reg_MPORT_5_data;
  assign CSR_Reg_MPORT_3_addr = 2'h3;
  assign CSR_Reg_MPORT_3_mask = 1'h1;
  assign CSR_Reg_MPORT_3_en = 1'h1;
  assign CSR_Reg_MPORT_6_data = _T_14 ? csr_wdata : CSR_Reg_MPORT_7_data;
  assign CSR_Reg_MPORT_6_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_MPORT_6_mask = 1'h1;
  assign CSR_Reg_MPORT_6_en = 1'h1;
  assign io_pc_next = pc_next; // @[EXU_AXI.scala 162:16]
  assign io_res2rd = _io_res2rd_T_208[63:0]; // @[EXU_AXI.scala 72:15]
  assign io_inst_store = io_ctrl_sign_Writemem_en; // @[EXU_AXI.scala 188:19]
  assign io_inst_load = io_ctrl_sign_Readmem_en; // @[EXU_AXI.scala 189:18]
  assign io_Mem_addr = add_res[31:0]; // @[EXU_AXI.scala 190:17]
  assign io_Mem_wdata = 32'h27 == io_inst_now ? {{32'd0}, _mem_wdata_T_9[31:0]} : _mem_wdata_T_16; // @[Mux.scala 81:58]
  assign io_Mem_wstrb = io_ctrl_sign_Wmask; // @[EXU_AXI.scala 192:18]
  assign reg_trace_input_reg_0 = Regfile_reg_trace_io_input_reg_0_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_1 = Regfile_reg_trace_io_input_reg_1_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_2 = Regfile_reg_trace_io_input_reg_2_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_3 = Regfile_reg_trace_io_input_reg_3_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_4 = Regfile_reg_trace_io_input_reg_4_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_5 = Regfile_reg_trace_io_input_reg_5_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_6 = Regfile_reg_trace_io_input_reg_6_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_7 = Regfile_reg_trace_io_input_reg_7_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_8 = Regfile_reg_trace_io_input_reg_8_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_9 = Regfile_reg_trace_io_input_reg_9_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_10 = Regfile_reg_trace_io_input_reg_10_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_11 = Regfile_reg_trace_io_input_reg_11_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_12 = Regfile_reg_trace_io_input_reg_12_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_13 = Regfile_reg_trace_io_input_reg_13_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_14 = Regfile_reg_trace_io_input_reg_14_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_15 = Regfile_reg_trace_io_input_reg_15_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_16 = Regfile_reg_trace_io_input_reg_16_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_17 = Regfile_reg_trace_io_input_reg_17_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_18 = Regfile_reg_trace_io_input_reg_18_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_19 = Regfile_reg_trace_io_input_reg_19_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_20 = Regfile_reg_trace_io_input_reg_20_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_21 = Regfile_reg_trace_io_input_reg_21_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_22 = Regfile_reg_trace_io_input_reg_22_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_23 = Regfile_reg_trace_io_input_reg_23_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_24 = Regfile_reg_trace_io_input_reg_24_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_25 = Regfile_reg_trace_io_input_reg_25_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_26 = Regfile_reg_trace_io_input_reg_26_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_27 = Regfile_reg_trace_io_input_reg_27_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_28 = Regfile_reg_trace_io_input_reg_28_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_29 = Regfile_reg_trace_io_input_reg_29_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_30 = Regfile_reg_trace_io_input_reg_30_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_31 = Regfile_reg_trace_io_input_reg_31_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_csr_reg_0 = CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_1 = CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_2 = CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_3 = 64'h0; // @[EXU_AXI.scala 167:{36,36}]
  assign reg_trace_pc = io_pc; // @[EXU_AXI.scala 166:21]
  always @(posedge clock) begin
    if (Regfile_MPORT_en & Regfile_MPORT_mask) begin
      Regfile[Regfile_MPORT_addr] <= Regfile_MPORT_data; // @[EXU_AXI.scala 37:22]
    end
    if (CSR_Reg_MPORT_1_en & CSR_Reg_MPORT_1_mask) begin
      CSR_Reg[CSR_Reg_MPORT_1_addr] <= CSR_Reg_MPORT_1_data; // @[EXU_AXI.scala 38:22]
    end
    if (CSR_Reg_MPORT_3_en & CSR_Reg_MPORT_3_mask) begin
      CSR_Reg[CSR_Reg_MPORT_3_addr] <= CSR_Reg_MPORT_3_data; // @[EXU_AXI.scala 38:22]
    end
    if (CSR_Reg_MPORT_6_en & CSR_Reg_MPORT_6_mask) begin
      CSR_Reg[CSR_Reg_MPORT_6_addr] <= CSR_Reg_MPORT_6_data; // @[EXU_AXI.scala 38:22]
    end
    if (reset) begin // @[EXU_AXI.scala 158:26]
      pc_next <= 64'h0; // @[EXU_AXI.scala 158:26]
    end else if (io_inst_valid) begin // @[EXU_AXI.scala 159:24]
      if (32'h3e == io_inst_now) begin // @[Mux.scala 81:58]
        pc_next <= _j_pc_T_46;
      end else if (32'h3d == io_inst_now) begin // @[Mux.scala 81:58]
        pc_next <= CSR_Reg_j_pc_MPORT_12_data;
      end else begin
        pc_next <= _j_pc_T_62;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    Regfile[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    CSR_Reg[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  pc_next = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top(
  input         clock,
  input         reset,
  output [31:0] io_inst,
  output [63:0] io_pc,
  output [63:0] io_pc_next,
  output [63:0] io_outval,
  output        io_step
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  axi_clock; // @[top.scala 18:21]
  wire  axi_reset; // @[top.scala 18:21]
  wire [31:0] axi_io_axi_in_araddr; // @[top.scala 18:21]
  wire  axi_io_axi_in_arvalid; // @[top.scala 18:21]
  wire  axi_io_axi_in_rready; // @[top.scala 18:21]
  wire [31:0] axi_io_axi_in_awaddr; // @[top.scala 18:21]
  wire  axi_io_axi_in_awvalid; // @[top.scala 18:21]
  wire [63:0] axi_io_axi_in_wdata; // @[top.scala 18:21]
  wire [7:0] axi_io_axi_in_wstrb; // @[top.scala 18:21]
  wire  axi_io_axi_in_wvalid; // @[top.scala 18:21]
  wire  axi_io_axi_in_bready; // @[top.scala 18:21]
  wire  axi_io_axi_out_arready; // @[top.scala 18:21]
  wire [63:0] axi_io_axi_out_rdata; // @[top.scala 18:21]
  wire  axi_io_axi_out_rvalid; // @[top.scala 18:21]
  wire  axi_io_axi_out_awready; // @[top.scala 18:21]
  wire  axi_io_axi_out_wready; // @[top.scala 18:21]
  wire  axi_io_axi_out_bvalid; // @[top.scala 18:21]
  wire  lsu_step_clock; // @[top.scala 19:26]
  wire  lsu_step_reset; // @[top.scala 19:26]
  wire  lsu_step_io_inst_store; // @[top.scala 19:26]
  wire  lsu_step_io_inst_load; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_mem_addr; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_mem_wdata; // @[top.scala 19:26]
  wire [7:0] lsu_step_io_mem_wstrb; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_mem_rdata; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_arready; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_axi_in_rdata; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_rvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_awready; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_wready; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_bvalid; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_axi_out_araddr; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_arvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_rready; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_axi_out_awaddr; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_awvalid; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_axi_out_wdata; // @[top.scala 19:26]
  wire [7:0] lsu_step_io_axi_out_wstrb; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_wvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_bready; // @[top.scala 19:26]
  wire  arbiter_clock; // @[top.scala 20:25]
  wire  arbiter_reset; // @[top.scala 20:25]
  wire [31:0] arbiter_io_ifu_axi_in_araddr; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_in_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_in_rready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_ifu_axi_out_rdata; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_out_rvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_lsu_axi_in_araddr; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_rready; // @[top.scala 20:25]
  wire [31:0] arbiter_io_lsu_axi_in_awaddr; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_awvalid; // @[top.scala 20:25]
  wire [63:0] arbiter_io_lsu_axi_in_wdata; // @[top.scala 20:25]
  wire [7:0] arbiter_io_lsu_axi_in_wstrb; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_wvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_bready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_arready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_lsu_axi_out_rdata; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_rvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_awready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_wready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_bvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_arready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_axi_in_rdata; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_rvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_awready; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_wready; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_bvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_axi_out_araddr; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_rready; // @[top.scala 20:25]
  wire [31:0] arbiter_io_axi_out_awaddr; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_awvalid; // @[top.scala 20:25]
  wire [63:0] arbiter_io_axi_out_wdata; // @[top.scala 20:25]
  wire [7:0] arbiter_io_axi_out_wstrb; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_wvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_bready; // @[top.scala 20:25]
  wire  ifu_step_clock; // @[top.scala 21:26]
  wire  ifu_step_reset; // @[top.scala 21:26]
  wire [63:0] ifu_step_io_pc; // @[top.scala 21:26]
  wire  ifu_step_io_pc_valid; // @[top.scala 21:26]
  wire  ifu_step_io_inst_valid; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_inst; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_inst_reg; // @[top.scala 21:26]
  wire [63:0] ifu_step_io_axi_in_rdata; // @[top.scala 21:26]
  wire  ifu_step_io_axi_in_rvalid; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_axi_out_araddr; // @[top.scala 21:26]
  wire  ifu_step_io_axi_out_arvalid; // @[top.scala 21:26]
  wire  ifu_step_io_axi_out_rready; // @[top.scala 21:26]
  wire  i_cache_clock; // @[top.scala 22:25]
  wire  i_cache_reset; // @[top.scala 22:25]
  wire [31:0] i_cache_io_from_ifu_araddr; // @[top.scala 22:25]
  wire  i_cache_io_from_ifu_arvalid; // @[top.scala 22:25]
  wire  i_cache_io_from_ifu_rready; // @[top.scala 22:25]
  wire [63:0] i_cache_io_to_ifu_rdata; // @[top.scala 22:25]
  wire  i_cache_io_to_ifu_rvalid; // @[top.scala 22:25]
  wire [31:0] i_cache_io_to_axi_araddr; // @[top.scala 22:25]
  wire  i_cache_io_to_axi_arvalid; // @[top.scala 22:25]
  wire  i_cache_io_to_axi_rready; // @[top.scala 22:25]
  wire [63:0] i_cache_io_from_axi_rdata; // @[top.scala 22:25]
  wire  i_cache_io_from_axi_rvalid; // @[top.scala 22:25]
  wire  d_cache_clock; // @[top.scala 23:25]
  wire  d_cache_reset; // @[top.scala 23:25]
  wire [63:0] d_cache_io_pc_now; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_araddr; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_arvalid; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_rready; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_awaddr; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_awvalid; // @[top.scala 23:25]
  wire [63:0] d_cache_io_from_lsu_wdata; // @[top.scala 23:25]
  wire [7:0] d_cache_io_from_lsu_wstrb; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_wvalid; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_bready; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_arready; // @[top.scala 23:25]
  wire [63:0] d_cache_io_to_lsu_rdata; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_rvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_awready; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_wready; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_bvalid; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_araddr; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_arvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_rready; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_awaddr; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_awvalid; // @[top.scala 23:25]
  wire [63:0] d_cache_io_to_axi_wdata; // @[top.scala 23:25]
  wire [7:0] d_cache_io_to_axi_wstrb; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_wvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_bready; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_arready; // @[top.scala 23:25]
  wire [63:0] d_cache_io_from_axi_rdata; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_rvalid; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_awready; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_wready; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_bvalid; // @[top.scala 23:25]
  wire [31:0] idu_step_io_inst; // @[top.scala 46:26]
  wire [31:0] idu_step_io_inst_now; // @[top.scala 46:26]
  wire [4:0] idu_step_io_rs1; // @[top.scala 46:26]
  wire [4:0] idu_step_io_rs2; // @[top.scala 46:26]
  wire [4:0] idu_step_io_rd; // @[top.scala 46:26]
  wire [63:0] idu_step_io_imm; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_reg_write; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_csr_write; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_Writemem_en; // @[top.scala 46:26]
  wire  idu_step_io_ctrl_sign_Readmem_en; // @[top.scala 46:26]
  wire [7:0] idu_step_io_ctrl_sign_Wmask; // @[top.scala 46:26]
  wire  exu_step_clock; // @[top.scala 51:26]
  wire  exu_step_reset; // @[top.scala 51:26]
  wire [63:0] exu_step_io_pc; // @[top.scala 51:26]
  wire [63:0] exu_step_io_pc_next; // @[top.scala 51:26]
  wire [31:0] exu_step_io_inst_now; // @[top.scala 51:26]
  wire [4:0] exu_step_io_rs1; // @[top.scala 51:26]
  wire [4:0] exu_step_io_rs2; // @[top.scala 51:26]
  wire [4:0] exu_step_io_rd; // @[top.scala 51:26]
  wire [63:0] exu_step_io_imm; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_reg_write; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_csr_write; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_Writemem_en; // @[top.scala 51:26]
  wire  exu_step_io_ctrl_sign_Readmem_en; // @[top.scala 51:26]
  wire [7:0] exu_step_io_ctrl_sign_Wmask; // @[top.scala 51:26]
  wire [63:0] exu_step_io_res2rd; // @[top.scala 51:26]
  wire  exu_step_io_inst_valid; // @[top.scala 51:26]
  wire  exu_step_io_inst_store; // @[top.scala 51:26]
  wire  exu_step_io_inst_load; // @[top.scala 51:26]
  wire [31:0] exu_step_io_Mem_addr; // @[top.scala 51:26]
  wire [63:0] exu_step_io_Mem_rdata; // @[top.scala 51:26]
  wire [63:0] exu_step_io_Mem_wdata; // @[top.scala 51:26]
  wire [7:0] exu_step_io_Mem_wstrb; // @[top.scala 51:26]
  wire  exu_step_io_rdata_valid; // @[top.scala 51:26]
  wire [31:0] dpi_flag; // @[top.scala 73:21]
  wire [31:0] dpi_ecall_flag; // @[top.scala 73:21]
  reg [63:0] pc_now; // @[top.scala 15:25]
  reg  execute_end; // @[top.scala 17:30]
  reg  pc_valid; // @[top.scala 87:27]
  reg  diff_step; // @[top.scala 90:28]
  AXI axi ( // @[top.scala 18:21]
    .clock(axi_clock),
    .reset(axi_reset),
    .io_axi_in_araddr(axi_io_axi_in_araddr),
    .io_axi_in_arvalid(axi_io_axi_in_arvalid),
    .io_axi_in_rready(axi_io_axi_in_rready),
    .io_axi_in_awaddr(axi_io_axi_in_awaddr),
    .io_axi_in_awvalid(axi_io_axi_in_awvalid),
    .io_axi_in_wdata(axi_io_axi_in_wdata),
    .io_axi_in_wstrb(axi_io_axi_in_wstrb),
    .io_axi_in_wvalid(axi_io_axi_in_wvalid),
    .io_axi_in_bready(axi_io_axi_in_bready),
    .io_axi_out_arready(axi_io_axi_out_arready),
    .io_axi_out_rdata(axi_io_axi_out_rdata),
    .io_axi_out_rvalid(axi_io_axi_out_rvalid),
    .io_axi_out_awready(axi_io_axi_out_awready),
    .io_axi_out_wready(axi_io_axi_out_wready),
    .io_axi_out_bvalid(axi_io_axi_out_bvalid)
  );
  LSU lsu_step ( // @[top.scala 19:26]
    .clock(lsu_step_clock),
    .reset(lsu_step_reset),
    .io_inst_store(lsu_step_io_inst_store),
    .io_inst_load(lsu_step_io_inst_load),
    .io_mem_addr(lsu_step_io_mem_addr),
    .io_mem_wdata(lsu_step_io_mem_wdata),
    .io_mem_wstrb(lsu_step_io_mem_wstrb),
    .io_mem_rdata(lsu_step_io_mem_rdata),
    .io_axi_in_arready(lsu_step_io_axi_in_arready),
    .io_axi_in_rdata(lsu_step_io_axi_in_rdata),
    .io_axi_in_rvalid(lsu_step_io_axi_in_rvalid),
    .io_axi_in_awready(lsu_step_io_axi_in_awready),
    .io_axi_in_wready(lsu_step_io_axi_in_wready),
    .io_axi_in_bvalid(lsu_step_io_axi_in_bvalid),
    .io_axi_out_araddr(lsu_step_io_axi_out_araddr),
    .io_axi_out_arvalid(lsu_step_io_axi_out_arvalid),
    .io_axi_out_rready(lsu_step_io_axi_out_rready),
    .io_axi_out_awaddr(lsu_step_io_axi_out_awaddr),
    .io_axi_out_awvalid(lsu_step_io_axi_out_awvalid),
    .io_axi_out_wdata(lsu_step_io_axi_out_wdata),
    .io_axi_out_wstrb(lsu_step_io_axi_out_wstrb),
    .io_axi_out_wvalid(lsu_step_io_axi_out_wvalid),
    .io_axi_out_bready(lsu_step_io_axi_out_bready)
  );
  AXI_ARBITER arbiter ( // @[top.scala 20:25]
    .clock(arbiter_clock),
    .reset(arbiter_reset),
    .io_ifu_axi_in_araddr(arbiter_io_ifu_axi_in_araddr),
    .io_ifu_axi_in_arvalid(arbiter_io_ifu_axi_in_arvalid),
    .io_ifu_axi_in_rready(arbiter_io_ifu_axi_in_rready),
    .io_ifu_axi_out_rdata(arbiter_io_ifu_axi_out_rdata),
    .io_ifu_axi_out_rvalid(arbiter_io_ifu_axi_out_rvalid),
    .io_lsu_axi_in_araddr(arbiter_io_lsu_axi_in_araddr),
    .io_lsu_axi_in_arvalid(arbiter_io_lsu_axi_in_arvalid),
    .io_lsu_axi_in_rready(arbiter_io_lsu_axi_in_rready),
    .io_lsu_axi_in_awaddr(arbiter_io_lsu_axi_in_awaddr),
    .io_lsu_axi_in_awvalid(arbiter_io_lsu_axi_in_awvalid),
    .io_lsu_axi_in_wdata(arbiter_io_lsu_axi_in_wdata),
    .io_lsu_axi_in_wstrb(arbiter_io_lsu_axi_in_wstrb),
    .io_lsu_axi_in_wvalid(arbiter_io_lsu_axi_in_wvalid),
    .io_lsu_axi_in_bready(arbiter_io_lsu_axi_in_bready),
    .io_lsu_axi_out_arready(arbiter_io_lsu_axi_out_arready),
    .io_lsu_axi_out_rdata(arbiter_io_lsu_axi_out_rdata),
    .io_lsu_axi_out_rvalid(arbiter_io_lsu_axi_out_rvalid),
    .io_lsu_axi_out_awready(arbiter_io_lsu_axi_out_awready),
    .io_lsu_axi_out_wready(arbiter_io_lsu_axi_out_wready),
    .io_lsu_axi_out_bvalid(arbiter_io_lsu_axi_out_bvalid),
    .io_axi_in_arready(arbiter_io_axi_in_arready),
    .io_axi_in_rdata(arbiter_io_axi_in_rdata),
    .io_axi_in_rvalid(arbiter_io_axi_in_rvalid),
    .io_axi_in_awready(arbiter_io_axi_in_awready),
    .io_axi_in_wready(arbiter_io_axi_in_wready),
    .io_axi_in_bvalid(arbiter_io_axi_in_bvalid),
    .io_axi_out_araddr(arbiter_io_axi_out_araddr),
    .io_axi_out_arvalid(arbiter_io_axi_out_arvalid),
    .io_axi_out_rready(arbiter_io_axi_out_rready),
    .io_axi_out_awaddr(arbiter_io_axi_out_awaddr),
    .io_axi_out_awvalid(arbiter_io_axi_out_awvalid),
    .io_axi_out_wdata(arbiter_io_axi_out_wdata),
    .io_axi_out_wstrb(arbiter_io_axi_out_wstrb),
    .io_axi_out_wvalid(arbiter_io_axi_out_wvalid),
    .io_axi_out_bready(arbiter_io_axi_out_bready)
  );
  IFU_AXI ifu_step ( // @[top.scala 21:26]
    .clock(ifu_step_clock),
    .reset(ifu_step_reset),
    .io_pc(ifu_step_io_pc),
    .io_pc_valid(ifu_step_io_pc_valid),
    .io_inst_valid(ifu_step_io_inst_valid),
    .io_inst(ifu_step_io_inst),
    .io_inst_reg(ifu_step_io_inst_reg),
    .io_axi_in_rdata(ifu_step_io_axi_in_rdata),
    .io_axi_in_rvalid(ifu_step_io_axi_in_rvalid),
    .io_axi_out_araddr(ifu_step_io_axi_out_araddr),
    .io_axi_out_arvalid(ifu_step_io_axi_out_arvalid),
    .io_axi_out_rready(ifu_step_io_axi_out_rready)
  );
  I_CACHE i_cache ( // @[top.scala 22:25]
    .clock(i_cache_clock),
    .reset(i_cache_reset),
    .io_from_ifu_araddr(i_cache_io_from_ifu_araddr),
    .io_from_ifu_arvalid(i_cache_io_from_ifu_arvalid),
    .io_from_ifu_rready(i_cache_io_from_ifu_rready),
    .io_to_ifu_rdata(i_cache_io_to_ifu_rdata),
    .io_to_ifu_rvalid(i_cache_io_to_ifu_rvalid),
    .io_to_axi_araddr(i_cache_io_to_axi_araddr),
    .io_to_axi_arvalid(i_cache_io_to_axi_arvalid),
    .io_to_axi_rready(i_cache_io_to_axi_rready),
    .io_from_axi_rdata(i_cache_io_from_axi_rdata),
    .io_from_axi_rvalid(i_cache_io_from_axi_rvalid)
  );
  D_CACHE d_cache ( // @[top.scala 23:25]
    .clock(d_cache_clock),
    .reset(d_cache_reset),
    .io_pc_now(d_cache_io_pc_now),
    .io_from_lsu_araddr(d_cache_io_from_lsu_araddr),
    .io_from_lsu_arvalid(d_cache_io_from_lsu_arvalid),
    .io_from_lsu_rready(d_cache_io_from_lsu_rready),
    .io_from_lsu_awaddr(d_cache_io_from_lsu_awaddr),
    .io_from_lsu_awvalid(d_cache_io_from_lsu_awvalid),
    .io_from_lsu_wdata(d_cache_io_from_lsu_wdata),
    .io_from_lsu_wstrb(d_cache_io_from_lsu_wstrb),
    .io_from_lsu_wvalid(d_cache_io_from_lsu_wvalid),
    .io_from_lsu_bready(d_cache_io_from_lsu_bready),
    .io_to_lsu_arready(d_cache_io_to_lsu_arready),
    .io_to_lsu_rdata(d_cache_io_to_lsu_rdata),
    .io_to_lsu_rvalid(d_cache_io_to_lsu_rvalid),
    .io_to_lsu_awready(d_cache_io_to_lsu_awready),
    .io_to_lsu_wready(d_cache_io_to_lsu_wready),
    .io_to_lsu_bvalid(d_cache_io_to_lsu_bvalid),
    .io_to_axi_araddr(d_cache_io_to_axi_araddr),
    .io_to_axi_arvalid(d_cache_io_to_axi_arvalid),
    .io_to_axi_rready(d_cache_io_to_axi_rready),
    .io_to_axi_awaddr(d_cache_io_to_axi_awaddr),
    .io_to_axi_awvalid(d_cache_io_to_axi_awvalid),
    .io_to_axi_wdata(d_cache_io_to_axi_wdata),
    .io_to_axi_wstrb(d_cache_io_to_axi_wstrb),
    .io_to_axi_wvalid(d_cache_io_to_axi_wvalid),
    .io_to_axi_bready(d_cache_io_to_axi_bready),
    .io_from_axi_arready(d_cache_io_from_axi_arready),
    .io_from_axi_rdata(d_cache_io_from_axi_rdata),
    .io_from_axi_rvalid(d_cache_io_from_axi_rvalid),
    .io_from_axi_awready(d_cache_io_from_axi_awready),
    .io_from_axi_wready(d_cache_io_from_axi_wready),
    .io_from_axi_bvalid(d_cache_io_from_axi_bvalid)
  );
  IDU idu_step ( // @[top.scala 46:26]
    .io_inst(idu_step_io_inst),
    .io_inst_now(idu_step_io_inst_now),
    .io_rs1(idu_step_io_rs1),
    .io_rs2(idu_step_io_rs2),
    .io_rd(idu_step_io_rd),
    .io_imm(idu_step_io_imm),
    .io_ctrl_sign_reg_write(idu_step_io_ctrl_sign_reg_write),
    .io_ctrl_sign_csr_write(idu_step_io_ctrl_sign_csr_write),
    .io_ctrl_sign_src2_is_imm(idu_step_io_ctrl_sign_src2_is_imm),
    .io_ctrl_sign_src1_is_pc(idu_step_io_ctrl_sign_src1_is_pc),
    .io_ctrl_sign_Writemem_en(idu_step_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(idu_step_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(idu_step_io_ctrl_sign_Wmask)
  );
  EXU_AXI exu_step ( // @[top.scala 51:26]
    .clock(exu_step_clock),
    .reset(exu_step_reset),
    .io_pc(exu_step_io_pc),
    .io_pc_next(exu_step_io_pc_next),
    .io_inst_now(exu_step_io_inst_now),
    .io_rs1(exu_step_io_rs1),
    .io_rs2(exu_step_io_rs2),
    .io_rd(exu_step_io_rd),
    .io_imm(exu_step_io_imm),
    .io_ctrl_sign_reg_write(exu_step_io_ctrl_sign_reg_write),
    .io_ctrl_sign_csr_write(exu_step_io_ctrl_sign_csr_write),
    .io_ctrl_sign_src2_is_imm(exu_step_io_ctrl_sign_src2_is_imm),
    .io_ctrl_sign_src1_is_pc(exu_step_io_ctrl_sign_src1_is_pc),
    .io_ctrl_sign_Writemem_en(exu_step_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(exu_step_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(exu_step_io_ctrl_sign_Wmask),
    .io_res2rd(exu_step_io_res2rd),
    .io_inst_valid(exu_step_io_inst_valid),
    .io_inst_store(exu_step_io_inst_store),
    .io_inst_load(exu_step_io_inst_load),
    .io_Mem_addr(exu_step_io_Mem_addr),
    .io_Mem_rdata(exu_step_io_Mem_rdata),
    .io_Mem_wdata(exu_step_io_Mem_wdata),
    .io_Mem_wstrb(exu_step_io_Mem_wstrb),
    .io_rdata_valid(exu_step_io_rdata_valid)
  );
  DPI dpi ( // @[top.scala 73:21]
    .flag(dpi_flag),
    .ecall_flag(dpi_ecall_flag)
  );
  assign io_inst = ifu_step_io_inst; // @[top.scala 25:13]
  assign io_pc = pc_now; // @[top.scala 16:11]
  assign io_pc_next = exu_step_io_pc_next; // @[top.scala 94:16]
  assign io_outval = exu_step_io_res2rd; // @[top.scala 69:15]
  assign io_step = diff_step; // @[top.scala 92:13]
  assign axi_clock = clock;
  assign axi_reset = reset;
  assign axi_io_axi_in_araddr = arbiter_io_axi_out_araddr; // @[top.scala 43:19]
  assign axi_io_axi_in_arvalid = arbiter_io_axi_out_arvalid; // @[top.scala 43:19]
  assign axi_io_axi_in_rready = arbiter_io_axi_out_rready; // @[top.scala 43:19]
  assign axi_io_axi_in_awaddr = arbiter_io_axi_out_awaddr; // @[top.scala 43:19]
  assign axi_io_axi_in_awvalid = arbiter_io_axi_out_awvalid; // @[top.scala 43:19]
  assign axi_io_axi_in_wdata = arbiter_io_axi_out_wdata; // @[top.scala 43:19]
  assign axi_io_axi_in_wstrb = arbiter_io_axi_out_wstrb; // @[top.scala 43:19]
  assign axi_io_axi_in_wvalid = arbiter_io_axi_out_wvalid; // @[top.scala 43:19]
  assign axi_io_axi_in_bready = arbiter_io_axi_out_bready; // @[top.scala 43:19]
  assign lsu_step_clock = clock;
  assign lsu_step_reset = reset;
  assign lsu_step_io_inst_store = exu_step_io_inst_store; // @[top.scala 61:28]
  assign lsu_step_io_inst_load = exu_step_io_inst_load; // @[top.scala 60:27]
  assign lsu_step_io_mem_addr = exu_step_io_Mem_addr; // @[top.scala 62:26]
  assign lsu_step_io_mem_wdata = exu_step_io_Mem_wdata; // @[top.scala 63:27]
  assign lsu_step_io_mem_wstrb = exu_step_io_Mem_wstrb; // @[top.scala 64:27]
  assign lsu_step_io_axi_in_arready = d_cache_io_to_lsu_arready; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_rdata = d_cache_io_to_lsu_rdata; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_rvalid = d_cache_io_to_lsu_rvalid; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_awready = d_cache_io_to_lsu_awready; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_wready = d_cache_io_to_lsu_wready; // @[top.scala 36:24]
  assign lsu_step_io_axi_in_bvalid = d_cache_io_to_lsu_bvalid; // @[top.scala 36:24]
  assign arbiter_clock = clock;
  assign arbiter_reset = reset;
  assign arbiter_io_ifu_axi_in_araddr = i_cache_io_to_axi_araddr; // @[top.scala 26:27]
  assign arbiter_io_ifu_axi_in_arvalid = i_cache_io_to_axi_arvalid; // @[top.scala 26:27]
  assign arbiter_io_ifu_axi_in_rready = i_cache_io_to_axi_rready; // @[top.scala 26:27]
  assign arbiter_io_lsu_axi_in_araddr = d_cache_io_to_axi_araddr; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_arvalid = d_cache_io_to_axi_arvalid; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_rready = d_cache_io_to_axi_rready; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_awaddr = d_cache_io_to_axi_awaddr; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_awvalid = d_cache_io_to_axi_awvalid; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_wdata = d_cache_io_to_axi_wdata; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_wstrb = d_cache_io_to_axi_wstrb; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_wvalid = d_cache_io_to_axi_wvalid; // @[top.scala 34:27]
  assign arbiter_io_lsu_axi_in_bready = d_cache_io_to_axi_bready; // @[top.scala 34:27]
  assign arbiter_io_axi_in_arready = axi_io_axi_out_arready; // @[top.scala 42:23]
  assign arbiter_io_axi_in_rdata = axi_io_axi_out_rdata; // @[top.scala 42:23]
  assign arbiter_io_axi_in_rvalid = axi_io_axi_out_rvalid; // @[top.scala 42:23]
  assign arbiter_io_axi_in_awready = axi_io_axi_out_awready; // @[top.scala 42:23]
  assign arbiter_io_axi_in_wready = axi_io_axi_out_wready; // @[top.scala 42:23]
  assign arbiter_io_axi_in_bvalid = axi_io_axi_out_bvalid; // @[top.scala 42:23]
  assign ifu_step_clock = clock;
  assign ifu_step_reset = reset;
  assign ifu_step_io_pc = pc_now; // @[top.scala 24:20]
  assign ifu_step_io_pc_valid = pc_valid; // @[top.scala 89:26]
  assign ifu_step_io_axi_in_rdata = i_cache_io_to_ifu_rdata; // @[top.scala 28:24]
  assign ifu_step_io_axi_in_rvalid = i_cache_io_to_ifu_rvalid; // @[top.scala 28:24]
  assign i_cache_clock = clock;
  assign i_cache_reset = reset;
  assign i_cache_io_from_ifu_araddr = ifu_step_io_axi_out_araddr; // @[top.scala 29:25]
  assign i_cache_io_from_ifu_arvalid = ifu_step_io_axi_out_arvalid; // @[top.scala 29:25]
  assign i_cache_io_from_ifu_rready = ifu_step_io_axi_out_rready; // @[top.scala 29:25]
  assign i_cache_io_from_axi_rdata = arbiter_io_ifu_axi_out_rdata; // @[top.scala 27:25]
  assign i_cache_io_from_axi_rvalid = arbiter_io_ifu_axi_out_rvalid; // @[top.scala 27:25]
  assign d_cache_clock = clock;
  assign d_cache_reset = reset;
  assign d_cache_io_pc_now = pc_now; // @[top.scala 38:23]
  assign d_cache_io_from_lsu_araddr = lsu_step_io_axi_out_araddr; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_arvalid = lsu_step_io_axi_out_arvalid; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_rready = lsu_step_io_axi_out_rready; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_awaddr = lsu_step_io_axi_out_awaddr; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_awvalid = lsu_step_io_axi_out_awvalid; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_wdata = lsu_step_io_axi_out_wdata; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_wstrb = lsu_step_io_axi_out_wstrb; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_wvalid = lsu_step_io_axi_out_wvalid; // @[top.scala 37:25]
  assign d_cache_io_from_lsu_bready = lsu_step_io_axi_out_bready; // @[top.scala 37:25]
  assign d_cache_io_from_axi_arready = arbiter_io_lsu_axi_out_arready; // @[top.scala 35:25]
  assign d_cache_io_from_axi_rdata = arbiter_io_lsu_axi_out_rdata; // @[top.scala 35:25]
  assign d_cache_io_from_axi_rvalid = arbiter_io_lsu_axi_out_rvalid; // @[top.scala 35:25]
  assign d_cache_io_from_axi_awready = arbiter_io_lsu_axi_out_awready; // @[top.scala 35:25]
  assign d_cache_io_from_axi_wready = arbiter_io_lsu_axi_out_wready; // @[top.scala 35:25]
  assign d_cache_io_from_axi_bvalid = arbiter_io_lsu_axi_out_bvalid; // @[top.scala 35:25]
  assign idu_step_io_inst = ~ifu_step_io_inst_valid & ~pc_valid & ~execute_end ? ifu_step_io_inst_reg : ifu_step_io_inst
    ; // @[top.scala 96:28]
  assign exu_step_clock = clock;
  assign exu_step_reset = reset;
  assign exu_step_io_pc = pc_now; // @[top.scala 52:20]
  assign exu_step_io_inst_now = idu_step_io_inst_now; // @[top.scala 53:26]
  assign exu_step_io_rs1 = idu_step_io_rs1; // @[top.scala 55:21]
  assign exu_step_io_rs2 = idu_step_io_rs2; // @[top.scala 56:21]
  assign exu_step_io_rd = idu_step_io_rd; // @[top.scala 57:20]
  assign exu_step_io_imm = idu_step_io_imm; // @[top.scala 58:21]
  assign exu_step_io_ctrl_sign_reg_write = idu_step_io_ctrl_sign_reg_write; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_csr_write = idu_step_io_ctrl_sign_csr_write; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_src2_is_imm = idu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_src1_is_pc = idu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_Writemem_en = idu_step_io_ctrl_sign_Writemem_en; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_Readmem_en = idu_step_io_ctrl_sign_Readmem_en; // @[top.scala 59:27]
  assign exu_step_io_ctrl_sign_Wmask = idu_step_io_ctrl_sign_Wmask; // @[top.scala 59:27]
  assign exu_step_io_inst_valid = ifu_step_io_inst_valid; // @[top.scala 68:28]
  assign exu_step_io_Mem_rdata = lsu_step_io_mem_rdata; // @[top.scala 65:27]
  assign exu_step_io_rdata_valid = lsu_step_io_axi_in_rvalid; // @[top.scala 66:29]
  assign dpi_flag = {{31'd0}, idu_step_io_inst_now == 32'h2}; // @[top.scala 74:17]
  assign dpi_ecall_flag = {{31'd0}, idu_step_io_inst_now == 32'h3d}; // @[top.scala 75:23]
  always @(posedge clock) begin
    if (reset) begin // @[top.scala 15:25]
      pc_now <= 64'h80000000; // @[top.scala 15:25]
    end else if (execute_end) begin // @[top.scala 93:18]
      pc_now <= exu_step_io_pc_next;
    end
    if (reset) begin // @[top.scala 17:30]
      execute_end <= 1'h0; // @[top.scala 17:30]
    end else if (exu_step_io_inst_store) begin // @[top.scala 85:23]
      execute_end <= lsu_step_io_axi_in_bvalid;
    end else if (exu_step_io_inst_load) begin // @[top.scala 85:76]
      execute_end <= lsu_step_io_axi_in_rvalid;
    end else begin
      execute_end <= ifu_step_io_inst_valid;
    end
    pc_valid <= reset | execute_end; // @[top.scala 87:{27,27} 88:14]
    if (reset) begin // @[top.scala 90:28]
      diff_step <= 1'h0; // @[top.scala 90:28]
    end else begin
      diff_step <= execute_end; // @[top.scala 91:15]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"pc : %x inst:%x execute_end : %d\n\n",pc_now,idu_step_io_inst,execute_end); // @[top.scala 86:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc_now = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  execute_end = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pc_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  diff_step = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
